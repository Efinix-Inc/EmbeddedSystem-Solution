// Generator : SpinalHDL dev    git head : 81793df2c4f55a20f7eff1130c4bb74a4b11319f
// Component : EfxDMA

`timescale 1ns/1ps

module EfxDMA (
  input  wire [13:0]   ctrl_PADDR,
  input  wire [0:0]    ctrl_PSEL,
  input  wire          ctrl_PENABLE,
  output wire          ctrl_PREADY,
  input  wire          ctrl_PWRITE,
  input  wire [31:0]   ctrl_PWDATA,
  output wire [31:0]   ctrl_PRDATA,
  output wire          ctrl_PSLVERROR,
  output wire [3:0]    ctrl_interrupts,
  output wire          read_arvalid,
  input  wire          read_arready,
  output wire [31:0]   read_araddr,
  output wire [3:0]    read_arregion,
  output wire [7:0]    read_arlen,
  output wire [2:0]    read_arsize,
  output wire [1:0]    read_arburst,
  output wire [0:0]    read_arlock,
  output wire [3:0]    read_arcache,
  output wire [3:0]    read_arqos,
  output wire [2:0]    read_arprot,
  input  wire          read_rvalid,
  output wire          read_rready,
  input  wire [255:0]  read_rdata,
  input  wire [1:0]    read_rresp,
  input  wire          read_rlast,
  output wire          write_awvalid,
  input  wire          write_awready,
  output wire [31:0]   write_awaddr,
  output wire [3:0]    write_awregion,
  output wire [7:0]    write_awlen,
  output wire [2:0]    write_awsize,
  output wire [1:0]    write_awburst,
  output wire [0:0]    write_awlock,
  output wire [3:0]    write_awcache,
  output wire [3:0]    write_awqos,
  output wire [2:0]    write_awprot,
  output wire          write_wvalid,
  input  wire          write_wready,
  output wire [255:0]  write_wdata,
  output wire [31:0]   write_wstrb,
  output wire          write_wlast,
  input  wire          write_bvalid,
  output wire          write_bready,
  input  wire [1:0]    write_bresp,
  input  wire          dat0_i_tvalid,
  output wire          dat0_i_tready,
  input  wire [63:0]   dat0_i_tdata,
  input  wire [7:0]    dat0_i_tkeep,
  input  wire [3:0]    dat0_i_tdest,
  input  wire          dat0_i_tlast,
  input  wire          dat2_i_tvalid,
  output wire          dat2_i_tready,
  input  wire [31:0]   dat2_i_tdata,
  input  wire [3:0]    dat2_i_tkeep,
  input  wire [3:0]    dat2_i_tdest,
  input  wire          dat2_i_tlast,
  output wire          dat1_o_tvalid,
  input  wire          dat1_o_tready,
  output wire [63:0]   dat1_o_tdata,
  output wire [7:0]    dat1_o_tkeep,
  output wire [3:0]    dat1_o_tdest,
  output wire          dat1_o_tlast,
  output wire          dat3_o_tvalid,
  input  wire          dat3_o_tready,
  output wire [31:0]   dat3_o_tdata,
  output wire [3:0]    dat3_o_tkeep,
  output wire [3:0]    dat3_o_tdest,
  output wire          dat3_o_tlast,
  input  wire          clk,
  input  wire          reset,
  input  wire          ctrl_clk,
  input  wire          ctrl_reset,
  input  wire          dat0_i_clk,
  input  wire          dat0_i_reset,
  input  wire          dat2_i_clk,
  input  wire          dat2_i_reset,
  input  wire          dat1_o_clk,
  input  wire          dat1_o_reset,
  input  wire          dat3_o_clk,
  input  wire          dat3_o_reset
);

  wire                core_io_read_cmd_valid;
  wire                core_io_read_cmd_payload_last;
  wire       [0:0]    core_io_read_cmd_payload_fragment_source;
  wire       [0:0]    core_io_read_cmd_payload_fragment_opcode;
  wire       [31:0]   core_io_read_cmd_payload_fragment_address;
  wire       [12:0]   core_io_read_cmd_payload_fragment_length;
  wire       [24:0]   core_io_read_cmd_payload_fragment_context;
  wire                core_io_read_rsp_ready;
  wire                core_io_write_cmd_valid;
  wire                core_io_write_cmd_payload_last;
  wire       [0:0]    core_io_write_cmd_payload_fragment_source;
  wire       [0:0]    core_io_write_cmd_payload_fragment_opcode;
  wire       [31:0]   core_io_write_cmd_payload_fragment_address;
  wire       [12:0]   core_io_write_cmd_payload_fragment_length;
  wire       [255:0]  core_io_write_cmd_payload_fragment_data;
  wire       [31:0]   core_io_write_cmd_payload_fragment_mask;
  wire       [14:0]   core_io_write_cmd_payload_fragment_context;
  wire                core_io_write_rsp_ready;
  wire                core_io_outputs_0_valid;
  wire       [127:0]  core_io_outputs_0_payload_data;
  wire       [15:0]   core_io_outputs_0_payload_mask;
  wire       [3:0]    core_io_outputs_0_payload_sink;
  wire                core_io_outputs_0_payload_last;
  wire                core_io_outputs_1_valid;
  wire       [127:0]  core_io_outputs_1_payload_data;
  wire       [15:0]   core_io_outputs_1_payload_mask;
  wire       [3:0]    core_io_outputs_1_payload_sink;
  wire                core_io_outputs_1_payload_last;
  wire                core_io_inputs_0_ready;
  wire                core_io_inputs_1_ready;
  wire       [3:0]    core_io_interrupts;
  wire                core_io_ctrl_PREADY;
  wire       [31:0]   core_io_ctrl_PRDATA;
  wire                core_io_ctrl_PSLVERROR;
  wire                withCtrlCc_apbCc_io_input_PREADY;
  wire       [31:0]   withCtrlCc_apbCc_io_input_PRDATA;
  wire                withCtrlCc_apbCc_io_input_PSLVERROR;
  wire       [13:0]   withCtrlCc_apbCc_io_output_PADDR;
  wire       [0:0]    withCtrlCc_apbCc_io_output_PSEL;
  wire                withCtrlCc_apbCc_io_output_PENABLE;
  wire                withCtrlCc_apbCc_io_output_PWRITE;
  wire       [31:0]   withCtrlCc_apbCc_io_output_PWDATA;
  wire       [3:0]    io_interrupts_buffercc_io_dataOut;
  wire                readLogic_sourceRemover_io_input_cmd_ready;
  wire                readLogic_sourceRemover_io_input_rsp_valid;
  wire                readLogic_sourceRemover_io_input_rsp_payload_last;
  wire       [0:0]    readLogic_sourceRemover_io_input_rsp_payload_fragment_source;
  wire       [0:0]    readLogic_sourceRemover_io_input_rsp_payload_fragment_opcode;
  wire       [255:0]  readLogic_sourceRemover_io_input_rsp_payload_fragment_data;
  wire       [24:0]   readLogic_sourceRemover_io_input_rsp_payload_fragment_context;
  wire                readLogic_sourceRemover_io_output_cmd_valid;
  wire                readLogic_sourceRemover_io_output_cmd_payload_last;
  wire       [0:0]    readLogic_sourceRemover_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   readLogic_sourceRemover_io_output_cmd_payload_fragment_address;
  wire       [12:0]   readLogic_sourceRemover_io_output_cmd_payload_fragment_length;
  wire       [25:0]   readLogic_sourceRemover_io_output_cmd_payload_fragment_context;
  wire                readLogic_sourceRemover_io_output_rsp_ready;
  wire                readLogic_bridge_io_input_cmd_ready;
  wire                readLogic_bridge_io_input_rsp_valid;
  wire                readLogic_bridge_io_input_rsp_payload_last;
  wire       [0:0]    readLogic_bridge_io_input_rsp_payload_fragment_opcode;
  wire       [255:0]  readLogic_bridge_io_input_rsp_payload_fragment_data;
  wire       [25:0]   readLogic_bridge_io_input_rsp_payload_fragment_context;
  wire                readLogic_bridge_io_output_ar_valid;
  wire       [31:0]   readLogic_bridge_io_output_ar_payload_addr;
  wire       [7:0]    readLogic_bridge_io_output_ar_payload_len;
  wire       [2:0]    readLogic_bridge_io_output_ar_payload_size;
  wire       [3:0]    readLogic_bridge_io_output_ar_payload_cache;
  wire       [2:0]    readLogic_bridge_io_output_ar_payload_prot;
  wire                readLogic_bridge_io_output_r_ready;
  wire                writeLogic_sourceRemover_io_input_cmd_ready;
  wire                writeLogic_sourceRemover_io_input_rsp_valid;
  wire                writeLogic_sourceRemover_io_input_rsp_payload_last;
  wire       [0:0]    writeLogic_sourceRemover_io_input_rsp_payload_fragment_source;
  wire       [0:0]    writeLogic_sourceRemover_io_input_rsp_payload_fragment_opcode;
  wire       [14:0]   writeLogic_sourceRemover_io_input_rsp_payload_fragment_context;
  wire                writeLogic_sourceRemover_io_output_cmd_valid;
  wire                writeLogic_sourceRemover_io_output_cmd_payload_last;
  wire       [0:0]    writeLogic_sourceRemover_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   writeLogic_sourceRemover_io_output_cmd_payload_fragment_address;
  wire       [12:0]   writeLogic_sourceRemover_io_output_cmd_payload_fragment_length;
  wire       [255:0]  writeLogic_sourceRemover_io_output_cmd_payload_fragment_data;
  wire       [31:0]   writeLogic_sourceRemover_io_output_cmd_payload_fragment_mask;
  wire       [15:0]   writeLogic_sourceRemover_io_output_cmd_payload_fragment_context;
  wire                writeLogic_sourceRemover_io_output_rsp_ready;
  wire                writeLogic_bridge_io_input_cmd_ready;
  wire                writeLogic_bridge_io_input_rsp_valid;
  wire                writeLogic_bridge_io_input_rsp_payload_last;
  wire       [0:0]    writeLogic_bridge_io_input_rsp_payload_fragment_opcode;
  wire       [15:0]   writeLogic_bridge_io_input_rsp_payload_fragment_context;
  wire                writeLogic_bridge_io_output_aw_valid;
  wire       [31:0]   writeLogic_bridge_io_output_aw_payload_addr;
  wire       [7:0]    writeLogic_bridge_io_output_aw_payload_len;
  wire       [2:0]    writeLogic_bridge_io_output_aw_payload_size;
  wire       [3:0]    writeLogic_bridge_io_output_aw_payload_cache;
  wire       [2:0]    writeLogic_bridge_io_output_aw_payload_prot;
  wire                writeLogic_bridge_io_output_w_valid;
  wire       [255:0]  writeLogic_bridge_io_output_w_payload_data;
  wire       [31:0]   writeLogic_bridge_io_output_w_payload_strb;
  wire                writeLogic_bridge_io_output_w_payload_last;
  wire                writeLogic_bridge_io_output_b_ready;
  wire                inputsAdapter_0_upsizer_logic_io_input_ready;
  wire                inputsAdapter_0_upsizer_logic_io_output_valid;
  wire       [127:0]  inputsAdapter_0_upsizer_logic_io_output_payload_data;
  wire       [15:0]   inputsAdapter_0_upsizer_logic_io_output_payload_mask;
  wire       [3:0]    inputsAdapter_0_upsizer_logic_io_output_payload_sink;
  wire                inputsAdapter_0_upsizer_logic_io_output_payload_last;
  wire                inputsAdapter_0_crossclock_fifo_io_push_ready;
  wire                inputsAdapter_0_crossclock_fifo_io_pop_valid;
  wire       [127:0]  inputsAdapter_0_crossclock_fifo_io_pop_payload_data;
  wire       [15:0]   inputsAdapter_0_crossclock_fifo_io_pop_payload_mask;
  wire       [3:0]    inputsAdapter_0_crossclock_fifo_io_pop_payload_sink;
  wire                inputsAdapter_0_crossclock_fifo_io_pop_payload_last;
  wire       [4:0]    inputsAdapter_0_crossclock_fifo_io_pushOccupancy;
  wire       [4:0]    inputsAdapter_0_crossclock_fifo_io_popOccupancy;
  wire                inputsAdapter_1_upsizer_logic_io_input_ready;
  wire                inputsAdapter_1_upsizer_logic_io_output_valid;
  wire       [127:0]  inputsAdapter_1_upsizer_logic_io_output_payload_data;
  wire       [15:0]   inputsAdapter_1_upsizer_logic_io_output_payload_mask;
  wire       [3:0]    inputsAdapter_1_upsizer_logic_io_output_payload_sink;
  wire                inputsAdapter_1_upsizer_logic_io_output_payload_last;
  wire                inputsAdapter_1_crossclock_fifo_io_push_ready;
  wire                inputsAdapter_1_crossclock_fifo_io_pop_valid;
  wire       [127:0]  inputsAdapter_1_crossclock_fifo_io_pop_payload_data;
  wire       [15:0]   inputsAdapter_1_crossclock_fifo_io_pop_payload_mask;
  wire       [3:0]    inputsAdapter_1_crossclock_fifo_io_pop_payload_sink;
  wire                inputsAdapter_1_crossclock_fifo_io_pop_payload_last;
  wire       [4:0]    inputsAdapter_1_crossclock_fifo_io_pushOccupancy;
  wire       [4:0]    inputsAdapter_1_crossclock_fifo_io_popOccupancy;
  wire                outputsAdapter_0_crossclock_fifo_io_push_ready;
  wire                outputsAdapter_0_crossclock_fifo_io_pop_valid;
  wire       [127:0]  outputsAdapter_0_crossclock_fifo_io_pop_payload_data;
  wire       [15:0]   outputsAdapter_0_crossclock_fifo_io_pop_payload_mask;
  wire       [3:0]    outputsAdapter_0_crossclock_fifo_io_pop_payload_sink;
  wire                outputsAdapter_0_crossclock_fifo_io_pop_payload_last;
  wire       [4:0]    outputsAdapter_0_crossclock_fifo_io_pushOccupancy;
  wire       [4:0]    outputsAdapter_0_crossclock_fifo_io_popOccupancy;
  wire                outputsAdapter_0_sparseDownsizer_logic_io_input_ready;
  wire                outputsAdapter_0_sparseDownsizer_logic_io_output_valid;
  wire       [63:0]   outputsAdapter_0_sparseDownsizer_logic_io_output_payload_data;
  wire       [7:0]    outputsAdapter_0_sparseDownsizer_logic_io_output_payload_mask;
  wire       [3:0]    outputsAdapter_0_sparseDownsizer_logic_io_output_payload_sink;
  wire                outputsAdapter_0_sparseDownsizer_logic_io_output_payload_last;
  wire                outputsAdapter_1_crossclock_fifo_io_push_ready;
  wire                outputsAdapter_1_crossclock_fifo_io_pop_valid;
  wire       [127:0]  outputsAdapter_1_crossclock_fifo_io_pop_payload_data;
  wire       [15:0]   outputsAdapter_1_crossclock_fifo_io_pop_payload_mask;
  wire       [3:0]    outputsAdapter_1_crossclock_fifo_io_pop_payload_sink;
  wire                outputsAdapter_1_crossclock_fifo_io_pop_payload_last;
  wire       [4:0]    outputsAdapter_1_crossclock_fifo_io_pushOccupancy;
  wire       [4:0]    outputsAdapter_1_crossclock_fifo_io_popOccupancy;
  wire                outputsAdapter_1_sparseDownsizer_logic_io_input_ready;
  wire                outputsAdapter_1_sparseDownsizer_logic_io_output_valid;
  wire       [31:0]   outputsAdapter_1_sparseDownsizer_logic_io_output_payload_data;
  wire       [3:0]    outputsAdapter_1_sparseDownsizer_logic_io_output_payload_mask;
  wire       [3:0]    outputsAdapter_1_sparseDownsizer_logic_io_output_payload_sink;
  wire                outputsAdapter_1_sparseDownsizer_logic_io_output_payload_last;
  wire                io_write_cmd_s2mPipe_valid;
  reg                 io_write_cmd_s2mPipe_ready;
  wire                io_write_cmd_s2mPipe_payload_last;
  wire       [0:0]    io_write_cmd_s2mPipe_payload_fragment_source;
  wire       [0:0]    io_write_cmd_s2mPipe_payload_fragment_opcode;
  wire       [31:0]   io_write_cmd_s2mPipe_payload_fragment_address;
  wire       [12:0]   io_write_cmd_s2mPipe_payload_fragment_length;
  wire       [255:0]  io_write_cmd_s2mPipe_payload_fragment_data;
  wire       [31:0]   io_write_cmd_s2mPipe_payload_fragment_mask;
  wire       [14:0]   io_write_cmd_s2mPipe_payload_fragment_context;
  reg                 io_write_cmd_rValidN;
  reg                 io_write_cmd_rData_last;
  reg        [0:0]    io_write_cmd_rData_fragment_source;
  reg        [0:0]    io_write_cmd_rData_fragment_opcode;
  reg        [31:0]   io_write_cmd_rData_fragment_address;
  reg        [12:0]   io_write_cmd_rData_fragment_length;
  reg        [255:0]  io_write_cmd_rData_fragment_data;
  reg        [31:0]   io_write_cmd_rData_fragment_mask;
  reg        [14:0]   io_write_cmd_rData_fragment_context;
  wire                io_write_cmd_s2mPipe_m2sPipe_valid;
  wire                io_write_cmd_s2mPipe_m2sPipe_ready;
  wire                io_write_cmd_s2mPipe_m2sPipe_payload_last;
  wire       [0:0]    io_write_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  wire       [0:0]    io_write_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   io_write_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  wire       [12:0]   io_write_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  wire       [255:0]  io_write_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  wire       [31:0]   io_write_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  wire       [14:0]   io_write_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  reg                 io_write_cmd_s2mPipe_rValid;
  reg                 io_write_cmd_s2mPipe_rData_last;
  reg        [0:0]    io_write_cmd_s2mPipe_rData_fragment_source;
  reg        [0:0]    io_write_cmd_s2mPipe_rData_fragment_opcode;
  reg        [31:0]   io_write_cmd_s2mPipe_rData_fragment_address;
  reg        [12:0]   io_write_cmd_s2mPipe_rData_fragment_length;
  reg        [255:0]  io_write_cmd_s2mPipe_rData_fragment_data;
  reg        [31:0]   io_write_cmd_s2mPipe_rData_fragment_mask;
  reg        [14:0]   io_write_cmd_s2mPipe_rData_fragment_context;
  wire                when_Stream_l375;
  wire                interconnect_read_aggregated_cmd_valid;
  wire                interconnect_read_aggregated_cmd_ready;
  wire                interconnect_read_aggregated_cmd_payload_last;
  wire       [0:0]    interconnect_read_aggregated_cmd_payload_fragment_source;
  wire       [0:0]    interconnect_read_aggregated_cmd_payload_fragment_opcode;
  wire       [31:0]   interconnect_read_aggregated_cmd_payload_fragment_address;
  wire       [12:0]   interconnect_read_aggregated_cmd_payload_fragment_length;
  wire       [24:0]   interconnect_read_aggregated_cmd_payload_fragment_context;
  wire                interconnect_read_aggregated_rsp_valid;
  wire                interconnect_read_aggregated_rsp_ready;
  wire                interconnect_read_aggregated_rsp_payload_last;
  wire       [0:0]    interconnect_read_aggregated_rsp_payload_fragment_source;
  wire       [0:0]    interconnect_read_aggregated_rsp_payload_fragment_opcode;
  wire       [255:0]  interconnect_read_aggregated_rsp_payload_fragment_data;
  wire       [24:0]   interconnect_read_aggregated_rsp_payload_fragment_context;
  wire                interconnect_write_aggregated_cmd_valid;
  reg                 interconnect_write_aggregated_cmd_ready;
  wire                interconnect_write_aggregated_cmd_payload_last;
  wire       [0:0]    interconnect_write_aggregated_cmd_payload_fragment_source;
  wire       [0:0]    interconnect_write_aggregated_cmd_payload_fragment_opcode;
  wire       [31:0]   interconnect_write_aggregated_cmd_payload_fragment_address;
  wire       [12:0]   interconnect_write_aggregated_cmd_payload_fragment_length;
  wire       [255:0]  interconnect_write_aggregated_cmd_payload_fragment_data;
  wire       [31:0]   interconnect_write_aggregated_cmd_payload_fragment_mask;
  wire       [14:0]   interconnect_write_aggregated_cmd_payload_fragment_context;
  wire                interconnect_write_aggregated_rsp_valid;
  wire                interconnect_write_aggregated_rsp_ready;
  wire                interconnect_write_aggregated_rsp_payload_last;
  wire       [0:0]    interconnect_write_aggregated_rsp_payload_fragment_source;
  wire       [0:0]    interconnect_write_aggregated_rsp_payload_fragment_opcode;
  wire       [14:0]   interconnect_write_aggregated_rsp_payload_fragment_context;
  wire                readLogic_resized_cmd_valid;
  wire                readLogic_resized_cmd_ready;
  wire                readLogic_resized_cmd_payload_last;
  wire       [0:0]    readLogic_resized_cmd_payload_fragment_source;
  wire       [0:0]    readLogic_resized_cmd_payload_fragment_opcode;
  wire       [31:0]   readLogic_resized_cmd_payload_fragment_address;
  wire       [12:0]   readLogic_resized_cmd_payload_fragment_length;
  wire       [24:0]   readLogic_resized_cmd_payload_fragment_context;
  wire                readLogic_resized_rsp_valid;
  wire                readLogic_resized_rsp_ready;
  wire                readLogic_resized_rsp_payload_last;
  wire       [0:0]    readLogic_resized_rsp_payload_fragment_source;
  wire       [0:0]    readLogic_resized_rsp_payload_fragment_opcode;
  wire       [255:0]  readLogic_resized_rsp_payload_fragment_data;
  wire       [24:0]   readLogic_resized_rsp_payload_fragment_context;
  wire                interconnect_read_aggregated_cmd_halfPipe_valid;
  wire                interconnect_read_aggregated_cmd_halfPipe_ready;
  wire                interconnect_read_aggregated_cmd_halfPipe_payload_last;
  wire       [0:0]    interconnect_read_aggregated_cmd_halfPipe_payload_fragment_source;
  wire       [0:0]    interconnect_read_aggregated_cmd_halfPipe_payload_fragment_opcode;
  wire       [31:0]   interconnect_read_aggregated_cmd_halfPipe_payload_fragment_address;
  wire       [12:0]   interconnect_read_aggregated_cmd_halfPipe_payload_fragment_length;
  wire       [24:0]   interconnect_read_aggregated_cmd_halfPipe_payload_fragment_context;
  reg                 interconnect_read_aggregated_cmd_rValid;
  wire                interconnect_read_aggregated_cmd_halfPipe_fire;
  reg                 interconnect_read_aggregated_cmd_rData_last;
  reg        [0:0]    interconnect_read_aggregated_cmd_rData_fragment_source;
  reg        [0:0]    interconnect_read_aggregated_cmd_rData_fragment_opcode;
  reg        [31:0]   interconnect_read_aggregated_cmd_rData_fragment_address;
  reg        [12:0]   interconnect_read_aggregated_cmd_rData_fragment_length;
  reg        [24:0]   interconnect_read_aggregated_cmd_rData_fragment_context;
  wire                readLogic_resized_rsp_combStage_valid;
  wire                readLogic_resized_rsp_combStage_ready;
  wire                readLogic_resized_rsp_combStage_payload_last;
  wire       [0:0]    readLogic_resized_rsp_combStage_payload_fragment_source;
  wire       [0:0]    readLogic_resized_rsp_combStage_payload_fragment_opcode;
  wire       [255:0]  readLogic_resized_rsp_combStage_payload_fragment_data;
  wire       [24:0]   readLogic_resized_rsp_combStage_payload_fragment_context;
  wire                readLogic_adapter_ar_valid;
  wire                readLogic_adapter_ar_ready;
  wire       [31:0]   readLogic_adapter_ar_payload_addr;
  wire       [3:0]    readLogic_adapter_ar_payload_region;
  wire       [7:0]    readLogic_adapter_ar_payload_len;
  wire       [2:0]    readLogic_adapter_ar_payload_size;
  wire       [1:0]    readLogic_adapter_ar_payload_burst;
  wire       [0:0]    readLogic_adapter_ar_payload_lock;
  wire       [3:0]    readLogic_adapter_ar_payload_cache;
  wire       [3:0]    readLogic_adapter_ar_payload_qos;
  wire       [2:0]    readLogic_adapter_ar_payload_prot;
  wire                readLogic_adapter_r_valid;
  wire                readLogic_adapter_r_ready;
  wire       [255:0]  readLogic_adapter_r_payload_data;
  wire       [1:0]    readLogic_adapter_r_payload_resp;
  wire                readLogic_adapter_r_payload_last;
  wire       [3:0]    _zz_readLogic_adapter_ar_payload_region;
  wire                readLogic_adapter_ar_halfPipe_valid;
  wire                readLogic_adapter_ar_halfPipe_ready;
  wire       [31:0]   readLogic_adapter_ar_halfPipe_payload_addr;
  wire       [3:0]    readLogic_adapter_ar_halfPipe_payload_region;
  wire       [7:0]    readLogic_adapter_ar_halfPipe_payload_len;
  wire       [2:0]    readLogic_adapter_ar_halfPipe_payload_size;
  wire       [1:0]    readLogic_adapter_ar_halfPipe_payload_burst;
  wire       [0:0]    readLogic_adapter_ar_halfPipe_payload_lock;
  wire       [3:0]    readLogic_adapter_ar_halfPipe_payload_cache;
  wire       [3:0]    readLogic_adapter_ar_halfPipe_payload_qos;
  wire       [2:0]    readLogic_adapter_ar_halfPipe_payload_prot;
  reg                 readLogic_adapter_ar_rValid;
  wire                readLogic_adapter_ar_halfPipe_fire;
  reg        [31:0]   readLogic_adapter_ar_rData_addr;
  reg        [3:0]    readLogic_adapter_ar_rData_region;
  reg        [7:0]    readLogic_adapter_ar_rData_len;
  reg        [2:0]    readLogic_adapter_ar_rData_size;
  reg        [1:0]    readLogic_adapter_ar_rData_burst;
  reg        [0:0]    readLogic_adapter_ar_rData_lock;
  reg        [3:0]    readLogic_adapter_ar_rData_cache;
  reg        [3:0]    readLogic_adapter_ar_rData_qos;
  reg        [2:0]    readLogic_adapter_ar_rData_prot;
  wire                read_r_s2mPipe_valid;
  reg                 read_r_s2mPipe_ready;
  wire       [255:0]  read_r_s2mPipe_payload_data;
  wire       [1:0]    read_r_s2mPipe_payload_resp;
  wire                read_r_s2mPipe_payload_last;
  reg                 read_r_rValidN;
  reg        [255:0]  read_r_rData_data;
  reg        [1:0]    read_r_rData_resp;
  reg                 read_r_rData_last;
  wire                readLogic_beforeQueue_valid;
  wire                readLogic_beforeQueue_ready;
  wire       [255:0]  readLogic_beforeQueue_payload_data;
  wire       [1:0]    readLogic_beforeQueue_payload_resp;
  wire                readLogic_beforeQueue_payload_last;
  reg                 read_r_s2mPipe_rValid;
  reg        [255:0]  read_r_s2mPipe_rData_data;
  reg        [1:0]    read_r_s2mPipe_rData_resp;
  reg                 read_r_s2mPipe_rData_last;
  wire                when_Stream_l375_1;
  wire                writeLogic_resized_cmd_valid;
  wire                writeLogic_resized_cmd_ready;
  wire                writeLogic_resized_cmd_payload_last;
  wire       [0:0]    writeLogic_resized_cmd_payload_fragment_source;
  wire       [0:0]    writeLogic_resized_cmd_payload_fragment_opcode;
  wire       [31:0]   writeLogic_resized_cmd_payload_fragment_address;
  wire       [12:0]   writeLogic_resized_cmd_payload_fragment_length;
  wire       [255:0]  writeLogic_resized_cmd_payload_fragment_data;
  wire       [31:0]   writeLogic_resized_cmd_payload_fragment_mask;
  wire       [14:0]   writeLogic_resized_cmd_payload_fragment_context;
  wire                writeLogic_resized_rsp_valid;
  wire                writeLogic_resized_rsp_ready;
  wire                writeLogic_resized_rsp_payload_last;
  wire       [0:0]    writeLogic_resized_rsp_payload_fragment_source;
  wire       [0:0]    writeLogic_resized_rsp_payload_fragment_opcode;
  wire       [14:0]   writeLogic_resized_rsp_payload_fragment_context;
  wire                interconnect_write_aggregated_cmd_m2sPipe_valid;
  wire                interconnect_write_aggregated_cmd_m2sPipe_ready;
  wire                interconnect_write_aggregated_cmd_m2sPipe_payload_last;
  wire       [0:0]    interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_source;
  wire       [0:0]    interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_address;
  wire       [12:0]   interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_length;
  wire       [255:0]  interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_data;
  wire       [31:0]   interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_mask;
  wire       [14:0]   interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_context;
  reg                 interconnect_write_aggregated_cmd_rValid;
  reg                 interconnect_write_aggregated_cmd_rData_last;
  reg        [0:0]    interconnect_write_aggregated_cmd_rData_fragment_source;
  reg        [0:0]    interconnect_write_aggregated_cmd_rData_fragment_opcode;
  reg        [31:0]   interconnect_write_aggregated_cmd_rData_fragment_address;
  reg        [12:0]   interconnect_write_aggregated_cmd_rData_fragment_length;
  reg        [255:0]  interconnect_write_aggregated_cmd_rData_fragment_data;
  reg        [31:0]   interconnect_write_aggregated_cmd_rData_fragment_mask;
  reg        [14:0]   interconnect_write_aggregated_cmd_rData_fragment_context;
  wire                when_Stream_l375_2;
  wire                writeLogic_resized_rsp_combStage_valid;
  wire                writeLogic_resized_rsp_combStage_ready;
  wire                writeLogic_resized_rsp_combStage_payload_last;
  wire       [0:0]    writeLogic_resized_rsp_combStage_payload_fragment_source;
  wire       [0:0]    writeLogic_resized_rsp_combStage_payload_fragment_opcode;
  wire       [14:0]   writeLogic_resized_rsp_combStage_payload_fragment_context;
  wire                writeLogic_adapter_aw_valid;
  wire                writeLogic_adapter_aw_ready;
  wire       [31:0]   writeLogic_adapter_aw_payload_addr;
  wire       [3:0]    writeLogic_adapter_aw_payload_region;
  wire       [7:0]    writeLogic_adapter_aw_payload_len;
  wire       [2:0]    writeLogic_adapter_aw_payload_size;
  wire       [1:0]    writeLogic_adapter_aw_payload_burst;
  wire       [0:0]    writeLogic_adapter_aw_payload_lock;
  wire       [3:0]    writeLogic_adapter_aw_payload_cache;
  wire       [3:0]    writeLogic_adapter_aw_payload_qos;
  wire       [2:0]    writeLogic_adapter_aw_payload_prot;
  wire                writeLogic_adapter_w_valid;
  wire                writeLogic_adapter_w_ready;
  wire       [255:0]  writeLogic_adapter_w_payload_data;
  wire       [31:0]   writeLogic_adapter_w_payload_strb;
  wire                writeLogic_adapter_w_payload_last;
  wire                writeLogic_adapter_b_valid;
  wire                writeLogic_adapter_b_ready;
  wire       [1:0]    writeLogic_adapter_b_payload_resp;
  wire       [3:0]    _zz_writeLogic_adapter_aw_payload_region;
  wire                writeLogic_adapter_aw_halfPipe_valid;
  wire                writeLogic_adapter_aw_halfPipe_ready;
  wire       [31:0]   writeLogic_adapter_aw_halfPipe_payload_addr;
  wire       [3:0]    writeLogic_adapter_aw_halfPipe_payload_region;
  wire       [7:0]    writeLogic_adapter_aw_halfPipe_payload_len;
  wire       [2:0]    writeLogic_adapter_aw_halfPipe_payload_size;
  wire       [1:0]    writeLogic_adapter_aw_halfPipe_payload_burst;
  wire       [0:0]    writeLogic_adapter_aw_halfPipe_payload_lock;
  wire       [3:0]    writeLogic_adapter_aw_halfPipe_payload_cache;
  wire       [3:0]    writeLogic_adapter_aw_halfPipe_payload_qos;
  wire       [2:0]    writeLogic_adapter_aw_halfPipe_payload_prot;
  reg                 writeLogic_adapter_aw_rValid;
  wire                writeLogic_adapter_aw_halfPipe_fire;
  reg        [31:0]   writeLogic_adapter_aw_rData_addr;
  reg        [3:0]    writeLogic_adapter_aw_rData_region;
  reg        [7:0]    writeLogic_adapter_aw_rData_len;
  reg        [2:0]    writeLogic_adapter_aw_rData_size;
  reg        [1:0]    writeLogic_adapter_aw_rData_burst;
  reg        [0:0]    writeLogic_adapter_aw_rData_lock;
  reg        [3:0]    writeLogic_adapter_aw_rData_cache;
  reg        [3:0]    writeLogic_adapter_aw_rData_qos;
  reg        [2:0]    writeLogic_adapter_aw_rData_prot;
  wire                writeLogic_adapter_w_s2mPipe_valid;
  reg                 writeLogic_adapter_w_s2mPipe_ready;
  wire       [255:0]  writeLogic_adapter_w_s2mPipe_payload_data;
  wire       [31:0]   writeLogic_adapter_w_s2mPipe_payload_strb;
  wire                writeLogic_adapter_w_s2mPipe_payload_last;
  reg                 writeLogic_adapter_w_rValidN;
  reg        [255:0]  writeLogic_adapter_w_rData_data;
  reg        [31:0]   writeLogic_adapter_w_rData_strb;
  reg                 writeLogic_adapter_w_rData_last;
  wire                writeLogic_adapter_w_s2mPipe_m2sPipe_valid;
  wire                writeLogic_adapter_w_s2mPipe_m2sPipe_ready;
  wire       [255:0]  writeLogic_adapter_w_s2mPipe_m2sPipe_payload_data;
  wire       [31:0]   writeLogic_adapter_w_s2mPipe_m2sPipe_payload_strb;
  wire                writeLogic_adapter_w_s2mPipe_m2sPipe_payload_last;
  reg                 writeLogic_adapter_w_s2mPipe_rValid;
  reg        [255:0]  writeLogic_adapter_w_s2mPipe_rData_data;
  reg        [31:0]   writeLogic_adapter_w_s2mPipe_rData_strb;
  reg                 writeLogic_adapter_w_s2mPipe_rData_last;
  wire                when_Stream_l375_3;
  wire                write_b_halfPipe_valid;
  wire                write_b_halfPipe_ready;
  wire       [1:0]    write_b_halfPipe_payload_resp;
  reg                 write_b_rValid;
  wire                write_b_halfPipe_fire;
  reg        [1:0]    write_b_rData_resp;
  wire                io_pop_s2mPipe_valid;
  reg                 io_pop_s2mPipe_ready;
  wire       [127:0]  io_pop_s2mPipe_payload_data;
  wire       [15:0]   io_pop_s2mPipe_payload_mask;
  wire       [3:0]    io_pop_s2mPipe_payload_sink;
  wire                io_pop_s2mPipe_payload_last;
  reg                 io_pop_rValidN;
  reg        [127:0]  io_pop_rData_data;
  reg        [15:0]   io_pop_rData_mask;
  reg        [3:0]    io_pop_rData_sink;
  reg                 io_pop_rData_last;
  wire                io_pop_s2mPipe_m2sPipe_valid;
  wire                io_pop_s2mPipe_m2sPipe_ready;
  wire       [127:0]  io_pop_s2mPipe_m2sPipe_payload_data;
  wire       [15:0]   io_pop_s2mPipe_m2sPipe_payload_mask;
  wire       [3:0]    io_pop_s2mPipe_m2sPipe_payload_sink;
  wire                io_pop_s2mPipe_m2sPipe_payload_last;
  reg                 io_pop_s2mPipe_rValid;
  reg        [127:0]  io_pop_s2mPipe_rData_data;
  reg        [15:0]   io_pop_s2mPipe_rData_mask;
  reg        [3:0]    io_pop_s2mPipe_rData_sink;
  reg                 io_pop_s2mPipe_rData_last;
  wire                when_Stream_l375_4;
  wire                io_pop_s2mPipe_valid_1;
  reg                 io_pop_s2mPipe_ready_1;
  wire       [127:0]  io_pop_s2mPipe_payload_data_1;
  wire       [15:0]   io_pop_s2mPipe_payload_mask_1;
  wire       [3:0]    io_pop_s2mPipe_payload_sink_1;
  wire                io_pop_s2mPipe_payload_last_1;
  reg                 io_pop_rValidN_1;
  reg        [127:0]  io_pop_rData_data_1;
  reg        [15:0]   io_pop_rData_mask_1;
  reg        [3:0]    io_pop_rData_sink_1;
  reg                 io_pop_rData_last_1;
  wire                io_pop_s2mPipe_m2sPipe_valid_1;
  wire                io_pop_s2mPipe_m2sPipe_ready_1;
  wire       [127:0]  io_pop_s2mPipe_m2sPipe_payload_data_1;
  wire       [15:0]   io_pop_s2mPipe_m2sPipe_payload_mask_1;
  wire       [3:0]    io_pop_s2mPipe_m2sPipe_payload_sink_1;
  wire                io_pop_s2mPipe_m2sPipe_payload_last_1;
  reg                 io_pop_s2mPipe_rValid_1;
  reg        [127:0]  io_pop_s2mPipe_rData_data_1;
  reg        [15:0]   io_pop_s2mPipe_rData_mask_1;
  reg        [3:0]    io_pop_s2mPipe_rData_sink_1;
  reg                 io_pop_s2mPipe_rData_last_1;
  wire                when_Stream_l375_5;
  wire                io_outputs_0_s2mPipe_valid;
  reg                 io_outputs_0_s2mPipe_ready;
  wire       [127:0]  io_outputs_0_s2mPipe_payload_data;
  wire       [15:0]   io_outputs_0_s2mPipe_payload_mask;
  wire       [3:0]    io_outputs_0_s2mPipe_payload_sink;
  wire                io_outputs_0_s2mPipe_payload_last;
  reg                 io_outputs_0_rValidN;
  reg        [127:0]  io_outputs_0_rData_data;
  reg        [15:0]   io_outputs_0_rData_mask;
  reg        [3:0]    io_outputs_0_rData_sink;
  reg                 io_outputs_0_rData_last;
  wire                outputsAdapter_0_ptr_valid;
  wire                outputsAdapter_0_ptr_ready;
  wire       [127:0]  outputsAdapter_0_ptr_payload_data;
  wire       [15:0]   outputsAdapter_0_ptr_payload_mask;
  wire       [3:0]    outputsAdapter_0_ptr_payload_sink;
  wire                outputsAdapter_0_ptr_payload_last;
  reg                 io_outputs_0_s2mPipe_rValid;
  reg        [127:0]  io_outputs_0_s2mPipe_rData_data;
  reg        [15:0]   io_outputs_0_s2mPipe_rData_mask;
  reg        [3:0]    io_outputs_0_s2mPipe_rData_sink;
  reg                 io_outputs_0_s2mPipe_rData_last;
  wire                when_Stream_l375_6;
  wire                io_outputs_1_s2mPipe_valid;
  reg                 io_outputs_1_s2mPipe_ready;
  wire       [127:0]  io_outputs_1_s2mPipe_payload_data;
  wire       [15:0]   io_outputs_1_s2mPipe_payload_mask;
  wire       [3:0]    io_outputs_1_s2mPipe_payload_sink;
  wire                io_outputs_1_s2mPipe_payload_last;
  reg                 io_outputs_1_rValidN;
  reg        [127:0]  io_outputs_1_rData_data;
  reg        [15:0]   io_outputs_1_rData_mask;
  reg        [3:0]    io_outputs_1_rData_sink;
  reg                 io_outputs_1_rData_last;
  wire                outputsAdapter_1_ptr_valid;
  wire                outputsAdapter_1_ptr_ready;
  wire       [127:0]  outputsAdapter_1_ptr_payload_data;
  wire       [15:0]   outputsAdapter_1_ptr_payload_mask;
  wire       [3:0]    outputsAdapter_1_ptr_payload_sink;
  wire                outputsAdapter_1_ptr_payload_last;
  reg                 io_outputs_1_s2mPipe_rValid;
  reg        [127:0]  io_outputs_1_s2mPipe_rData_data;
  reg        [15:0]   io_outputs_1_s2mPipe_rData_mask;
  reg        [3:0]    io_outputs_1_s2mPipe_rData_sink;
  reg                 io_outputs_1_s2mPipe_rData_last;
  wire                when_Stream_l375_7;
  wire                interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  wire       [0:0]    interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [31:0]   interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [12:0]   interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [24:0]   interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [255:0]  interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [24:0]   interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  wire       [0:0]    interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [31:0]   interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [12:0]   interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [255:0]  interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [31:0]   interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [14:0]   interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [14:0]   interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;

  EfxDMA_Core core (
    .io_read_cmd_valid                     (core_io_read_cmd_valid                                                                                 ), //o
    .io_read_cmd_ready                     (interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready                          ), //i
    .io_read_cmd_payload_last              (core_io_read_cmd_payload_last                                                                          ), //o
    .io_read_cmd_payload_fragment_source   (core_io_read_cmd_payload_fragment_source                                                               ), //o
    .io_read_cmd_payload_fragment_opcode   (core_io_read_cmd_payload_fragment_opcode                                                               ), //o
    .io_read_cmd_payload_fragment_address  (core_io_read_cmd_payload_fragment_address[31:0]                                                        ), //o
    .io_read_cmd_payload_fragment_length   (core_io_read_cmd_payload_fragment_length[12:0]                                                         ), //o
    .io_read_cmd_payload_fragment_context  (core_io_read_cmd_payload_fragment_context[24:0]                                                        ), //o
    .io_read_rsp_valid                     (interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid                          ), //i
    .io_read_rsp_ready                     (core_io_read_rsp_ready                                                                                 ), //o
    .io_read_rsp_payload_last              (interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last                   ), //i
    .io_read_rsp_payload_fragment_source   (interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source        ), //i
    .io_read_rsp_payload_fragment_opcode   (interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode        ), //i
    .io_read_rsp_payload_fragment_data     (interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data[255:0]   ), //i
    .io_read_rsp_payload_fragment_context  (interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context[24:0] ), //i
    .io_write_cmd_valid                    (core_io_write_cmd_valid                                                                                ), //o
    .io_write_cmd_ready                    (io_write_cmd_rValidN                                                                                   ), //i
    .io_write_cmd_payload_last             (core_io_write_cmd_payload_last                                                                         ), //o
    .io_write_cmd_payload_fragment_source  (core_io_write_cmd_payload_fragment_source                                                              ), //o
    .io_write_cmd_payload_fragment_opcode  (core_io_write_cmd_payload_fragment_opcode                                                              ), //o
    .io_write_cmd_payload_fragment_address (core_io_write_cmd_payload_fragment_address[31:0]                                                       ), //o
    .io_write_cmd_payload_fragment_length  (core_io_write_cmd_payload_fragment_length[12:0]                                                        ), //o
    .io_write_cmd_payload_fragment_data    (core_io_write_cmd_payload_fragment_data[255:0]                                                         ), //o
    .io_write_cmd_payload_fragment_mask    (core_io_write_cmd_payload_fragment_mask[31:0]                                                          ), //o
    .io_write_cmd_payload_fragment_context (core_io_write_cmd_payload_fragment_context[14:0]                                                       ), //o
    .io_write_rsp_valid                    (interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid                         ), //i
    .io_write_rsp_ready                    (core_io_write_rsp_ready                                                                                ), //o
    .io_write_rsp_payload_last             (interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last                  ), //i
    .io_write_rsp_payload_fragment_source  (interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source       ), //i
    .io_write_rsp_payload_fragment_opcode  (interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode       ), //i
    .io_write_rsp_payload_fragment_context (interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context[14:0]), //i
    .io_outputs_0_valid                    (core_io_outputs_0_valid                                                                                ), //o
    .io_outputs_0_ready                    (io_outputs_0_rValidN                                                                                   ), //i
    .io_outputs_0_payload_data             (core_io_outputs_0_payload_data[127:0]                                                                  ), //o
    .io_outputs_0_payload_mask             (core_io_outputs_0_payload_mask[15:0]                                                                   ), //o
    .io_outputs_0_payload_sink             (core_io_outputs_0_payload_sink[3:0]                                                                    ), //o
    .io_outputs_0_payload_last             (core_io_outputs_0_payload_last                                                                         ), //o
    .io_outputs_1_valid                    (core_io_outputs_1_valid                                                                                ), //o
    .io_outputs_1_ready                    (io_outputs_1_rValidN                                                                                   ), //i
    .io_outputs_1_payload_data             (core_io_outputs_1_payload_data[127:0]                                                                  ), //o
    .io_outputs_1_payload_mask             (core_io_outputs_1_payload_mask[15:0]                                                                   ), //o
    .io_outputs_1_payload_sink             (core_io_outputs_1_payload_sink[3:0]                                                                    ), //o
    .io_outputs_1_payload_last             (core_io_outputs_1_payload_last                                                                         ), //o
    .io_inputs_0_valid                     (io_pop_s2mPipe_m2sPipe_valid                                                                           ), //i
    .io_inputs_0_ready                     (core_io_inputs_0_ready                                                                                 ), //o
    .io_inputs_0_payload_data              (io_pop_s2mPipe_m2sPipe_payload_data[127:0]                                                             ), //i
    .io_inputs_0_payload_mask              (io_pop_s2mPipe_m2sPipe_payload_mask[15:0]                                                              ), //i
    .io_inputs_0_payload_sink              (io_pop_s2mPipe_m2sPipe_payload_sink[3:0]                                                               ), //i
    .io_inputs_0_payload_last              (io_pop_s2mPipe_m2sPipe_payload_last                                                                    ), //i
    .io_inputs_1_valid                     (io_pop_s2mPipe_m2sPipe_valid_1                                                                         ), //i
    .io_inputs_1_ready                     (core_io_inputs_1_ready                                                                                 ), //o
    .io_inputs_1_payload_data              (io_pop_s2mPipe_m2sPipe_payload_data_1[127:0]                                                           ), //i
    .io_inputs_1_payload_mask              (io_pop_s2mPipe_m2sPipe_payload_mask_1[15:0]                                                            ), //i
    .io_inputs_1_payload_sink              (io_pop_s2mPipe_m2sPipe_payload_sink_1[3:0]                                                             ), //i
    .io_inputs_1_payload_last              (io_pop_s2mPipe_m2sPipe_payload_last_1                                                                  ), //i
    .io_interrupts                         (core_io_interrupts[3:0]                                                                                ), //o
    .io_ctrl_PADDR                         (withCtrlCc_apbCc_io_output_PADDR[13:0]                                                                 ), //i
    .io_ctrl_PSEL                          (withCtrlCc_apbCc_io_output_PSEL                                                                        ), //i
    .io_ctrl_PENABLE                       (withCtrlCc_apbCc_io_output_PENABLE                                                                     ), //i
    .io_ctrl_PREADY                        (core_io_ctrl_PREADY                                                                                    ), //o
    .io_ctrl_PWRITE                        (withCtrlCc_apbCc_io_output_PWRITE                                                                      ), //i
    .io_ctrl_PWDATA                        (withCtrlCc_apbCc_io_output_PWDATA[31:0]                                                                ), //i
    .io_ctrl_PRDATA                        (core_io_ctrl_PRDATA[31:0]                                                                              ), //o
    .io_ctrl_PSLVERROR                     (core_io_ctrl_PSLVERROR                                                                                 ), //o
    .clk                                   (clk                                                                                                    ), //i
    .reset                                 (reset                                                                                                  )  //i
  );
  EfxDMA_Apb3CC withCtrlCc_apbCc (
    .io_input_PADDR      (ctrl_PADDR[13:0]                       ), //i
    .io_input_PSEL       (ctrl_PSEL                              ), //i
    .io_input_PENABLE    (ctrl_PENABLE                           ), //i
    .io_input_PREADY     (withCtrlCc_apbCc_io_input_PREADY       ), //o
    .io_input_PWRITE     (ctrl_PWRITE                            ), //i
    .io_input_PWDATA     (ctrl_PWDATA[31:0]                      ), //i
    .io_input_PRDATA     (withCtrlCc_apbCc_io_input_PRDATA[31:0] ), //o
    .io_input_PSLVERROR  (withCtrlCc_apbCc_io_input_PSLVERROR    ), //o
    .io_output_PADDR     (withCtrlCc_apbCc_io_output_PADDR[13:0] ), //o
    .io_output_PSEL      (withCtrlCc_apbCc_io_output_PSEL        ), //o
    .io_output_PENABLE   (withCtrlCc_apbCc_io_output_PENABLE     ), //o
    .io_output_PREADY    (core_io_ctrl_PREADY                    ), //i
    .io_output_PWRITE    (withCtrlCc_apbCc_io_output_PWRITE      ), //o
    .io_output_PWDATA    (withCtrlCc_apbCc_io_output_PWDATA[31:0]), //o
    .io_output_PRDATA    (core_io_ctrl_PRDATA[31:0]              ), //i
    .io_output_PSLVERROR (core_io_ctrl_PSLVERROR                 ), //i
    .ctrl_clk            (ctrl_clk                               ), //i
    .ctrl_reset          (ctrl_reset                             ), //i
    .clk                 (clk                                    ), //i
    .reset               (reset                                  )  //i
  );
  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_10 io_interrupts_buffercc (
    .io_dataIn  (core_io_interrupts[3:0]               ), //i
    .io_dataOut (io_interrupts_buffercc_io_dataOut[3:0]), //o
    .ctrl_clk   (ctrl_clk                              ), //i
    .ctrl_reset (ctrl_reset                            )  //i
  );
  EfxDMA_BmbSourceRemover readLogic_sourceRemover (
    .io_input_cmd_valid                     (readLogic_resized_cmd_valid                                         ), //i
    .io_input_cmd_ready                     (readLogic_sourceRemover_io_input_cmd_ready                          ), //o
    .io_input_cmd_payload_last              (readLogic_resized_cmd_payload_last                                  ), //i
    .io_input_cmd_payload_fragment_source   (readLogic_resized_cmd_payload_fragment_source                       ), //i
    .io_input_cmd_payload_fragment_opcode   (readLogic_resized_cmd_payload_fragment_opcode                       ), //i
    .io_input_cmd_payload_fragment_address  (readLogic_resized_cmd_payload_fragment_address[31:0]                ), //i
    .io_input_cmd_payload_fragment_length   (readLogic_resized_cmd_payload_fragment_length[12:0]                 ), //i
    .io_input_cmd_payload_fragment_context  (readLogic_resized_cmd_payload_fragment_context[24:0]                ), //i
    .io_input_rsp_valid                     (readLogic_sourceRemover_io_input_rsp_valid                          ), //o
    .io_input_rsp_ready                     (readLogic_resized_rsp_ready                                         ), //i
    .io_input_rsp_payload_last              (readLogic_sourceRemover_io_input_rsp_payload_last                   ), //o
    .io_input_rsp_payload_fragment_source   (readLogic_sourceRemover_io_input_rsp_payload_fragment_source        ), //o
    .io_input_rsp_payload_fragment_opcode   (readLogic_sourceRemover_io_input_rsp_payload_fragment_opcode        ), //o
    .io_input_rsp_payload_fragment_data     (readLogic_sourceRemover_io_input_rsp_payload_fragment_data[255:0]   ), //o
    .io_input_rsp_payload_fragment_context  (readLogic_sourceRemover_io_input_rsp_payload_fragment_context[24:0] ), //o
    .io_output_cmd_valid                    (readLogic_sourceRemover_io_output_cmd_valid                         ), //o
    .io_output_cmd_ready                    (readLogic_bridge_io_input_cmd_ready                                 ), //i
    .io_output_cmd_payload_last             (readLogic_sourceRemover_io_output_cmd_payload_last                  ), //o
    .io_output_cmd_payload_fragment_opcode  (readLogic_sourceRemover_io_output_cmd_payload_fragment_opcode       ), //o
    .io_output_cmd_payload_fragment_address (readLogic_sourceRemover_io_output_cmd_payload_fragment_address[31:0]), //o
    .io_output_cmd_payload_fragment_length  (readLogic_sourceRemover_io_output_cmd_payload_fragment_length[12:0] ), //o
    .io_output_cmd_payload_fragment_context (readLogic_sourceRemover_io_output_cmd_payload_fragment_context[25:0]), //o
    .io_output_rsp_valid                    (readLogic_bridge_io_input_rsp_valid                                 ), //i
    .io_output_rsp_ready                    (readLogic_sourceRemover_io_output_rsp_ready                         ), //o
    .io_output_rsp_payload_last             (readLogic_bridge_io_input_rsp_payload_last                          ), //i
    .io_output_rsp_payload_fragment_opcode  (readLogic_bridge_io_input_rsp_payload_fragment_opcode               ), //i
    .io_output_rsp_payload_fragment_data    (readLogic_bridge_io_input_rsp_payload_fragment_data[255:0]          ), //i
    .io_output_rsp_payload_fragment_context (readLogic_bridge_io_input_rsp_payload_fragment_context[25:0]        )  //i
  );
  EfxDMA_BmbToAxi4ReadOnlyBridge readLogic_bridge (
    .io_input_cmd_valid                    (readLogic_sourceRemover_io_output_cmd_valid                         ), //i
    .io_input_cmd_ready                    (readLogic_bridge_io_input_cmd_ready                                 ), //o
    .io_input_cmd_payload_last             (readLogic_sourceRemover_io_output_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_opcode  (readLogic_sourceRemover_io_output_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (readLogic_sourceRemover_io_output_cmd_payload_fragment_address[31:0]), //i
    .io_input_cmd_payload_fragment_length  (readLogic_sourceRemover_io_output_cmd_payload_fragment_length[12:0] ), //i
    .io_input_cmd_payload_fragment_context (readLogic_sourceRemover_io_output_cmd_payload_fragment_context[25:0]), //i
    .io_input_rsp_valid                    (readLogic_bridge_io_input_rsp_valid                                 ), //o
    .io_input_rsp_ready                    (readLogic_sourceRemover_io_output_rsp_ready                         ), //i
    .io_input_rsp_payload_last             (readLogic_bridge_io_input_rsp_payload_last                          ), //o
    .io_input_rsp_payload_fragment_opcode  (readLogic_bridge_io_input_rsp_payload_fragment_opcode               ), //o
    .io_input_rsp_payload_fragment_data    (readLogic_bridge_io_input_rsp_payload_fragment_data[255:0]          ), //o
    .io_input_rsp_payload_fragment_context (readLogic_bridge_io_input_rsp_payload_fragment_context[25:0]        ), //o
    .io_output_ar_valid                    (readLogic_bridge_io_output_ar_valid                                 ), //o
    .io_output_ar_ready                    (readLogic_adapter_ar_ready                                          ), //i
    .io_output_ar_payload_addr             (readLogic_bridge_io_output_ar_payload_addr[31:0]                    ), //o
    .io_output_ar_payload_len              (readLogic_bridge_io_output_ar_payload_len[7:0]                      ), //o
    .io_output_ar_payload_size             (readLogic_bridge_io_output_ar_payload_size[2:0]                     ), //o
    .io_output_ar_payload_cache            (readLogic_bridge_io_output_ar_payload_cache[3:0]                    ), //o
    .io_output_ar_payload_prot             (readLogic_bridge_io_output_ar_payload_prot[2:0]                     ), //o
    .io_output_r_valid                     (readLogic_adapter_r_valid                                           ), //i
    .io_output_r_ready                     (readLogic_bridge_io_output_r_ready                                  ), //o
    .io_output_r_payload_data              (readLogic_adapter_r_payload_data[255:0]                             ), //i
    .io_output_r_payload_resp              (readLogic_adapter_r_payload_resp[1:0]                               ), //i
    .io_output_r_payload_last              (readLogic_adapter_r_payload_last                                    ), //i
    .clk                                   (clk                                                                 ), //i
    .reset                                 (reset                                                               )  //i
  );
  EfxDMA_BmbSourceRemover_1 writeLogic_sourceRemover (
    .io_input_cmd_valid                     (writeLogic_resized_cmd_valid                                         ), //i
    .io_input_cmd_ready                     (writeLogic_sourceRemover_io_input_cmd_ready                          ), //o
    .io_input_cmd_payload_last              (writeLogic_resized_cmd_payload_last                                  ), //i
    .io_input_cmd_payload_fragment_source   (writeLogic_resized_cmd_payload_fragment_source                       ), //i
    .io_input_cmd_payload_fragment_opcode   (writeLogic_resized_cmd_payload_fragment_opcode                       ), //i
    .io_input_cmd_payload_fragment_address  (writeLogic_resized_cmd_payload_fragment_address[31:0]                ), //i
    .io_input_cmd_payload_fragment_length   (writeLogic_resized_cmd_payload_fragment_length[12:0]                 ), //i
    .io_input_cmd_payload_fragment_data     (writeLogic_resized_cmd_payload_fragment_data[255:0]                  ), //i
    .io_input_cmd_payload_fragment_mask     (writeLogic_resized_cmd_payload_fragment_mask[31:0]                   ), //i
    .io_input_cmd_payload_fragment_context  (writeLogic_resized_cmd_payload_fragment_context[14:0]                ), //i
    .io_input_rsp_valid                     (writeLogic_sourceRemover_io_input_rsp_valid                          ), //o
    .io_input_rsp_ready                     (writeLogic_resized_rsp_ready                                         ), //i
    .io_input_rsp_payload_last              (writeLogic_sourceRemover_io_input_rsp_payload_last                   ), //o
    .io_input_rsp_payload_fragment_source   (writeLogic_sourceRemover_io_input_rsp_payload_fragment_source        ), //o
    .io_input_rsp_payload_fragment_opcode   (writeLogic_sourceRemover_io_input_rsp_payload_fragment_opcode        ), //o
    .io_input_rsp_payload_fragment_context  (writeLogic_sourceRemover_io_input_rsp_payload_fragment_context[14:0] ), //o
    .io_output_cmd_valid                    (writeLogic_sourceRemover_io_output_cmd_valid                         ), //o
    .io_output_cmd_ready                    (writeLogic_bridge_io_input_cmd_ready                                 ), //i
    .io_output_cmd_payload_last             (writeLogic_sourceRemover_io_output_cmd_payload_last                  ), //o
    .io_output_cmd_payload_fragment_opcode  (writeLogic_sourceRemover_io_output_cmd_payload_fragment_opcode       ), //o
    .io_output_cmd_payload_fragment_address (writeLogic_sourceRemover_io_output_cmd_payload_fragment_address[31:0]), //o
    .io_output_cmd_payload_fragment_length  (writeLogic_sourceRemover_io_output_cmd_payload_fragment_length[12:0] ), //o
    .io_output_cmd_payload_fragment_data    (writeLogic_sourceRemover_io_output_cmd_payload_fragment_data[255:0]  ), //o
    .io_output_cmd_payload_fragment_mask    (writeLogic_sourceRemover_io_output_cmd_payload_fragment_mask[31:0]   ), //o
    .io_output_cmd_payload_fragment_context (writeLogic_sourceRemover_io_output_cmd_payload_fragment_context[15:0]), //o
    .io_output_rsp_valid                    (writeLogic_bridge_io_input_rsp_valid                                 ), //i
    .io_output_rsp_ready                    (writeLogic_sourceRemover_io_output_rsp_ready                         ), //o
    .io_output_rsp_payload_last             (writeLogic_bridge_io_input_rsp_payload_last                          ), //i
    .io_output_rsp_payload_fragment_opcode  (writeLogic_bridge_io_input_rsp_payload_fragment_opcode               ), //i
    .io_output_rsp_payload_fragment_context (writeLogic_bridge_io_input_rsp_payload_fragment_context[15:0]        )  //i
  );
  EfxDMA_BmbToAxi4WriteOnlyBridge writeLogic_bridge (
    .io_input_cmd_valid                    (writeLogic_sourceRemover_io_output_cmd_valid                         ), //i
    .io_input_cmd_ready                    (writeLogic_bridge_io_input_cmd_ready                                 ), //o
    .io_input_cmd_payload_last             (writeLogic_sourceRemover_io_output_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_opcode  (writeLogic_sourceRemover_io_output_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (writeLogic_sourceRemover_io_output_cmd_payload_fragment_address[31:0]), //i
    .io_input_cmd_payload_fragment_length  (writeLogic_sourceRemover_io_output_cmd_payload_fragment_length[12:0] ), //i
    .io_input_cmd_payload_fragment_data    (writeLogic_sourceRemover_io_output_cmd_payload_fragment_data[255:0]  ), //i
    .io_input_cmd_payload_fragment_mask    (writeLogic_sourceRemover_io_output_cmd_payload_fragment_mask[31:0]   ), //i
    .io_input_cmd_payload_fragment_context (writeLogic_sourceRemover_io_output_cmd_payload_fragment_context[15:0]), //i
    .io_input_rsp_valid                    (writeLogic_bridge_io_input_rsp_valid                                 ), //o
    .io_input_rsp_ready                    (writeLogic_sourceRemover_io_output_rsp_ready                         ), //i
    .io_input_rsp_payload_last             (writeLogic_bridge_io_input_rsp_payload_last                          ), //o
    .io_input_rsp_payload_fragment_opcode  (writeLogic_bridge_io_input_rsp_payload_fragment_opcode               ), //o
    .io_input_rsp_payload_fragment_context (writeLogic_bridge_io_input_rsp_payload_fragment_context[15:0]        ), //o
    .io_output_aw_valid                    (writeLogic_bridge_io_output_aw_valid                                 ), //o
    .io_output_aw_ready                    (writeLogic_adapter_aw_ready                                          ), //i
    .io_output_aw_payload_addr             (writeLogic_bridge_io_output_aw_payload_addr[31:0]                    ), //o
    .io_output_aw_payload_len              (writeLogic_bridge_io_output_aw_payload_len[7:0]                      ), //o
    .io_output_aw_payload_size             (writeLogic_bridge_io_output_aw_payload_size[2:0]                     ), //o
    .io_output_aw_payload_cache            (writeLogic_bridge_io_output_aw_payload_cache[3:0]                    ), //o
    .io_output_aw_payload_prot             (writeLogic_bridge_io_output_aw_payload_prot[2:0]                     ), //o
    .io_output_w_valid                     (writeLogic_bridge_io_output_w_valid                                  ), //o
    .io_output_w_ready                     (writeLogic_adapter_w_ready                                           ), //i
    .io_output_w_payload_data              (writeLogic_bridge_io_output_w_payload_data[255:0]                    ), //o
    .io_output_w_payload_strb              (writeLogic_bridge_io_output_w_payload_strb[31:0]                     ), //o
    .io_output_w_payload_last              (writeLogic_bridge_io_output_w_payload_last                           ), //o
    .io_output_b_valid                     (writeLogic_adapter_b_valid                                           ), //i
    .io_output_b_ready                     (writeLogic_bridge_io_output_b_ready                                  ), //o
    .io_output_b_payload_resp              (writeLogic_adapter_b_payload_resp[1:0]                               ), //i
    .clk                                   (clk                                                                  ), //i
    .reset                                 (reset                                                                )  //i
  );
  EfxDMA_BsbUpSizerDense inputsAdapter_0_upsizer_logic (
    .io_input_valid         (dat0_i_tvalid                                              ), //i
    .io_input_ready         (inputsAdapter_0_upsizer_logic_io_input_ready               ), //o
    .io_input_payload_data  (dat0_i_tdata[63:0]                                         ), //i
    .io_input_payload_mask  (dat0_i_tkeep[7:0]                                          ), //i
    .io_input_payload_sink  (dat0_i_tdest[3:0]                                          ), //i
    .io_input_payload_last  (dat0_i_tlast                                               ), //i
    .io_output_valid        (inputsAdapter_0_upsizer_logic_io_output_valid              ), //o
    .io_output_ready        (inputsAdapter_0_crossclock_fifo_io_push_ready              ), //i
    .io_output_payload_data (inputsAdapter_0_upsizer_logic_io_output_payload_data[127:0]), //o
    .io_output_payload_mask (inputsAdapter_0_upsizer_logic_io_output_payload_mask[15:0] ), //o
    .io_output_payload_sink (inputsAdapter_0_upsizer_logic_io_output_payload_sink[3:0]  ), //o
    .io_output_payload_last (inputsAdapter_0_upsizer_logic_io_output_payload_last       ), //o
    .dat0_i_clk             (dat0_i_clk                                                 ), //i
    .dat0_i_reset           (dat0_i_reset                                               )  //i
  );
  EfxDMA_StreamFifoCC inputsAdapter_0_crossclock_fifo (
    .io_push_valid        (inputsAdapter_0_upsizer_logic_io_output_valid              ), //i
    .io_push_ready        (inputsAdapter_0_crossclock_fifo_io_push_ready              ), //o
    .io_push_payload_data (inputsAdapter_0_upsizer_logic_io_output_payload_data[127:0]), //i
    .io_push_payload_mask (inputsAdapter_0_upsizer_logic_io_output_payload_mask[15:0] ), //i
    .io_push_payload_sink (inputsAdapter_0_upsizer_logic_io_output_payload_sink[3:0]  ), //i
    .io_push_payload_last (inputsAdapter_0_upsizer_logic_io_output_payload_last       ), //i
    .io_pop_valid         (inputsAdapter_0_crossclock_fifo_io_pop_valid               ), //o
    .io_pop_ready         (io_pop_rValidN                                             ), //i
    .io_pop_payload_data  (inputsAdapter_0_crossclock_fifo_io_pop_payload_data[127:0] ), //o
    .io_pop_payload_mask  (inputsAdapter_0_crossclock_fifo_io_pop_payload_mask[15:0]  ), //o
    .io_pop_payload_sink  (inputsAdapter_0_crossclock_fifo_io_pop_payload_sink[3:0]   ), //o
    .io_pop_payload_last  (inputsAdapter_0_crossclock_fifo_io_pop_payload_last        ), //o
    .io_pushOccupancy     (inputsAdapter_0_crossclock_fifo_io_pushOccupancy[4:0]      ), //o
    .io_popOccupancy      (inputsAdapter_0_crossclock_fifo_io_popOccupancy[4:0]       ), //o
    .dat0_i_clk           (dat0_i_clk                                                 ), //i
    .dat0_i_reset         (dat0_i_reset                                               ), //i
    .clk                  (clk                                                        ), //i
    .reset                (reset                                                      )  //i
  );
  EfxDMA_BsbUpSizerDense_1 inputsAdapter_1_upsizer_logic (
    .io_input_valid         (dat2_i_tvalid                                              ), //i
    .io_input_ready         (inputsAdapter_1_upsizer_logic_io_input_ready               ), //o
    .io_input_payload_data  (dat2_i_tdata[31:0]                                         ), //i
    .io_input_payload_mask  (dat2_i_tkeep[3:0]                                          ), //i
    .io_input_payload_sink  (dat2_i_tdest[3:0]                                          ), //i
    .io_input_payload_last  (dat2_i_tlast                                               ), //i
    .io_output_valid        (inputsAdapter_1_upsizer_logic_io_output_valid              ), //o
    .io_output_ready        (inputsAdapter_1_crossclock_fifo_io_push_ready              ), //i
    .io_output_payload_data (inputsAdapter_1_upsizer_logic_io_output_payload_data[127:0]), //o
    .io_output_payload_mask (inputsAdapter_1_upsizer_logic_io_output_payload_mask[15:0] ), //o
    .io_output_payload_sink (inputsAdapter_1_upsizer_logic_io_output_payload_sink[3:0]  ), //o
    .io_output_payload_last (inputsAdapter_1_upsizer_logic_io_output_payload_last       ), //o
    .dat2_i_clk             (dat2_i_clk                                                 ), //i
    .dat2_i_reset           (dat2_i_reset                                               )  //i
  );
  EfxDMA_StreamFifoCC_1 inputsAdapter_1_crossclock_fifo (
    .io_push_valid        (inputsAdapter_1_upsizer_logic_io_output_valid              ), //i
    .io_push_ready        (inputsAdapter_1_crossclock_fifo_io_push_ready              ), //o
    .io_push_payload_data (inputsAdapter_1_upsizer_logic_io_output_payload_data[127:0]), //i
    .io_push_payload_mask (inputsAdapter_1_upsizer_logic_io_output_payload_mask[15:0] ), //i
    .io_push_payload_sink (inputsAdapter_1_upsizer_logic_io_output_payload_sink[3:0]  ), //i
    .io_push_payload_last (inputsAdapter_1_upsizer_logic_io_output_payload_last       ), //i
    .io_pop_valid         (inputsAdapter_1_crossclock_fifo_io_pop_valid               ), //o
    .io_pop_ready         (io_pop_rValidN_1                                           ), //i
    .io_pop_payload_data  (inputsAdapter_1_crossclock_fifo_io_pop_payload_data[127:0] ), //o
    .io_pop_payload_mask  (inputsAdapter_1_crossclock_fifo_io_pop_payload_mask[15:0]  ), //o
    .io_pop_payload_sink  (inputsAdapter_1_crossclock_fifo_io_pop_payload_sink[3:0]   ), //o
    .io_pop_payload_last  (inputsAdapter_1_crossclock_fifo_io_pop_payload_last        ), //o
    .io_pushOccupancy     (inputsAdapter_1_crossclock_fifo_io_pushOccupancy[4:0]      ), //o
    .io_popOccupancy      (inputsAdapter_1_crossclock_fifo_io_popOccupancy[4:0]       ), //o
    .dat2_i_clk           (dat2_i_clk                                                 ), //i
    .dat2_i_reset         (dat2_i_reset                                               ), //i
    .clk                  (clk                                                        ), //i
    .reset                (reset                                                      )  //i
  );
  EfxDMA_StreamFifoCC_2 outputsAdapter_0_crossclock_fifo (
    .io_push_valid        (outputsAdapter_0_ptr_valid                                 ), //i
    .io_push_ready        (outputsAdapter_0_crossclock_fifo_io_push_ready             ), //o
    .io_push_payload_data (outputsAdapter_0_ptr_payload_data[127:0]                   ), //i
    .io_push_payload_mask (outputsAdapter_0_ptr_payload_mask[15:0]                    ), //i
    .io_push_payload_sink (outputsAdapter_0_ptr_payload_sink[3:0]                     ), //i
    .io_push_payload_last (outputsAdapter_0_ptr_payload_last                          ), //i
    .io_pop_valid         (outputsAdapter_0_crossclock_fifo_io_pop_valid              ), //o
    .io_pop_ready         (outputsAdapter_0_sparseDownsizer_logic_io_input_ready      ), //i
    .io_pop_payload_data  (outputsAdapter_0_crossclock_fifo_io_pop_payload_data[127:0]), //o
    .io_pop_payload_mask  (outputsAdapter_0_crossclock_fifo_io_pop_payload_mask[15:0] ), //o
    .io_pop_payload_sink  (outputsAdapter_0_crossclock_fifo_io_pop_payload_sink[3:0]  ), //o
    .io_pop_payload_last  (outputsAdapter_0_crossclock_fifo_io_pop_payload_last       ), //o
    .io_pushOccupancy     (outputsAdapter_0_crossclock_fifo_io_pushOccupancy[4:0]     ), //o
    .io_popOccupancy      (outputsAdapter_0_crossclock_fifo_io_popOccupancy[4:0]      ), //o
    .clk                  (clk                                                        ), //i
    .reset                (reset                                                      ), //i
    .dat1_o_clk           (dat1_o_clk                                                 ), //i
    .dat1_o_reset         (dat1_o_reset                                               )  //i
  );
  EfxDMA_BsbDownSizerSparse outputsAdapter_0_sparseDownsizer_logic (
    .io_input_valid         (outputsAdapter_0_crossclock_fifo_io_pop_valid                      ), //i
    .io_input_ready         (outputsAdapter_0_sparseDownsizer_logic_io_input_ready              ), //o
    .io_input_payload_data  (outputsAdapter_0_crossclock_fifo_io_pop_payload_data[127:0]        ), //i
    .io_input_payload_mask  (outputsAdapter_0_crossclock_fifo_io_pop_payload_mask[15:0]         ), //i
    .io_input_payload_sink  (outputsAdapter_0_crossclock_fifo_io_pop_payload_sink[3:0]          ), //i
    .io_input_payload_last  (outputsAdapter_0_crossclock_fifo_io_pop_payload_last               ), //i
    .io_output_valid        (outputsAdapter_0_sparseDownsizer_logic_io_output_valid             ), //o
    .io_output_ready        (dat1_o_tready                                                      ), //i
    .io_output_payload_data (outputsAdapter_0_sparseDownsizer_logic_io_output_payload_data[63:0]), //o
    .io_output_payload_mask (outputsAdapter_0_sparseDownsizer_logic_io_output_payload_mask[7:0] ), //o
    .io_output_payload_sink (outputsAdapter_0_sparseDownsizer_logic_io_output_payload_sink[3:0] ), //o
    .io_output_payload_last (outputsAdapter_0_sparseDownsizer_logic_io_output_payload_last      ), //o
    .dat1_o_clk             (dat1_o_clk                                                         ), //i
    .dat1_o_reset           (dat1_o_reset                                                       )  //i
  );
  EfxDMA_StreamFifoCC_3 outputsAdapter_1_crossclock_fifo (
    .io_push_valid        (outputsAdapter_1_ptr_valid                                 ), //i
    .io_push_ready        (outputsAdapter_1_crossclock_fifo_io_push_ready             ), //o
    .io_push_payload_data (outputsAdapter_1_ptr_payload_data[127:0]                   ), //i
    .io_push_payload_mask (outputsAdapter_1_ptr_payload_mask[15:0]                    ), //i
    .io_push_payload_sink (outputsAdapter_1_ptr_payload_sink[3:0]                     ), //i
    .io_push_payload_last (outputsAdapter_1_ptr_payload_last                          ), //i
    .io_pop_valid         (outputsAdapter_1_crossclock_fifo_io_pop_valid              ), //o
    .io_pop_ready         (outputsAdapter_1_sparseDownsizer_logic_io_input_ready      ), //i
    .io_pop_payload_data  (outputsAdapter_1_crossclock_fifo_io_pop_payload_data[127:0]), //o
    .io_pop_payload_mask  (outputsAdapter_1_crossclock_fifo_io_pop_payload_mask[15:0] ), //o
    .io_pop_payload_sink  (outputsAdapter_1_crossclock_fifo_io_pop_payload_sink[3:0]  ), //o
    .io_pop_payload_last  (outputsAdapter_1_crossclock_fifo_io_pop_payload_last       ), //o
    .io_pushOccupancy     (outputsAdapter_1_crossclock_fifo_io_pushOccupancy[4:0]     ), //o
    .io_popOccupancy      (outputsAdapter_1_crossclock_fifo_io_popOccupancy[4:0]      ), //o
    .clk                  (clk                                                        ), //i
    .reset                (reset                                                      ), //i
    .dat3_o_clk           (dat3_o_clk                                                 ), //i
    .dat3_o_reset         (dat3_o_reset                                               )  //i
  );
  EfxDMA_BsbDownSizerSparse_1 outputsAdapter_1_sparseDownsizer_logic (
    .io_input_valid         (outputsAdapter_1_crossclock_fifo_io_pop_valid                      ), //i
    .io_input_ready         (outputsAdapter_1_sparseDownsizer_logic_io_input_ready              ), //o
    .io_input_payload_data  (outputsAdapter_1_crossclock_fifo_io_pop_payload_data[127:0]        ), //i
    .io_input_payload_mask  (outputsAdapter_1_crossclock_fifo_io_pop_payload_mask[15:0]         ), //i
    .io_input_payload_sink  (outputsAdapter_1_crossclock_fifo_io_pop_payload_sink[3:0]          ), //i
    .io_input_payload_last  (outputsAdapter_1_crossclock_fifo_io_pop_payload_last               ), //i
    .io_output_valid        (outputsAdapter_1_sparseDownsizer_logic_io_output_valid             ), //o
    .io_output_ready        (dat3_o_tready                                                      ), //i
    .io_output_payload_data (outputsAdapter_1_sparseDownsizer_logic_io_output_payload_data[31:0]), //o
    .io_output_payload_mask (outputsAdapter_1_sparseDownsizer_logic_io_output_payload_mask[3:0] ), //o
    .io_output_payload_sink (outputsAdapter_1_sparseDownsizer_logic_io_output_payload_sink[3:0] ), //o
    .io_output_payload_last (outputsAdapter_1_sparseDownsizer_logic_io_output_payload_last      ), //o
    .dat3_o_clk             (dat3_o_clk                                                         ), //i
    .dat3_o_reset           (dat3_o_reset                                                       )  //i
  );
  assign ctrl_PREADY = withCtrlCc_apbCc_io_input_PREADY;
  assign ctrl_PRDATA = withCtrlCc_apbCc_io_input_PRDATA;
  assign ctrl_PSLVERROR = withCtrlCc_apbCc_io_input_PSLVERROR;
  assign ctrl_interrupts = io_interrupts_buffercc_io_dataOut;
  assign io_write_cmd_s2mPipe_valid = (core_io_write_cmd_valid || (! io_write_cmd_rValidN));
  assign io_write_cmd_s2mPipe_payload_last = (io_write_cmd_rValidN ? core_io_write_cmd_payload_last : io_write_cmd_rData_last);
  assign io_write_cmd_s2mPipe_payload_fragment_source = (io_write_cmd_rValidN ? core_io_write_cmd_payload_fragment_source : io_write_cmd_rData_fragment_source);
  assign io_write_cmd_s2mPipe_payload_fragment_opcode = (io_write_cmd_rValidN ? core_io_write_cmd_payload_fragment_opcode : io_write_cmd_rData_fragment_opcode);
  assign io_write_cmd_s2mPipe_payload_fragment_address = (io_write_cmd_rValidN ? core_io_write_cmd_payload_fragment_address : io_write_cmd_rData_fragment_address);
  assign io_write_cmd_s2mPipe_payload_fragment_length = (io_write_cmd_rValidN ? core_io_write_cmd_payload_fragment_length : io_write_cmd_rData_fragment_length);
  assign io_write_cmd_s2mPipe_payload_fragment_data = (io_write_cmd_rValidN ? core_io_write_cmd_payload_fragment_data : io_write_cmd_rData_fragment_data);
  assign io_write_cmd_s2mPipe_payload_fragment_mask = (io_write_cmd_rValidN ? core_io_write_cmd_payload_fragment_mask : io_write_cmd_rData_fragment_mask);
  assign io_write_cmd_s2mPipe_payload_fragment_context = (io_write_cmd_rValidN ? core_io_write_cmd_payload_fragment_context : io_write_cmd_rData_fragment_context);
  always @(*) begin
    io_write_cmd_s2mPipe_ready = io_write_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375) begin
      io_write_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! io_write_cmd_s2mPipe_m2sPipe_valid);
  assign io_write_cmd_s2mPipe_m2sPipe_valid = io_write_cmd_s2mPipe_rValid;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_last = io_write_cmd_s2mPipe_rData_last;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_fragment_source = io_write_cmd_s2mPipe_rData_fragment_source;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_fragment_opcode = io_write_cmd_s2mPipe_rData_fragment_opcode;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_fragment_address = io_write_cmd_s2mPipe_rData_fragment_address;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_fragment_length = io_write_cmd_s2mPipe_rData_fragment_length;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_fragment_data = io_write_cmd_s2mPipe_rData_fragment_data;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_fragment_mask = io_write_cmd_s2mPipe_rData_fragment_mask;
  assign io_write_cmd_s2mPipe_m2sPipe_payload_fragment_context = io_write_cmd_s2mPipe_rData_fragment_context;
  assign io_write_cmd_s2mPipe_m2sPipe_ready = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign interconnect_read_aggregated_cmd_halfPipe_fire = (interconnect_read_aggregated_cmd_halfPipe_valid && interconnect_read_aggregated_cmd_halfPipe_ready);
  assign interconnect_read_aggregated_cmd_ready = (! interconnect_read_aggregated_cmd_rValid);
  assign interconnect_read_aggregated_cmd_halfPipe_valid = interconnect_read_aggregated_cmd_rValid;
  assign interconnect_read_aggregated_cmd_halfPipe_payload_last = interconnect_read_aggregated_cmd_rData_last;
  assign interconnect_read_aggregated_cmd_halfPipe_payload_fragment_source = interconnect_read_aggregated_cmd_rData_fragment_source;
  assign interconnect_read_aggregated_cmd_halfPipe_payload_fragment_opcode = interconnect_read_aggregated_cmd_rData_fragment_opcode;
  assign interconnect_read_aggregated_cmd_halfPipe_payload_fragment_address = interconnect_read_aggregated_cmd_rData_fragment_address;
  assign interconnect_read_aggregated_cmd_halfPipe_payload_fragment_length = interconnect_read_aggregated_cmd_rData_fragment_length;
  assign interconnect_read_aggregated_cmd_halfPipe_payload_fragment_context = interconnect_read_aggregated_cmd_rData_fragment_context;
  assign readLogic_resized_cmd_valid = interconnect_read_aggregated_cmd_halfPipe_valid;
  assign interconnect_read_aggregated_cmd_halfPipe_ready = readLogic_resized_cmd_ready;
  assign readLogic_resized_cmd_payload_last = interconnect_read_aggregated_cmd_halfPipe_payload_last;
  assign readLogic_resized_cmd_payload_fragment_source = interconnect_read_aggregated_cmd_halfPipe_payload_fragment_source;
  assign readLogic_resized_cmd_payload_fragment_opcode = interconnect_read_aggregated_cmd_halfPipe_payload_fragment_opcode;
  assign readLogic_resized_cmd_payload_fragment_address = interconnect_read_aggregated_cmd_halfPipe_payload_fragment_address;
  assign readLogic_resized_cmd_payload_fragment_length = interconnect_read_aggregated_cmd_halfPipe_payload_fragment_length;
  assign readLogic_resized_cmd_payload_fragment_context = interconnect_read_aggregated_cmd_halfPipe_payload_fragment_context;
  assign readLogic_resized_rsp_combStage_valid = readLogic_resized_rsp_valid;
  assign readLogic_resized_rsp_ready = readLogic_resized_rsp_combStage_ready;
  assign readLogic_resized_rsp_combStage_payload_last = readLogic_resized_rsp_payload_last;
  assign readLogic_resized_rsp_combStage_payload_fragment_source = readLogic_resized_rsp_payload_fragment_source;
  assign readLogic_resized_rsp_combStage_payload_fragment_opcode = readLogic_resized_rsp_payload_fragment_opcode;
  assign readLogic_resized_rsp_combStage_payload_fragment_data = readLogic_resized_rsp_payload_fragment_data;
  assign readLogic_resized_rsp_combStage_payload_fragment_context = readLogic_resized_rsp_payload_fragment_context;
  assign interconnect_read_aggregated_rsp_valid = readLogic_resized_rsp_combStage_valid;
  assign readLogic_resized_rsp_combStage_ready = interconnect_read_aggregated_rsp_ready;
  assign interconnect_read_aggregated_rsp_payload_last = readLogic_resized_rsp_combStage_payload_last;
  assign interconnect_read_aggregated_rsp_payload_fragment_source = readLogic_resized_rsp_combStage_payload_fragment_source;
  assign interconnect_read_aggregated_rsp_payload_fragment_opcode = readLogic_resized_rsp_combStage_payload_fragment_opcode;
  assign interconnect_read_aggregated_rsp_payload_fragment_data = readLogic_resized_rsp_combStage_payload_fragment_data;
  assign interconnect_read_aggregated_rsp_payload_fragment_context = readLogic_resized_rsp_combStage_payload_fragment_context;
  assign readLogic_resized_cmd_ready = readLogic_sourceRemover_io_input_cmd_ready;
  assign readLogic_resized_rsp_valid = readLogic_sourceRemover_io_input_rsp_valid;
  assign readLogic_resized_rsp_payload_last = readLogic_sourceRemover_io_input_rsp_payload_last;
  assign readLogic_resized_rsp_payload_fragment_source = readLogic_sourceRemover_io_input_rsp_payload_fragment_source;
  assign readLogic_resized_rsp_payload_fragment_opcode = readLogic_sourceRemover_io_input_rsp_payload_fragment_opcode;
  assign readLogic_resized_rsp_payload_fragment_data = readLogic_sourceRemover_io_input_rsp_payload_fragment_data;
  assign readLogic_resized_rsp_payload_fragment_context = readLogic_sourceRemover_io_input_rsp_payload_fragment_context;
  assign readLogic_adapter_ar_valid = readLogic_bridge_io_output_ar_valid;
  assign readLogic_adapter_ar_payload_addr = readLogic_bridge_io_output_ar_payload_addr;
  assign _zz_readLogic_adapter_ar_payload_region[3 : 0] = 4'b0000;
  assign readLogic_adapter_ar_payload_region = _zz_readLogic_adapter_ar_payload_region;
  assign readLogic_adapter_ar_payload_len = readLogic_bridge_io_output_ar_payload_len;
  assign readLogic_adapter_ar_payload_size = readLogic_bridge_io_output_ar_payload_size;
  assign readLogic_adapter_ar_payload_burst = 2'b01;
  assign readLogic_adapter_ar_payload_lock = 1'b0;
  assign readLogic_adapter_ar_payload_cache = readLogic_bridge_io_output_ar_payload_cache;
  assign readLogic_adapter_ar_payload_qos = 4'b0000;
  assign readLogic_adapter_ar_payload_prot = readLogic_bridge_io_output_ar_payload_prot;
  assign readLogic_adapter_r_ready = readLogic_bridge_io_output_r_ready;
  assign readLogic_adapter_ar_halfPipe_fire = (readLogic_adapter_ar_halfPipe_valid && readLogic_adapter_ar_halfPipe_ready);
  assign readLogic_adapter_ar_ready = (! readLogic_adapter_ar_rValid);
  assign readLogic_adapter_ar_halfPipe_valid = readLogic_adapter_ar_rValid;
  assign readLogic_adapter_ar_halfPipe_payload_addr = readLogic_adapter_ar_rData_addr;
  assign readLogic_adapter_ar_halfPipe_payload_region = readLogic_adapter_ar_rData_region;
  assign readLogic_adapter_ar_halfPipe_payload_len = readLogic_adapter_ar_rData_len;
  assign readLogic_adapter_ar_halfPipe_payload_size = readLogic_adapter_ar_rData_size;
  assign readLogic_adapter_ar_halfPipe_payload_burst = readLogic_adapter_ar_rData_burst;
  assign readLogic_adapter_ar_halfPipe_payload_lock = readLogic_adapter_ar_rData_lock;
  assign readLogic_adapter_ar_halfPipe_payload_cache = readLogic_adapter_ar_rData_cache;
  assign readLogic_adapter_ar_halfPipe_payload_qos = readLogic_adapter_ar_rData_qos;
  assign readLogic_adapter_ar_halfPipe_payload_prot = readLogic_adapter_ar_rData_prot;
  assign read_arvalid = readLogic_adapter_ar_halfPipe_valid;
  assign readLogic_adapter_ar_halfPipe_ready = read_arready;
  assign read_araddr = readLogic_adapter_ar_halfPipe_payload_addr;
  assign read_arregion = readLogic_adapter_ar_halfPipe_payload_region;
  assign read_arlen = readLogic_adapter_ar_halfPipe_payload_len;
  assign read_arsize = readLogic_adapter_ar_halfPipe_payload_size;
  assign read_arburst = readLogic_adapter_ar_halfPipe_payload_burst;
  assign read_arlock = readLogic_adapter_ar_halfPipe_payload_lock;
  assign read_arcache = readLogic_adapter_ar_halfPipe_payload_cache;
  assign read_arqos = readLogic_adapter_ar_halfPipe_payload_qos;
  assign read_arprot = readLogic_adapter_ar_halfPipe_payload_prot;
  assign read_rready = read_r_rValidN;
  assign read_r_s2mPipe_valid = (read_rvalid || (! read_r_rValidN));
  assign read_r_s2mPipe_payload_data = (read_r_rValidN ? read_rdata : read_r_rData_data);
  assign read_r_s2mPipe_payload_resp = (read_r_rValidN ? read_rresp : read_r_rData_resp);
  assign read_r_s2mPipe_payload_last = (read_r_rValidN ? read_rlast : read_r_rData_last);
  always @(*) begin
    read_r_s2mPipe_ready = readLogic_beforeQueue_ready;
    if(when_Stream_l375_1) begin
      read_r_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! readLogic_beforeQueue_valid);
  assign readLogic_beforeQueue_valid = read_r_s2mPipe_rValid;
  assign readLogic_beforeQueue_payload_data = read_r_s2mPipe_rData_data;
  assign readLogic_beforeQueue_payload_resp = read_r_s2mPipe_rData_resp;
  assign readLogic_beforeQueue_payload_last = read_r_s2mPipe_rData_last;
  assign readLogic_adapter_r_valid = readLogic_beforeQueue_valid;
  assign readLogic_beforeQueue_ready = readLogic_adapter_r_ready;
  assign readLogic_adapter_r_payload_data = readLogic_beforeQueue_payload_data;
  assign readLogic_adapter_r_payload_resp = readLogic_beforeQueue_payload_resp;
  assign readLogic_adapter_r_payload_last = readLogic_beforeQueue_payload_last;
  always @(*) begin
    interconnect_write_aggregated_cmd_ready = interconnect_write_aggregated_cmd_m2sPipe_ready;
    if(when_Stream_l375_2) begin
      interconnect_write_aggregated_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l375_2 = (! interconnect_write_aggregated_cmd_m2sPipe_valid);
  assign interconnect_write_aggregated_cmd_m2sPipe_valid = interconnect_write_aggregated_cmd_rValid;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_last = interconnect_write_aggregated_cmd_rData_last;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_source = interconnect_write_aggregated_cmd_rData_fragment_source;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_opcode = interconnect_write_aggregated_cmd_rData_fragment_opcode;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_address = interconnect_write_aggregated_cmd_rData_fragment_address;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_length = interconnect_write_aggregated_cmd_rData_fragment_length;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_data = interconnect_write_aggregated_cmd_rData_fragment_data;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_mask = interconnect_write_aggregated_cmd_rData_fragment_mask;
  assign interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_context = interconnect_write_aggregated_cmd_rData_fragment_context;
  assign writeLogic_resized_cmd_valid = interconnect_write_aggregated_cmd_m2sPipe_valid;
  assign interconnect_write_aggregated_cmd_m2sPipe_ready = writeLogic_resized_cmd_ready;
  assign writeLogic_resized_cmd_payload_last = interconnect_write_aggregated_cmd_m2sPipe_payload_last;
  assign writeLogic_resized_cmd_payload_fragment_source = interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_source;
  assign writeLogic_resized_cmd_payload_fragment_opcode = interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_opcode;
  assign writeLogic_resized_cmd_payload_fragment_address = interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_address;
  assign writeLogic_resized_cmd_payload_fragment_length = interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_length;
  assign writeLogic_resized_cmd_payload_fragment_data = interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_data;
  assign writeLogic_resized_cmd_payload_fragment_mask = interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_mask;
  assign writeLogic_resized_cmd_payload_fragment_context = interconnect_write_aggregated_cmd_m2sPipe_payload_fragment_context;
  assign writeLogic_resized_rsp_combStage_valid = writeLogic_resized_rsp_valid;
  assign writeLogic_resized_rsp_ready = writeLogic_resized_rsp_combStage_ready;
  assign writeLogic_resized_rsp_combStage_payload_last = writeLogic_resized_rsp_payload_last;
  assign writeLogic_resized_rsp_combStage_payload_fragment_source = writeLogic_resized_rsp_payload_fragment_source;
  assign writeLogic_resized_rsp_combStage_payload_fragment_opcode = writeLogic_resized_rsp_payload_fragment_opcode;
  assign writeLogic_resized_rsp_combStage_payload_fragment_context = writeLogic_resized_rsp_payload_fragment_context;
  assign interconnect_write_aggregated_rsp_valid = writeLogic_resized_rsp_combStage_valid;
  assign writeLogic_resized_rsp_combStage_ready = interconnect_write_aggregated_rsp_ready;
  assign interconnect_write_aggregated_rsp_payload_last = writeLogic_resized_rsp_combStage_payload_last;
  assign interconnect_write_aggregated_rsp_payload_fragment_source = writeLogic_resized_rsp_combStage_payload_fragment_source;
  assign interconnect_write_aggregated_rsp_payload_fragment_opcode = writeLogic_resized_rsp_combStage_payload_fragment_opcode;
  assign interconnect_write_aggregated_rsp_payload_fragment_context = writeLogic_resized_rsp_combStage_payload_fragment_context;
  assign writeLogic_resized_cmd_ready = writeLogic_sourceRemover_io_input_cmd_ready;
  assign writeLogic_resized_rsp_valid = writeLogic_sourceRemover_io_input_rsp_valid;
  assign writeLogic_resized_rsp_payload_last = writeLogic_sourceRemover_io_input_rsp_payload_last;
  assign writeLogic_resized_rsp_payload_fragment_source = writeLogic_sourceRemover_io_input_rsp_payload_fragment_source;
  assign writeLogic_resized_rsp_payload_fragment_opcode = writeLogic_sourceRemover_io_input_rsp_payload_fragment_opcode;
  assign writeLogic_resized_rsp_payload_fragment_context = writeLogic_sourceRemover_io_input_rsp_payload_fragment_context;
  assign writeLogic_adapter_aw_valid = writeLogic_bridge_io_output_aw_valid;
  assign writeLogic_adapter_aw_payload_addr = writeLogic_bridge_io_output_aw_payload_addr;
  assign _zz_writeLogic_adapter_aw_payload_region[3 : 0] = 4'b0000;
  assign writeLogic_adapter_aw_payload_region = _zz_writeLogic_adapter_aw_payload_region;
  assign writeLogic_adapter_aw_payload_len = writeLogic_bridge_io_output_aw_payload_len;
  assign writeLogic_adapter_aw_payload_size = writeLogic_bridge_io_output_aw_payload_size;
  assign writeLogic_adapter_aw_payload_burst = 2'b01;
  assign writeLogic_adapter_aw_payload_lock = 1'b0;
  assign writeLogic_adapter_aw_payload_cache = writeLogic_bridge_io_output_aw_payload_cache;
  assign writeLogic_adapter_aw_payload_qos = 4'b0000;
  assign writeLogic_adapter_aw_payload_prot = writeLogic_bridge_io_output_aw_payload_prot;
  assign writeLogic_adapter_w_valid = writeLogic_bridge_io_output_w_valid;
  assign writeLogic_adapter_w_payload_data = writeLogic_bridge_io_output_w_payload_data;
  assign writeLogic_adapter_w_payload_strb = writeLogic_bridge_io_output_w_payload_strb;
  assign writeLogic_adapter_w_payload_last = writeLogic_bridge_io_output_w_payload_last;
  assign writeLogic_adapter_b_ready = writeLogic_bridge_io_output_b_ready;
  assign writeLogic_adapter_aw_halfPipe_fire = (writeLogic_adapter_aw_halfPipe_valid && writeLogic_adapter_aw_halfPipe_ready);
  assign writeLogic_adapter_aw_ready = (! writeLogic_adapter_aw_rValid);
  assign writeLogic_adapter_aw_halfPipe_valid = writeLogic_adapter_aw_rValid;
  assign writeLogic_adapter_aw_halfPipe_payload_addr = writeLogic_adapter_aw_rData_addr;
  assign writeLogic_adapter_aw_halfPipe_payload_region = writeLogic_adapter_aw_rData_region;
  assign writeLogic_adapter_aw_halfPipe_payload_len = writeLogic_adapter_aw_rData_len;
  assign writeLogic_adapter_aw_halfPipe_payload_size = writeLogic_adapter_aw_rData_size;
  assign writeLogic_adapter_aw_halfPipe_payload_burst = writeLogic_adapter_aw_rData_burst;
  assign writeLogic_adapter_aw_halfPipe_payload_lock = writeLogic_adapter_aw_rData_lock;
  assign writeLogic_adapter_aw_halfPipe_payload_cache = writeLogic_adapter_aw_rData_cache;
  assign writeLogic_adapter_aw_halfPipe_payload_qos = writeLogic_adapter_aw_rData_qos;
  assign writeLogic_adapter_aw_halfPipe_payload_prot = writeLogic_adapter_aw_rData_prot;
  assign write_awvalid = writeLogic_adapter_aw_halfPipe_valid;
  assign writeLogic_adapter_aw_halfPipe_ready = write_awready;
  assign write_awaddr = writeLogic_adapter_aw_halfPipe_payload_addr;
  assign write_awregion = writeLogic_adapter_aw_halfPipe_payload_region;
  assign write_awlen = writeLogic_adapter_aw_halfPipe_payload_len;
  assign write_awsize = writeLogic_adapter_aw_halfPipe_payload_size;
  assign write_awburst = writeLogic_adapter_aw_halfPipe_payload_burst;
  assign write_awlock = writeLogic_adapter_aw_halfPipe_payload_lock;
  assign write_awcache = writeLogic_adapter_aw_halfPipe_payload_cache;
  assign write_awqos = writeLogic_adapter_aw_halfPipe_payload_qos;
  assign write_awprot = writeLogic_adapter_aw_halfPipe_payload_prot;
  assign writeLogic_adapter_w_ready = writeLogic_adapter_w_rValidN;
  assign writeLogic_adapter_w_s2mPipe_valid = (writeLogic_adapter_w_valid || (! writeLogic_adapter_w_rValidN));
  assign writeLogic_adapter_w_s2mPipe_payload_data = (writeLogic_adapter_w_rValidN ? writeLogic_adapter_w_payload_data : writeLogic_adapter_w_rData_data);
  assign writeLogic_adapter_w_s2mPipe_payload_strb = (writeLogic_adapter_w_rValidN ? writeLogic_adapter_w_payload_strb : writeLogic_adapter_w_rData_strb);
  assign writeLogic_adapter_w_s2mPipe_payload_last = (writeLogic_adapter_w_rValidN ? writeLogic_adapter_w_payload_last : writeLogic_adapter_w_rData_last);
  always @(*) begin
    writeLogic_adapter_w_s2mPipe_ready = writeLogic_adapter_w_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_3) begin
      writeLogic_adapter_w_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_3 = (! writeLogic_adapter_w_s2mPipe_m2sPipe_valid);
  assign writeLogic_adapter_w_s2mPipe_m2sPipe_valid = writeLogic_adapter_w_s2mPipe_rValid;
  assign writeLogic_adapter_w_s2mPipe_m2sPipe_payload_data = writeLogic_adapter_w_s2mPipe_rData_data;
  assign writeLogic_adapter_w_s2mPipe_m2sPipe_payload_strb = writeLogic_adapter_w_s2mPipe_rData_strb;
  assign writeLogic_adapter_w_s2mPipe_m2sPipe_payload_last = writeLogic_adapter_w_s2mPipe_rData_last;
  assign write_wvalid = writeLogic_adapter_w_s2mPipe_m2sPipe_valid;
  assign writeLogic_adapter_w_s2mPipe_m2sPipe_ready = write_wready;
  assign write_wdata = writeLogic_adapter_w_s2mPipe_m2sPipe_payload_data;
  assign write_wstrb = writeLogic_adapter_w_s2mPipe_m2sPipe_payload_strb;
  assign write_wlast = writeLogic_adapter_w_s2mPipe_m2sPipe_payload_last;
  assign write_b_halfPipe_fire = (write_b_halfPipe_valid && write_b_halfPipe_ready);
  assign write_bready = (! write_b_rValid);
  assign write_b_halfPipe_valid = write_b_rValid;
  assign write_b_halfPipe_payload_resp = write_b_rData_resp;
  assign writeLogic_adapter_b_valid = write_b_halfPipe_valid;
  assign write_b_halfPipe_ready = writeLogic_adapter_b_ready;
  assign writeLogic_adapter_b_payload_resp = write_b_halfPipe_payload_resp;
  assign dat0_i_tready = inputsAdapter_0_upsizer_logic_io_input_ready;
  assign io_pop_s2mPipe_valid = (inputsAdapter_0_crossclock_fifo_io_pop_valid || (! io_pop_rValidN));
  assign io_pop_s2mPipe_payload_data = (io_pop_rValidN ? inputsAdapter_0_crossclock_fifo_io_pop_payload_data : io_pop_rData_data);
  assign io_pop_s2mPipe_payload_mask = (io_pop_rValidN ? inputsAdapter_0_crossclock_fifo_io_pop_payload_mask : io_pop_rData_mask);
  assign io_pop_s2mPipe_payload_sink = (io_pop_rValidN ? inputsAdapter_0_crossclock_fifo_io_pop_payload_sink : io_pop_rData_sink);
  assign io_pop_s2mPipe_payload_last = (io_pop_rValidN ? inputsAdapter_0_crossclock_fifo_io_pop_payload_last : io_pop_rData_last);
  always @(*) begin
    io_pop_s2mPipe_ready = io_pop_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_4) begin
      io_pop_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_4 = (! io_pop_s2mPipe_m2sPipe_valid);
  assign io_pop_s2mPipe_m2sPipe_valid = io_pop_s2mPipe_rValid;
  assign io_pop_s2mPipe_m2sPipe_payload_data = io_pop_s2mPipe_rData_data;
  assign io_pop_s2mPipe_m2sPipe_payload_mask = io_pop_s2mPipe_rData_mask;
  assign io_pop_s2mPipe_m2sPipe_payload_sink = io_pop_s2mPipe_rData_sink;
  assign io_pop_s2mPipe_m2sPipe_payload_last = io_pop_s2mPipe_rData_last;
  assign io_pop_s2mPipe_m2sPipe_ready = core_io_inputs_0_ready;
  assign dat2_i_tready = inputsAdapter_1_upsizer_logic_io_input_ready;
  assign io_pop_s2mPipe_valid_1 = (inputsAdapter_1_crossclock_fifo_io_pop_valid || (! io_pop_rValidN_1));
  assign io_pop_s2mPipe_payload_data_1 = (io_pop_rValidN_1 ? inputsAdapter_1_crossclock_fifo_io_pop_payload_data : io_pop_rData_data_1);
  assign io_pop_s2mPipe_payload_mask_1 = (io_pop_rValidN_1 ? inputsAdapter_1_crossclock_fifo_io_pop_payload_mask : io_pop_rData_mask_1);
  assign io_pop_s2mPipe_payload_sink_1 = (io_pop_rValidN_1 ? inputsAdapter_1_crossclock_fifo_io_pop_payload_sink : io_pop_rData_sink_1);
  assign io_pop_s2mPipe_payload_last_1 = (io_pop_rValidN_1 ? inputsAdapter_1_crossclock_fifo_io_pop_payload_last : io_pop_rData_last_1);
  always @(*) begin
    io_pop_s2mPipe_ready_1 = io_pop_s2mPipe_m2sPipe_ready_1;
    if(when_Stream_l375_5) begin
      io_pop_s2mPipe_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_5 = (! io_pop_s2mPipe_m2sPipe_valid_1);
  assign io_pop_s2mPipe_m2sPipe_valid_1 = io_pop_s2mPipe_rValid_1;
  assign io_pop_s2mPipe_m2sPipe_payload_data_1 = io_pop_s2mPipe_rData_data_1;
  assign io_pop_s2mPipe_m2sPipe_payload_mask_1 = io_pop_s2mPipe_rData_mask_1;
  assign io_pop_s2mPipe_m2sPipe_payload_sink_1 = io_pop_s2mPipe_rData_sink_1;
  assign io_pop_s2mPipe_m2sPipe_payload_last_1 = io_pop_s2mPipe_rData_last_1;
  assign io_pop_s2mPipe_m2sPipe_ready_1 = core_io_inputs_1_ready;
  assign io_outputs_0_s2mPipe_valid = (core_io_outputs_0_valid || (! io_outputs_0_rValidN));
  assign io_outputs_0_s2mPipe_payload_data = (io_outputs_0_rValidN ? core_io_outputs_0_payload_data : io_outputs_0_rData_data);
  assign io_outputs_0_s2mPipe_payload_mask = (io_outputs_0_rValidN ? core_io_outputs_0_payload_mask : io_outputs_0_rData_mask);
  assign io_outputs_0_s2mPipe_payload_sink = (io_outputs_0_rValidN ? core_io_outputs_0_payload_sink : io_outputs_0_rData_sink);
  assign io_outputs_0_s2mPipe_payload_last = (io_outputs_0_rValidN ? core_io_outputs_0_payload_last : io_outputs_0_rData_last);
  always @(*) begin
    io_outputs_0_s2mPipe_ready = outputsAdapter_0_ptr_ready;
    if(when_Stream_l375_6) begin
      io_outputs_0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_6 = (! outputsAdapter_0_ptr_valid);
  assign outputsAdapter_0_ptr_valid = io_outputs_0_s2mPipe_rValid;
  assign outputsAdapter_0_ptr_payload_data = io_outputs_0_s2mPipe_rData_data;
  assign outputsAdapter_0_ptr_payload_mask = io_outputs_0_s2mPipe_rData_mask;
  assign outputsAdapter_0_ptr_payload_sink = io_outputs_0_s2mPipe_rData_sink;
  assign outputsAdapter_0_ptr_payload_last = io_outputs_0_s2mPipe_rData_last;
  assign outputsAdapter_0_ptr_ready = outputsAdapter_0_crossclock_fifo_io_push_ready;
  assign dat1_o_tvalid = outputsAdapter_0_sparseDownsizer_logic_io_output_valid;
  assign dat1_o_tdata = outputsAdapter_0_sparseDownsizer_logic_io_output_payload_data;
  assign dat1_o_tkeep = outputsAdapter_0_sparseDownsizer_logic_io_output_payload_mask;
  assign dat1_o_tdest = outputsAdapter_0_sparseDownsizer_logic_io_output_payload_sink;
  assign dat1_o_tlast = outputsAdapter_0_sparseDownsizer_logic_io_output_payload_last;
  assign io_outputs_1_s2mPipe_valid = (core_io_outputs_1_valid || (! io_outputs_1_rValidN));
  assign io_outputs_1_s2mPipe_payload_data = (io_outputs_1_rValidN ? core_io_outputs_1_payload_data : io_outputs_1_rData_data);
  assign io_outputs_1_s2mPipe_payload_mask = (io_outputs_1_rValidN ? core_io_outputs_1_payload_mask : io_outputs_1_rData_mask);
  assign io_outputs_1_s2mPipe_payload_sink = (io_outputs_1_rValidN ? core_io_outputs_1_payload_sink : io_outputs_1_rData_sink);
  assign io_outputs_1_s2mPipe_payload_last = (io_outputs_1_rValidN ? core_io_outputs_1_payload_last : io_outputs_1_rData_last);
  always @(*) begin
    io_outputs_1_s2mPipe_ready = outputsAdapter_1_ptr_ready;
    if(when_Stream_l375_7) begin
      io_outputs_1_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_7 = (! outputsAdapter_1_ptr_valid);
  assign outputsAdapter_1_ptr_valid = io_outputs_1_s2mPipe_rValid;
  assign outputsAdapter_1_ptr_payload_data = io_outputs_1_s2mPipe_rData_data;
  assign outputsAdapter_1_ptr_payload_mask = io_outputs_1_s2mPipe_rData_mask;
  assign outputsAdapter_1_ptr_payload_sink = io_outputs_1_s2mPipe_rData_sink;
  assign outputsAdapter_1_ptr_payload_last = io_outputs_1_s2mPipe_rData_last;
  assign outputsAdapter_1_ptr_ready = outputsAdapter_1_crossclock_fifo_io_push_ready;
  assign dat3_o_tvalid = outputsAdapter_1_sparseDownsizer_logic_io_output_valid;
  assign dat3_o_tdata = outputsAdapter_1_sparseDownsizer_logic_io_output_payload_data;
  assign dat3_o_tkeep = outputsAdapter_1_sparseDownsizer_logic_io_output_payload_mask;
  assign dat3_o_tdest = outputsAdapter_1_sparseDownsizer_logic_io_output_payload_sink;
  assign dat3_o_tlast = outputsAdapter_1_sparseDownsizer_logic_io_output_payload_last;
  assign interconnect_read_aggregated_cmd_valid = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = interconnect_read_aggregated_cmd_ready;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = interconnect_read_aggregated_rsp_valid;
  assign interconnect_read_aggregated_rsp_ready = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  assign interconnect_read_aggregated_cmd_payload_last = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = interconnect_read_aggregated_rsp_payload_last;
  assign interconnect_read_aggregated_cmd_payload_fragment_source = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  assign interconnect_read_aggregated_cmd_payload_fragment_opcode = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  assign interconnect_read_aggregated_cmd_payload_fragment_address = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  assign interconnect_read_aggregated_cmd_payload_fragment_length = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  assign interconnect_read_aggregated_cmd_payload_fragment_context = interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = interconnect_read_aggregated_rsp_payload_fragment_source;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = interconnect_read_aggregated_rsp_payload_fragment_opcode;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = interconnect_read_aggregated_rsp_payload_fragment_data;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = interconnect_read_aggregated_rsp_payload_fragment_context;
  assign interconnect_write_aggregated_cmd_valid = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = interconnect_write_aggregated_cmd_ready;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = interconnect_write_aggregated_rsp_valid;
  assign interconnect_write_aggregated_rsp_ready = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  assign interconnect_write_aggregated_cmd_payload_last = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = interconnect_write_aggregated_rsp_payload_last;
  assign interconnect_write_aggregated_cmd_payload_fragment_source = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  assign interconnect_write_aggregated_cmd_payload_fragment_opcode = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  assign interconnect_write_aggregated_cmd_payload_fragment_address = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  assign interconnect_write_aggregated_cmd_payload_fragment_length = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  assign interconnect_write_aggregated_cmd_payload_fragment_data = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  assign interconnect_write_aggregated_cmd_payload_fragment_mask = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  assign interconnect_write_aggregated_cmd_payload_fragment_context = interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = interconnect_write_aggregated_rsp_payload_fragment_source;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = interconnect_write_aggregated_rsp_payload_fragment_opcode;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = interconnect_write_aggregated_rsp_payload_fragment_context;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = core_io_read_cmd_valid;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = core_io_read_rsp_ready;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = core_io_read_cmd_payload_last;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source = core_io_read_cmd_payload_fragment_source;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = core_io_read_cmd_payload_fragment_opcode;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = core_io_read_cmd_payload_fragment_address;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = core_io_read_cmd_payload_fragment_length;
  assign interconnect_read_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = core_io_read_cmd_payload_fragment_context;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = io_write_cmd_s2mPipe_m2sPipe_valid;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = core_io_write_rsp_ready;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = io_write_cmd_s2mPipe_m2sPipe_payload_last;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source = io_write_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = io_write_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = io_write_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = io_write_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = io_write_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = io_write_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  assign interconnect_write_aggregated_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = io_write_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  always @(posedge clk) begin
    if(reset) begin
      io_write_cmd_rValidN <= 1'b1;
      io_write_cmd_s2mPipe_rValid <= 1'b0;
      interconnect_read_aggregated_cmd_rValid <= 1'b0;
      readLogic_adapter_ar_rValid <= 1'b0;
      read_r_rValidN <= 1'b1;
      read_r_s2mPipe_rValid <= 1'b0;
      interconnect_write_aggregated_cmd_rValid <= 1'b0;
      writeLogic_adapter_aw_rValid <= 1'b0;
      writeLogic_adapter_w_rValidN <= 1'b1;
      writeLogic_adapter_w_s2mPipe_rValid <= 1'b0;
      write_b_rValid <= 1'b0;
      io_pop_rValidN <= 1'b1;
      io_pop_s2mPipe_rValid <= 1'b0;
      io_pop_rValidN_1 <= 1'b1;
      io_pop_s2mPipe_rValid_1 <= 1'b0;
      io_outputs_0_rValidN <= 1'b1;
      io_outputs_0_s2mPipe_rValid <= 1'b0;
      io_outputs_1_rValidN <= 1'b1;
      io_outputs_1_s2mPipe_rValid <= 1'b0;
    end else begin
      if(core_io_write_cmd_valid) begin
        io_write_cmd_rValidN <= 1'b0;
      end
      if(io_write_cmd_s2mPipe_ready) begin
        io_write_cmd_rValidN <= 1'b1;
      end
      if(io_write_cmd_s2mPipe_ready) begin
        io_write_cmd_s2mPipe_rValid <= io_write_cmd_s2mPipe_valid;
      end
      if(interconnect_read_aggregated_cmd_valid) begin
        interconnect_read_aggregated_cmd_rValid <= 1'b1;
      end
      if(interconnect_read_aggregated_cmd_halfPipe_fire) begin
        interconnect_read_aggregated_cmd_rValid <= 1'b0;
      end
      if(readLogic_adapter_ar_valid) begin
        readLogic_adapter_ar_rValid <= 1'b1;
      end
      if(readLogic_adapter_ar_halfPipe_fire) begin
        readLogic_adapter_ar_rValid <= 1'b0;
      end
      if(read_rvalid) begin
        read_r_rValidN <= 1'b0;
      end
      if(read_r_s2mPipe_ready) begin
        read_r_rValidN <= 1'b1;
      end
      if(read_r_s2mPipe_ready) begin
        read_r_s2mPipe_rValid <= read_r_s2mPipe_valid;
      end
      if(interconnect_write_aggregated_cmd_ready) begin
        interconnect_write_aggregated_cmd_rValid <= interconnect_write_aggregated_cmd_valid;
      end
      if(writeLogic_adapter_aw_valid) begin
        writeLogic_adapter_aw_rValid <= 1'b1;
      end
      if(writeLogic_adapter_aw_halfPipe_fire) begin
        writeLogic_adapter_aw_rValid <= 1'b0;
      end
      if(writeLogic_adapter_w_valid) begin
        writeLogic_adapter_w_rValidN <= 1'b0;
      end
      if(writeLogic_adapter_w_s2mPipe_ready) begin
        writeLogic_adapter_w_rValidN <= 1'b1;
      end
      if(writeLogic_adapter_w_s2mPipe_ready) begin
        writeLogic_adapter_w_s2mPipe_rValid <= writeLogic_adapter_w_s2mPipe_valid;
      end
      if(write_bvalid) begin
        write_b_rValid <= 1'b1;
      end
      if(write_b_halfPipe_fire) begin
        write_b_rValid <= 1'b0;
      end
      if(inputsAdapter_0_crossclock_fifo_io_pop_valid) begin
        io_pop_rValidN <= 1'b0;
      end
      if(io_pop_s2mPipe_ready) begin
        io_pop_rValidN <= 1'b1;
      end
      if(io_pop_s2mPipe_ready) begin
        io_pop_s2mPipe_rValid <= io_pop_s2mPipe_valid;
      end
      if(inputsAdapter_1_crossclock_fifo_io_pop_valid) begin
        io_pop_rValidN_1 <= 1'b0;
      end
      if(io_pop_s2mPipe_ready_1) begin
        io_pop_rValidN_1 <= 1'b1;
      end
      if(io_pop_s2mPipe_ready_1) begin
        io_pop_s2mPipe_rValid_1 <= io_pop_s2mPipe_valid_1;
      end
      if(core_io_outputs_0_valid) begin
        io_outputs_0_rValidN <= 1'b0;
      end
      if(io_outputs_0_s2mPipe_ready) begin
        io_outputs_0_rValidN <= 1'b1;
      end
      if(io_outputs_0_s2mPipe_ready) begin
        io_outputs_0_s2mPipe_rValid <= io_outputs_0_s2mPipe_valid;
      end
      if(core_io_outputs_1_valid) begin
        io_outputs_1_rValidN <= 1'b0;
      end
      if(io_outputs_1_s2mPipe_ready) begin
        io_outputs_1_rValidN <= 1'b1;
      end
      if(io_outputs_1_s2mPipe_ready) begin
        io_outputs_1_s2mPipe_rValid <= io_outputs_1_s2mPipe_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(io_write_cmd_rValidN) begin
      io_write_cmd_rData_last <= core_io_write_cmd_payload_last;
      io_write_cmd_rData_fragment_source <= core_io_write_cmd_payload_fragment_source;
      io_write_cmd_rData_fragment_opcode <= core_io_write_cmd_payload_fragment_opcode;
      io_write_cmd_rData_fragment_address <= core_io_write_cmd_payload_fragment_address;
      io_write_cmd_rData_fragment_length <= core_io_write_cmd_payload_fragment_length;
      io_write_cmd_rData_fragment_data <= core_io_write_cmd_payload_fragment_data;
      io_write_cmd_rData_fragment_mask <= core_io_write_cmd_payload_fragment_mask;
      io_write_cmd_rData_fragment_context <= core_io_write_cmd_payload_fragment_context;
    end
    if(io_write_cmd_s2mPipe_ready) begin
      io_write_cmd_s2mPipe_rData_last <= io_write_cmd_s2mPipe_payload_last;
      io_write_cmd_s2mPipe_rData_fragment_source <= io_write_cmd_s2mPipe_payload_fragment_source;
      io_write_cmd_s2mPipe_rData_fragment_opcode <= io_write_cmd_s2mPipe_payload_fragment_opcode;
      io_write_cmd_s2mPipe_rData_fragment_address <= io_write_cmd_s2mPipe_payload_fragment_address;
      io_write_cmd_s2mPipe_rData_fragment_length <= io_write_cmd_s2mPipe_payload_fragment_length;
      io_write_cmd_s2mPipe_rData_fragment_data <= io_write_cmd_s2mPipe_payload_fragment_data;
      io_write_cmd_s2mPipe_rData_fragment_mask <= io_write_cmd_s2mPipe_payload_fragment_mask;
      io_write_cmd_s2mPipe_rData_fragment_context <= io_write_cmd_s2mPipe_payload_fragment_context;
    end
    if(interconnect_read_aggregated_cmd_ready) begin
      interconnect_read_aggregated_cmd_rData_last <= interconnect_read_aggregated_cmd_payload_last;
      interconnect_read_aggregated_cmd_rData_fragment_source <= interconnect_read_aggregated_cmd_payload_fragment_source;
      interconnect_read_aggregated_cmd_rData_fragment_opcode <= interconnect_read_aggregated_cmd_payload_fragment_opcode;
      interconnect_read_aggregated_cmd_rData_fragment_address <= interconnect_read_aggregated_cmd_payload_fragment_address;
      interconnect_read_aggregated_cmd_rData_fragment_length <= interconnect_read_aggregated_cmd_payload_fragment_length;
      interconnect_read_aggregated_cmd_rData_fragment_context <= interconnect_read_aggregated_cmd_payload_fragment_context;
    end
    if(readLogic_adapter_ar_ready) begin
      readLogic_adapter_ar_rData_addr <= readLogic_adapter_ar_payload_addr;
      readLogic_adapter_ar_rData_region <= readLogic_adapter_ar_payload_region;
      readLogic_adapter_ar_rData_len <= readLogic_adapter_ar_payload_len;
      readLogic_adapter_ar_rData_size <= readLogic_adapter_ar_payload_size;
      readLogic_adapter_ar_rData_burst <= readLogic_adapter_ar_payload_burst;
      readLogic_adapter_ar_rData_lock <= readLogic_adapter_ar_payload_lock;
      readLogic_adapter_ar_rData_cache <= readLogic_adapter_ar_payload_cache;
      readLogic_adapter_ar_rData_qos <= readLogic_adapter_ar_payload_qos;
      readLogic_adapter_ar_rData_prot <= readLogic_adapter_ar_payload_prot;
    end
    if(read_rready) begin
      read_r_rData_data <= read_rdata;
      read_r_rData_resp <= read_rresp;
      read_r_rData_last <= read_rlast;
    end
    if(read_r_s2mPipe_ready) begin
      read_r_s2mPipe_rData_data <= read_r_s2mPipe_payload_data;
      read_r_s2mPipe_rData_resp <= read_r_s2mPipe_payload_resp;
      read_r_s2mPipe_rData_last <= read_r_s2mPipe_payload_last;
    end
    if(interconnect_write_aggregated_cmd_ready) begin
      interconnect_write_aggregated_cmd_rData_last <= interconnect_write_aggregated_cmd_payload_last;
      interconnect_write_aggregated_cmd_rData_fragment_source <= interconnect_write_aggregated_cmd_payload_fragment_source;
      interconnect_write_aggregated_cmd_rData_fragment_opcode <= interconnect_write_aggregated_cmd_payload_fragment_opcode;
      interconnect_write_aggregated_cmd_rData_fragment_address <= interconnect_write_aggregated_cmd_payload_fragment_address;
      interconnect_write_aggregated_cmd_rData_fragment_length <= interconnect_write_aggregated_cmd_payload_fragment_length;
      interconnect_write_aggregated_cmd_rData_fragment_data <= interconnect_write_aggregated_cmd_payload_fragment_data;
      interconnect_write_aggregated_cmd_rData_fragment_mask <= interconnect_write_aggregated_cmd_payload_fragment_mask;
      interconnect_write_aggregated_cmd_rData_fragment_context <= interconnect_write_aggregated_cmd_payload_fragment_context;
    end
    if(writeLogic_adapter_aw_ready) begin
      writeLogic_adapter_aw_rData_addr <= writeLogic_adapter_aw_payload_addr;
      writeLogic_adapter_aw_rData_region <= writeLogic_adapter_aw_payload_region;
      writeLogic_adapter_aw_rData_len <= writeLogic_adapter_aw_payload_len;
      writeLogic_adapter_aw_rData_size <= writeLogic_adapter_aw_payload_size;
      writeLogic_adapter_aw_rData_burst <= writeLogic_adapter_aw_payload_burst;
      writeLogic_adapter_aw_rData_lock <= writeLogic_adapter_aw_payload_lock;
      writeLogic_adapter_aw_rData_cache <= writeLogic_adapter_aw_payload_cache;
      writeLogic_adapter_aw_rData_qos <= writeLogic_adapter_aw_payload_qos;
      writeLogic_adapter_aw_rData_prot <= writeLogic_adapter_aw_payload_prot;
    end
    if(writeLogic_adapter_w_ready) begin
      writeLogic_adapter_w_rData_data <= writeLogic_adapter_w_payload_data;
      writeLogic_adapter_w_rData_strb <= writeLogic_adapter_w_payload_strb;
      writeLogic_adapter_w_rData_last <= writeLogic_adapter_w_payload_last;
    end
    if(writeLogic_adapter_w_s2mPipe_ready) begin
      writeLogic_adapter_w_s2mPipe_rData_data <= writeLogic_adapter_w_s2mPipe_payload_data;
      writeLogic_adapter_w_s2mPipe_rData_strb <= writeLogic_adapter_w_s2mPipe_payload_strb;
      writeLogic_adapter_w_s2mPipe_rData_last <= writeLogic_adapter_w_s2mPipe_payload_last;
    end
    if(write_bready) begin
      write_b_rData_resp <= write_bresp;
    end
    if(io_pop_rValidN) begin
      io_pop_rData_data <= inputsAdapter_0_crossclock_fifo_io_pop_payload_data;
      io_pop_rData_mask <= inputsAdapter_0_crossclock_fifo_io_pop_payload_mask;
      io_pop_rData_sink <= inputsAdapter_0_crossclock_fifo_io_pop_payload_sink;
      io_pop_rData_last <= inputsAdapter_0_crossclock_fifo_io_pop_payload_last;
    end
    if(io_pop_s2mPipe_ready) begin
      io_pop_s2mPipe_rData_data <= io_pop_s2mPipe_payload_data;
      io_pop_s2mPipe_rData_mask <= io_pop_s2mPipe_payload_mask;
      io_pop_s2mPipe_rData_sink <= io_pop_s2mPipe_payload_sink;
      io_pop_s2mPipe_rData_last <= io_pop_s2mPipe_payload_last;
    end
    if(io_pop_rValidN_1) begin
      io_pop_rData_data_1 <= inputsAdapter_1_crossclock_fifo_io_pop_payload_data;
      io_pop_rData_mask_1 <= inputsAdapter_1_crossclock_fifo_io_pop_payload_mask;
      io_pop_rData_sink_1 <= inputsAdapter_1_crossclock_fifo_io_pop_payload_sink;
      io_pop_rData_last_1 <= inputsAdapter_1_crossclock_fifo_io_pop_payload_last;
    end
    if(io_pop_s2mPipe_ready_1) begin
      io_pop_s2mPipe_rData_data_1 <= io_pop_s2mPipe_payload_data_1;
      io_pop_s2mPipe_rData_mask_1 <= io_pop_s2mPipe_payload_mask_1;
      io_pop_s2mPipe_rData_sink_1 <= io_pop_s2mPipe_payload_sink_1;
      io_pop_s2mPipe_rData_last_1 <= io_pop_s2mPipe_payload_last_1;
    end
    if(io_outputs_0_rValidN) begin
      io_outputs_0_rData_data <= core_io_outputs_0_payload_data;
      io_outputs_0_rData_mask <= core_io_outputs_0_payload_mask;
      io_outputs_0_rData_sink <= core_io_outputs_0_payload_sink;
      io_outputs_0_rData_last <= core_io_outputs_0_payload_last;
    end
    if(io_outputs_0_s2mPipe_ready) begin
      io_outputs_0_s2mPipe_rData_data <= io_outputs_0_s2mPipe_payload_data;
      io_outputs_0_s2mPipe_rData_mask <= io_outputs_0_s2mPipe_payload_mask;
      io_outputs_0_s2mPipe_rData_sink <= io_outputs_0_s2mPipe_payload_sink;
      io_outputs_0_s2mPipe_rData_last <= io_outputs_0_s2mPipe_payload_last;
    end
    if(io_outputs_1_rValidN) begin
      io_outputs_1_rData_data <= core_io_outputs_1_payload_data;
      io_outputs_1_rData_mask <= core_io_outputs_1_payload_mask;
      io_outputs_1_rData_sink <= core_io_outputs_1_payload_sink;
      io_outputs_1_rData_last <= core_io_outputs_1_payload_last;
    end
    if(io_outputs_1_s2mPipe_ready) begin
      io_outputs_1_s2mPipe_rData_data <= io_outputs_1_s2mPipe_payload_data;
      io_outputs_1_s2mPipe_rData_mask <= io_outputs_1_s2mPipe_payload_mask;
      io_outputs_1_s2mPipe_rData_sink <= io_outputs_1_s2mPipe_payload_sink;
      io_outputs_1_s2mPipe_rData_last <= io_outputs_1_s2mPipe_payload_last;
    end
  end


endmodule

module EfxDMA_BsbDownSizerSparse_1 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [127:0]  io_input_payload_data,
  input  wire [15:0]   io_input_payload_mask,
  input  wire [3:0]    io_input_payload_sink,
  input  wire          io_input_payload_last,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_data,
  output wire [3:0]    io_output_payload_mask,
  output wire [3:0]    io_output_payload_sink,
  output wire          io_output_payload_last,
  input  wire          dat3_o_clk,
  input  wire          dat3_o_reset
);

  reg        [31:0]   _zz_io_output_payload_data;
  reg        [3:0]    _zz_io_output_payload_mask;
  reg        [1:0]    counter;
  wire                end_1;
  wire                io_output_fire;

  always @(*) begin
    case(counter)
      2'b00 : begin
        _zz_io_output_payload_data = io_input_payload_data[31 : 0];
        _zz_io_output_payload_mask = io_input_payload_mask[3 : 0];
      end
      2'b01 : begin
        _zz_io_output_payload_data = io_input_payload_data[63 : 32];
        _zz_io_output_payload_mask = io_input_payload_mask[7 : 4];
      end
      2'b10 : begin
        _zz_io_output_payload_data = io_input_payload_data[95 : 64];
        _zz_io_output_payload_mask = io_input_payload_mask[11 : 8];
      end
      default : begin
        _zz_io_output_payload_data = io_input_payload_data[127 : 96];
        _zz_io_output_payload_mask = io_input_payload_mask[15 : 12];
      end
    endcase
  end

  assign end_1 = (counter == 2'b11);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_ready = (io_output_ready && end_1);
  assign io_output_valid = io_input_valid;
  assign io_output_payload_data = _zz_io_output_payload_data;
  assign io_output_payload_mask = _zz_io_output_payload_mask;
  assign io_output_payload_sink = io_input_payload_sink;
  assign io_output_payload_last = (io_input_payload_last && end_1);
  always @(posedge dat3_o_clk) begin
    if(dat3_o_reset) begin
      counter <= 2'b00;
    end else begin
      if(io_output_fire) begin
        counter <= (counter + 2'b01);
      end
    end
  end


endmodule

module EfxDMA_StreamFifoCC_3 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [127:0]  io_push_payload_data,
  input  wire [15:0]   io_push_payload_mask,
  input  wire [3:0]    io_push_payload_sink,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [127:0]  io_pop_payload_data,
  output wire [15:0]   io_pop_payload_mask,
  output wire [3:0]    io_pop_payload_sink,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          clk,
  input  wire          reset,
  input  wire          dat3_o_clk,
  input  wire          dat3_o_reset
);

  reg        [148:0]  ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [148:0]  _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [127:0]  popCC_readPort_rsp_data;
  wire       [15:0]   popCC_readPort_rsp_mask;
  wire       [3:0]    popCC_readPort_rsp_sink;
  wire                popCC_readPort_rsp_last;
  wire       [148:0]  _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [127:0]  popCC_readArbitation_translated_payload_data;
  wire       [15:0]   popCC_readArbitation_translated_payload_mask;
  wire       [3:0]    popCC_readArbitation_translated_payload_sink;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [148:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_sink,{io_push_payload_mask,io_push_payload_data}}};
  always @(posedge clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge dat3_o_clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_3 popToPushGray_buffercc (
    .io_dataIn  (popToPushGray[4:0]                    ), //i
    .io_dataOut (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .clk        (clk                                   ), //i
    .reset      (reset                                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_9 pushToPopGray_buffercc (
    .io_dataIn    (pushToPopGray[4:0]                    ), //i
    .io_dataOut   (pushToPopGray_buffercc_io_dataOut[4:0]), //o
    .dat3_o_clk   (dat3_o_clk                            ), //i
    .dat3_o_reset (dat3_o_reset                          )  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[127 : 0];
  assign popCC_readPort_rsp_mask = _zz_popCC_readPort_rsp_data[143 : 128];
  assign popCC_readPort_rsp_sink = _zz_popCC_readPort_rsp_data[147 : 144];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[148];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_mask = popCC_readPort_rsp_mask;
  assign popCC_readArbitation_translated_payload_sink = popCC_readPort_rsp_sink;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_mask = popCC_readArbitation_translated_payload_mask;
  assign io_pop_payload_sink = popCC_readArbitation_translated_payload_sink;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge clk) begin
    if(reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge dat3_o_clk) begin
    if(dat3_o_reset) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge dat3_o_clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module EfxDMA_BsbDownSizerSparse (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [127:0]  io_input_payload_data,
  input  wire [15:0]   io_input_payload_mask,
  input  wire [3:0]    io_input_payload_sink,
  input  wire          io_input_payload_last,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [63:0]   io_output_payload_data,
  output wire [7:0]    io_output_payload_mask,
  output wire [3:0]    io_output_payload_sink,
  output wire          io_output_payload_last,
  input  wire          dat1_o_clk,
  input  wire          dat1_o_reset
);

  reg        [63:0]   _zz_io_output_payload_data;
  reg        [7:0]    _zz_io_output_payload_mask;
  reg        [0:0]    counter;
  wire                end_1;
  wire                io_output_fire;

  always @(*) begin
    case(counter)
      1'b0 : begin
        _zz_io_output_payload_data = io_input_payload_data[63 : 0];
        _zz_io_output_payload_mask = io_input_payload_mask[7 : 0];
      end
      default : begin
        _zz_io_output_payload_data = io_input_payload_data[127 : 64];
        _zz_io_output_payload_mask = io_input_payload_mask[15 : 8];
      end
    endcase
  end

  assign end_1 = (counter == 1'b1);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_ready = (io_output_ready && end_1);
  assign io_output_valid = io_input_valid;
  assign io_output_payload_data = _zz_io_output_payload_data;
  assign io_output_payload_mask = _zz_io_output_payload_mask;
  assign io_output_payload_sink = io_input_payload_sink;
  assign io_output_payload_last = (io_input_payload_last && end_1);
  always @(posedge dat1_o_clk) begin
    if(dat1_o_reset) begin
      counter <= 1'b0;
    end else begin
      if(io_output_fire) begin
        counter <= (counter + 1'b1);
      end
    end
  end


endmodule

module EfxDMA_StreamFifoCC_2 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [127:0]  io_push_payload_data,
  input  wire [15:0]   io_push_payload_mask,
  input  wire [3:0]    io_push_payload_sink,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [127:0]  io_pop_payload_data,
  output wire [15:0]   io_pop_payload_mask,
  output wire [3:0]    io_pop_payload_sink,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          clk,
  input  wire          reset,
  input  wire          dat1_o_clk,
  input  wire          dat1_o_reset
);

  reg        [148:0]  ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [148:0]  _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [127:0]  popCC_readPort_rsp_data;
  wire       [15:0]   popCC_readPort_rsp_mask;
  wire       [3:0]    popCC_readPort_rsp_sink;
  wire                popCC_readPort_rsp_last;
  wire       [148:0]  _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [127:0]  popCC_readArbitation_translated_payload_data;
  wire       [15:0]   popCC_readArbitation_translated_payload_mask;
  wire       [3:0]    popCC_readArbitation_translated_payload_sink;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [148:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_sink,{io_push_payload_mask,io_push_payload_data}}};
  always @(posedge clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge dat1_o_clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_3 popToPushGray_buffercc (
    .io_dataIn  (popToPushGray[4:0]                    ), //i
    .io_dataOut (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .clk        (clk                                   ), //i
    .reset      (reset                                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_7 pushToPopGray_buffercc (
    .io_dataIn    (pushToPopGray[4:0]                    ), //i
    .io_dataOut   (pushToPopGray_buffercc_io_dataOut[4:0]), //o
    .dat1_o_clk   (dat1_o_clk                            ), //i
    .dat1_o_reset (dat1_o_reset                          )  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[127 : 0];
  assign popCC_readPort_rsp_mask = _zz_popCC_readPort_rsp_data[143 : 128];
  assign popCC_readPort_rsp_sink = _zz_popCC_readPort_rsp_data[147 : 144];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[148];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_mask = popCC_readPort_rsp_mask;
  assign popCC_readArbitation_translated_payload_sink = popCC_readPort_rsp_sink;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_mask = popCC_readArbitation_translated_payload_mask;
  assign io_pop_payload_sink = popCC_readArbitation_translated_payload_sink;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge clk) begin
    if(reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge dat1_o_clk) begin
    if(dat1_o_reset) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge dat1_o_clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module EfxDMA_StreamFifoCC_1 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [127:0]  io_push_payload_data,
  input  wire [15:0]   io_push_payload_mask,
  input  wire [3:0]    io_push_payload_sink,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [127:0]  io_pop_payload_data,
  output wire [15:0]   io_pop_payload_mask,
  output wire [3:0]    io_pop_payload_sink,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          dat2_i_clk,
  input  wire          dat2_i_reset,
  input  wire          clk,
  input  wire          reset
);

  reg        [148:0]  ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [148:0]  _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [127:0]  popCC_readPort_rsp_data;
  wire       [15:0]   popCC_readPort_rsp_mask;
  wire       [3:0]    popCC_readPort_rsp_sink;
  wire                popCC_readPort_rsp_last;
  wire       [148:0]  _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [127:0]  popCC_readArbitation_translated_payload_data;
  wire       [15:0]   popCC_readArbitation_translated_payload_mask;
  wire       [3:0]    popCC_readArbitation_translated_payload_sink;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [148:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_sink,{io_push_payload_mask,io_push_payload_data}}};
  always @(posedge dat2_i_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_4 popToPushGray_buffercc (
    .io_dataIn    (popToPushGray[4:0]                    ), //i
    .io_dataOut   (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .dat2_i_clk   (dat2_i_clk                            ), //i
    .dat2_i_reset (dat2_i_reset                          )  //i
  );
  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_3 pushToPopGray_buffercc (
    .io_dataIn  (pushToPopGray[4:0]                    ), //i
    .io_dataOut (pushToPopGray_buffercc_io_dataOut[4:0]), //o
    .clk        (clk                                   ), //i
    .reset      (reset                                 )  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[127 : 0];
  assign popCC_readPort_rsp_mask = _zz_popCC_readPort_rsp_data[143 : 128];
  assign popCC_readPort_rsp_sink = _zz_popCC_readPort_rsp_data[147 : 144];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[148];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_mask = popCC_readPort_rsp_mask;
  assign popCC_readArbitation_translated_payload_sink = popCC_readPort_rsp_sink;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_mask = popCC_readArbitation_translated_payload_mask;
  assign io_pop_payload_sink = popCC_readArbitation_translated_payload_sink;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge dat2_i_clk) begin
    if(dat2_i_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module EfxDMA_BsbUpSizerDense_1 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [31:0]   io_input_payload_data,
  input  wire [3:0]    io_input_payload_mask,
  input  wire [3:0]    io_input_payload_sink,
  input  wire          io_input_payload_last,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [127:0]  io_output_payload_data,
  output wire [15:0]   io_output_payload_mask,
  output wire [3:0]    io_output_payload_sink,
  output wire          io_output_payload_last,
  input  wire          dat2_i_clk,
  input  wire          dat2_i_reset
);

  reg                 valid;
  reg        [1:0]    counter;
  reg        [127:0]  buffer_data;
  reg        [15:0]   buffer_mask;
  reg        [3:0]    buffer_sink;
  reg                 buffer_last;
  wire                full;
  wire                canAggregate;
  wire                onOutput;
  wire       [1:0]    counterSample;
  wire                io_output_fire;
  wire                io_input_fire;
  wire       [3:0]    _zz_1;
  wire       [3:0]    _zz_2;

  assign full = ((counter == 2'b00) || buffer_last);
  assign canAggregate = ((((valid && (! buffer_last)) && (! full)) && 1'b1) && (buffer_sink == io_input_payload_sink));
  assign counterSample = (canAggregate ? counter : 2'b00);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign _zz_1 = ({3'd0,1'b1} <<< counterSample);
  assign _zz_2 = ({3'd0,1'b1} <<< counterSample);
  assign io_output_valid = (valid && ((valid && full) || (io_input_valid && (! canAggregate))));
  assign io_output_payload_data = buffer_data;
  assign io_output_payload_mask = buffer_mask;
  assign io_output_payload_sink = buffer_sink;
  assign io_output_payload_last = buffer_last;
  assign io_input_ready = (((! valid) || canAggregate) || io_output_ready);
  always @(posedge dat2_i_clk) begin
    if(dat2_i_reset) begin
      valid <= 1'b0;
      counter <= 2'b00;
      buffer_last <= 1'b0;
      buffer_mask <= 16'h0;
    end else begin
      if(io_output_fire) begin
        valid <= 1'b0;
        buffer_mask <= 16'h0;
      end
      if(io_input_fire) begin
        valid <= 1'b1;
        if(_zz_2[0]) begin
          buffer_mask[3 : 0] <= io_input_payload_mask;
        end
        if(_zz_2[1]) begin
          buffer_mask[7 : 4] <= io_input_payload_mask;
        end
        if(_zz_2[2]) begin
          buffer_mask[11 : 8] <= io_input_payload_mask;
        end
        if(_zz_2[3]) begin
          buffer_mask[15 : 12] <= io_input_payload_mask;
        end
        buffer_last <= io_input_payload_last;
        counter <= (counterSample + 2'b01);
      end
    end
  end

  always @(posedge dat2_i_clk) begin
    if(io_input_fire) begin
      buffer_sink <= io_input_payload_sink;
      if(_zz_1[0]) begin
        buffer_data[31 : 0] <= io_input_payload_data;
      end
      if(_zz_1[1]) begin
        buffer_data[63 : 32] <= io_input_payload_data;
      end
      if(_zz_1[2]) begin
        buffer_data[95 : 64] <= io_input_payload_data;
      end
      if(_zz_1[3]) begin
        buffer_data[127 : 96] <= io_input_payload_data;
      end
    end
  end


endmodule

module EfxDMA_StreamFifoCC (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [127:0]  io_push_payload_data,
  input  wire [15:0]   io_push_payload_mask,
  input  wire [3:0]    io_push_payload_sink,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [127:0]  io_pop_payload_data,
  output wire [15:0]   io_pop_payload_mask,
  output wire [3:0]    io_pop_payload_sink,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          dat0_i_clk,
  input  wire          dat0_i_reset,
  input  wire          clk,
  input  wire          reset
);

  reg        [148:0]  ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [148:0]  _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [127:0]  popCC_readPort_rsp_data;
  wire       [15:0]   popCC_readPort_rsp_mask;
  wire       [3:0]    popCC_readPort_rsp_sink;
  wire                popCC_readPort_rsp_last;
  wire       [148:0]  _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [127:0]  popCC_readArbitation_translated_payload_data;
  wire       [15:0]   popCC_readArbitation_translated_payload_mask;
  wire       [3:0]    popCC_readArbitation_translated_payload_sink;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [148:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_sink,{io_push_payload_mask,io_push_payload_data}}};
  always @(posedge dat0_i_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_2 popToPushGray_buffercc (
    .io_dataIn    (popToPushGray[4:0]                    ), //i
    .io_dataOut   (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .dat0_i_clk   (dat0_i_clk                            ), //i
    .dat0_i_reset (dat0_i_reset                          )  //i
  );
  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_3 pushToPopGray_buffercc (
    .io_dataIn  (pushToPopGray[4:0]                    ), //i
    .io_dataOut (pushToPopGray_buffercc_io_dataOut[4:0]), //o
    .clk        (clk                                   ), //i
    .reset      (reset                                 )  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[127 : 0];
  assign popCC_readPort_rsp_mask = _zz_popCC_readPort_rsp_data[143 : 128];
  assign popCC_readPort_rsp_sink = _zz_popCC_readPort_rsp_data[147 : 144];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[148];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_mask = popCC_readPort_rsp_mask;
  assign popCC_readArbitation_translated_payload_sink = popCC_readPort_rsp_sink;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_mask = popCC_readArbitation_translated_payload_mask;
  assign io_pop_payload_sink = popCC_readArbitation_translated_payload_sink;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge dat0_i_clk) begin
    if(dat0_i_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module EfxDMA_BsbUpSizerDense (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [63:0]   io_input_payload_data,
  input  wire [7:0]    io_input_payload_mask,
  input  wire [3:0]    io_input_payload_sink,
  input  wire          io_input_payload_last,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [127:0]  io_output_payload_data,
  output wire [15:0]   io_output_payload_mask,
  output wire [3:0]    io_output_payload_sink,
  output wire          io_output_payload_last,
  input  wire          dat0_i_clk,
  input  wire          dat0_i_reset
);

  reg                 valid;
  reg        [0:0]    counter;
  reg        [127:0]  buffer_data;
  reg        [15:0]   buffer_mask;
  reg        [3:0]    buffer_sink;
  reg                 buffer_last;
  wire                full;
  wire                canAggregate;
  wire                onOutput;
  wire       [0:0]    counterSample;
  wire                io_output_fire;
  wire                io_input_fire;
  wire       [1:0]    _zz_1;
  wire       [1:0]    _zz_2;

  assign full = ((counter == 1'b0) || buffer_last);
  assign canAggregate = ((((valid && (! buffer_last)) && (! full)) && 1'b1) && (buffer_sink == io_input_payload_sink));
  assign counterSample = (canAggregate ? counter : 1'b0);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign _zz_1 = ({1'd0,1'b1} <<< counterSample);
  assign _zz_2 = ({1'd0,1'b1} <<< counterSample);
  assign io_output_valid = (valid && ((valid && full) || (io_input_valid && (! canAggregate))));
  assign io_output_payload_data = buffer_data;
  assign io_output_payload_mask = buffer_mask;
  assign io_output_payload_sink = buffer_sink;
  assign io_output_payload_last = buffer_last;
  assign io_input_ready = (((! valid) || canAggregate) || io_output_ready);
  always @(posedge dat0_i_clk) begin
    if(dat0_i_reset) begin
      valid <= 1'b0;
      counter <= 1'b0;
      buffer_last <= 1'b0;
      buffer_mask <= 16'h0;
    end else begin
      if(io_output_fire) begin
        valid <= 1'b0;
        buffer_mask <= 16'h0;
      end
      if(io_input_fire) begin
        valid <= 1'b1;
        if(_zz_2[0]) begin
          buffer_mask[7 : 0] <= io_input_payload_mask;
        end
        if(_zz_2[1]) begin
          buffer_mask[15 : 8] <= io_input_payload_mask;
        end
        buffer_last <= io_input_payload_last;
        counter <= (counterSample + 1'b1);
      end
    end
  end

  always @(posedge dat0_i_clk) begin
    if(io_input_fire) begin
      buffer_sink <= io_input_payload_sink;
      if(_zz_1[0]) begin
        buffer_data[63 : 0] <= io_input_payload_data;
      end
      if(_zz_1[1]) begin
        buffer_data[127 : 64] <= io_input_payload_data;
      end
    end
  end


endmodule

module EfxDMA_BmbToAxi4WriteOnlyBridge (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [12:0]   io_input_cmd_payload_fragment_length,
  input  wire [255:0]  io_input_cmd_payload_fragment_data,
  input  wire [31:0]   io_input_cmd_payload_fragment_mask,
  input  wire [15:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [15:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [7:0]    io_output_aw_payload_len,
  output wire [2:0]    io_output_aw_payload_size,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [255:0]  io_output_w_payload_data,
  output wire [31:0]   io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  reg                 contextRemover_io_output_cmd_ready;
  reg        [0:0]    contextRemover_io_output_rsp_payload_fragment_opcode;
  wire                contextRemover_io_input_cmd_ready;
  wire                contextRemover_io_input_rsp_valid;
  wire                contextRemover_io_input_rsp_payload_last;
  wire       [0:0]    contextRemover_io_input_rsp_payload_fragment_opcode;
  wire       [15:0]   contextRemover_io_input_rsp_payload_fragment_context;
  wire                contextRemover_io_output_cmd_valid;
  wire                contextRemover_io_output_cmd_payload_last;
  wire       [0:0]    contextRemover_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   contextRemover_io_output_cmd_payload_fragment_address;
  wire       [12:0]   contextRemover_io_output_cmd_payload_fragment_length;
  wire       [255:0]  contextRemover_io_output_cmd_payload_fragment_data;
  wire       [31:0]   contextRemover_io_output_cmd_payload_fragment_mask;
  wire                contextRemover_io_output_rsp_ready;
  wire       [8:0]    _zz_io_output_aw_payload_len;
  wire       [13:0]   _zz_io_output_aw_payload_len_1;
  wire       [13:0]   _zz_io_output_aw_payload_len_2;
  wire       [4:0]    _zz_io_output_aw_payload_len_3;
  wire                cmdFork_valid;
  reg                 cmdFork_ready;
  wire                cmdFork_payload_last;
  wire       [0:0]    cmdFork_payload_fragment_opcode;
  wire       [31:0]   cmdFork_payload_fragment_address;
  wire       [12:0]   cmdFork_payload_fragment_length;
  wire       [255:0]  cmdFork_payload_fragment_data;
  wire       [31:0]   cmdFork_payload_fragment_mask;
  wire                dataFork_valid;
  wire                dataFork_ready;
  wire                dataFork_payload_last;
  wire       [0:0]    dataFork_payload_fragment_opcode;
  wire       [31:0]   dataFork_payload_fragment_address;
  wire       [12:0]   dataFork_payload_fragment_length;
  wire       [255:0]  dataFork_payload_fragment_data;
  wire       [31:0]   dataFork_payload_fragment_mask;
  reg                 contextRemover_io_output_cmd_fork2_logic_linkEnable_0;
  reg                 contextRemover_io_output_cmd_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdFork_fire;
  wire                dataFork_fire;
  wire                contextRemover_io_output_cmd_fire;
  reg                 contextRemover_io_output_cmd_payload_first;
  wire                when_Stream_l445;
  reg                 cmdStage_valid;
  wire                cmdStage_ready;
  wire                cmdStage_payload_last;
  wire       [0:0]    cmdStage_payload_fragment_opcode;
  wire       [31:0]   cmdStage_payload_fragment_address;
  wire       [12:0]   cmdStage_payload_fragment_length;
  wire       [255:0]  cmdStage_payload_fragment_data;
  wire       [31:0]   cmdStage_payload_fragment_mask;
  wire                when_BmbToAxi4Bridge_l297;

  assign _zz_io_output_aw_payload_len = _zz_io_output_aw_payload_len_1[13 : 5];
  assign _zz_io_output_aw_payload_len_1 = ({1'b0,cmdStage_payload_fragment_length} + _zz_io_output_aw_payload_len_2);
  assign _zz_io_output_aw_payload_len_3 = cmdStage_payload_fragment_address[4 : 0];
  assign _zz_io_output_aw_payload_len_2 = {9'd0, _zz_io_output_aw_payload_len_3};
  EfxDMA_BmbContextRemover_1 contextRemover (
    .io_input_cmd_valid                     (io_input_cmd_valid                                         ), //i
    .io_input_cmd_ready                     (contextRemover_io_input_cmd_ready                          ), //o
    .io_input_cmd_payload_last              (io_input_cmd_payload_last                                  ), //i
    .io_input_cmd_payload_fragment_opcode   (io_input_cmd_payload_fragment_opcode                       ), //i
    .io_input_cmd_payload_fragment_address  (io_input_cmd_payload_fragment_address[31:0]                ), //i
    .io_input_cmd_payload_fragment_length   (io_input_cmd_payload_fragment_length[12:0]                 ), //i
    .io_input_cmd_payload_fragment_data     (io_input_cmd_payload_fragment_data[255:0]                  ), //i
    .io_input_cmd_payload_fragment_mask     (io_input_cmd_payload_fragment_mask[31:0]                   ), //i
    .io_input_cmd_payload_fragment_context  (io_input_cmd_payload_fragment_context[15:0]                ), //i
    .io_input_rsp_valid                     (contextRemover_io_input_rsp_valid                          ), //o
    .io_input_rsp_ready                     (io_input_rsp_ready                                         ), //i
    .io_input_rsp_payload_last              (contextRemover_io_input_rsp_payload_last                   ), //o
    .io_input_rsp_payload_fragment_opcode   (contextRemover_io_input_rsp_payload_fragment_opcode        ), //o
    .io_input_rsp_payload_fragment_context  (contextRemover_io_input_rsp_payload_fragment_context[15:0] ), //o
    .io_output_cmd_valid                    (contextRemover_io_output_cmd_valid                         ), //o
    .io_output_cmd_ready                    (contextRemover_io_output_cmd_ready                         ), //i
    .io_output_cmd_payload_last             (contextRemover_io_output_cmd_payload_last                  ), //o
    .io_output_cmd_payload_fragment_opcode  (contextRemover_io_output_cmd_payload_fragment_opcode       ), //o
    .io_output_cmd_payload_fragment_address (contextRemover_io_output_cmd_payload_fragment_address[31:0]), //o
    .io_output_cmd_payload_fragment_length  (contextRemover_io_output_cmd_payload_fragment_length[12:0] ), //o
    .io_output_cmd_payload_fragment_data    (contextRemover_io_output_cmd_payload_fragment_data[255:0]  ), //o
    .io_output_cmd_payload_fragment_mask    (contextRemover_io_output_cmd_payload_fragment_mask[31:0]   ), //o
    .io_output_rsp_valid                    (io_output_b_valid                                          ), //i
    .io_output_rsp_ready                    (contextRemover_io_output_rsp_ready                         ), //o
    .io_output_rsp_payload_last             (1'b1                                                       ), //i
    .io_output_rsp_payload_fragment_opcode  (contextRemover_io_output_rsp_payload_fragment_opcode       ), //i
    .clk                                    (clk                                                        ), //i
    .reset                                  (reset                                                      )  //i
  );
  assign io_input_cmd_ready = contextRemover_io_input_cmd_ready;
  assign io_input_rsp_valid = contextRemover_io_input_rsp_valid;
  assign io_input_rsp_payload_last = contextRemover_io_input_rsp_payload_last;
  assign io_input_rsp_payload_fragment_opcode = contextRemover_io_input_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_context = contextRemover_io_input_rsp_payload_fragment_context;
  always @(*) begin
    contextRemover_io_output_cmd_ready = 1'b1;
    if(when_Stream_l1063) begin
      contextRemover_io_output_cmd_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      contextRemover_io_output_cmd_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdFork_ready) && contextRemover_io_output_cmd_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! dataFork_ready) && contextRemover_io_output_cmd_fork2_logic_linkEnable_1);
  assign cmdFork_valid = (contextRemover_io_output_cmd_valid && contextRemover_io_output_cmd_fork2_logic_linkEnable_0);
  assign cmdFork_payload_last = contextRemover_io_output_cmd_payload_last;
  assign cmdFork_payload_fragment_opcode = contextRemover_io_output_cmd_payload_fragment_opcode;
  assign cmdFork_payload_fragment_address = contextRemover_io_output_cmd_payload_fragment_address;
  assign cmdFork_payload_fragment_length = contextRemover_io_output_cmd_payload_fragment_length;
  assign cmdFork_payload_fragment_data = contextRemover_io_output_cmd_payload_fragment_data;
  assign cmdFork_payload_fragment_mask = contextRemover_io_output_cmd_payload_fragment_mask;
  assign cmdFork_fire = (cmdFork_valid && cmdFork_ready);
  assign dataFork_valid = (contextRemover_io_output_cmd_valid && contextRemover_io_output_cmd_fork2_logic_linkEnable_1);
  assign dataFork_payload_last = contextRemover_io_output_cmd_payload_last;
  assign dataFork_payload_fragment_opcode = contextRemover_io_output_cmd_payload_fragment_opcode;
  assign dataFork_payload_fragment_address = contextRemover_io_output_cmd_payload_fragment_address;
  assign dataFork_payload_fragment_length = contextRemover_io_output_cmd_payload_fragment_length;
  assign dataFork_payload_fragment_data = contextRemover_io_output_cmd_payload_fragment_data;
  assign dataFork_payload_fragment_mask = contextRemover_io_output_cmd_payload_fragment_mask;
  assign dataFork_fire = (dataFork_valid && dataFork_ready);
  assign contextRemover_io_output_cmd_fire = (contextRemover_io_output_cmd_valid && contextRemover_io_output_cmd_ready);
  assign when_Stream_l445 = (! contextRemover_io_output_cmd_payload_first);
  always @(*) begin
    cmdStage_valid = cmdFork_valid;
    if(when_Stream_l445) begin
      cmdStage_valid = 1'b0;
    end
  end

  always @(*) begin
    cmdFork_ready = cmdStage_ready;
    if(when_Stream_l445) begin
      cmdFork_ready = 1'b1;
    end
  end

  assign cmdStage_payload_last = cmdFork_payload_last;
  assign cmdStage_payload_fragment_opcode = cmdFork_payload_fragment_opcode;
  assign cmdStage_payload_fragment_address = cmdFork_payload_fragment_address;
  assign cmdStage_payload_fragment_length = cmdFork_payload_fragment_length;
  assign cmdStage_payload_fragment_data = cmdFork_payload_fragment_data;
  assign cmdStage_payload_fragment_mask = cmdFork_payload_fragment_mask;
  assign io_output_aw_valid = cmdStage_valid;
  assign cmdStage_ready = io_output_aw_ready;
  assign io_output_aw_payload_addr = cmdStage_payload_fragment_address;
  assign io_output_aw_payload_len = _zz_io_output_aw_payload_len[7:0];
  assign io_output_aw_payload_size = 3'b101;
  assign io_output_aw_payload_prot = 3'b010;
  assign io_output_aw_payload_cache = 4'b1111;
  assign io_output_w_valid = dataFork_valid;
  assign dataFork_ready = io_output_w_ready;
  assign io_output_w_payload_data = dataFork_payload_fragment_data;
  assign io_output_w_payload_strb = dataFork_payload_fragment_mask;
  assign io_output_w_payload_last = dataFork_payload_last;
  assign io_output_b_ready = contextRemover_io_output_rsp_ready;
  assign when_BmbToAxi4Bridge_l297 = (io_output_b_payload_resp == 2'b00);
  always @(*) begin
    if(when_BmbToAxi4Bridge_l297) begin
      contextRemover_io_output_rsp_payload_fragment_opcode = 1'b0;
    end else begin
      contextRemover_io_output_rsp_payload_fragment_opcode = 1'b1;
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      contextRemover_io_output_cmd_fork2_logic_linkEnable_0 <= 1'b1;
      contextRemover_io_output_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      contextRemover_io_output_cmd_payload_first <= 1'b1;
    end else begin
      if(cmdFork_fire) begin
        contextRemover_io_output_cmd_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(dataFork_fire) begin
        contextRemover_io_output_cmd_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(contextRemover_io_output_cmd_ready) begin
        contextRemover_io_output_cmd_fork2_logic_linkEnable_0 <= 1'b1;
        contextRemover_io_output_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(contextRemover_io_output_cmd_fire) begin
        contextRemover_io_output_cmd_payload_first <= contextRemover_io_output_cmd_payload_last;
      end
    end
  end


endmodule

module EfxDMA_BmbSourceRemover_1 (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [12:0]   io_input_cmd_payload_fragment_length,
  input  wire [255:0]  io_input_cmd_payload_fragment_data,
  input  wire [31:0]   io_input_cmd_payload_fragment_mask,
  input  wire [14:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [14:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [12:0]   io_output_cmd_payload_fragment_length,
  output wire [255:0]  io_output_cmd_payload_fragment_data,
  output wire [31:0]   io_output_cmd_payload_fragment_mask,
  output wire [15:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [15:0]   io_output_rsp_payload_fragment_context
);

  wire       [0:0]    cmdContext_source;
  wire       [14:0]   cmdContext_context;
  wire       [0:0]    rspContext_source;
  wire       [14:0]   rspContext_context;
  wire       [15:0]   _zz_rspContext_source;

  assign cmdContext_source = io_input_cmd_payload_fragment_source;
  assign cmdContext_context = io_input_cmd_payload_fragment_context;
  assign io_output_cmd_valid = io_input_cmd_valid;
  assign io_input_cmd_ready = io_output_cmd_ready;
  assign io_output_cmd_payload_last = io_input_cmd_payload_last;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_output_cmd_payload_fragment_context = {cmdContext_context,cmdContext_source};
  assign _zz_rspContext_source = io_output_rsp_payload_fragment_context;
  assign rspContext_source = _zz_rspContext_source[0 : 0];
  assign rspContext_context = _zz_rspContext_source[15 : 1];
  assign io_input_rsp_valid = io_output_rsp_valid;
  assign io_output_rsp_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = io_output_rsp_payload_last;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_source = rspContext_source;
  assign io_input_rsp_payload_fragment_context = rspContext_context;

endmodule

module EfxDMA_BmbToAxi4ReadOnlyBridge (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [12:0]   io_input_cmd_payload_fragment_length,
  input  wire [25:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [255:0]  io_input_rsp_payload_fragment_data,
  output wire [25:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [7:0]    io_output_ar_payload_len,
  output wire [2:0]    io_output_ar_payload_size,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [255:0]  io_output_r_payload_data,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  reg        [0:0]    contextRemover_io_output_rsp_payload_fragment_opcode;
  wire                contextRemover_io_input_cmd_ready;
  wire                contextRemover_io_input_rsp_valid;
  wire                contextRemover_io_input_rsp_payload_last;
  wire       [0:0]    contextRemover_io_input_rsp_payload_fragment_opcode;
  wire       [255:0]  contextRemover_io_input_rsp_payload_fragment_data;
  wire       [25:0]   contextRemover_io_input_rsp_payload_fragment_context;
  wire                contextRemover_io_output_cmd_valid;
  wire                contextRemover_io_output_cmd_payload_last;
  wire       [0:0]    contextRemover_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   contextRemover_io_output_cmd_payload_fragment_address;
  wire       [12:0]   contextRemover_io_output_cmd_payload_fragment_length;
  wire                contextRemover_io_output_rsp_ready;
  wire       [8:0]    _zz_io_output_ar_payload_len;
  wire       [13:0]   _zz_io_output_ar_payload_len_1;
  wire       [13:0]   _zz_io_output_ar_payload_len_2;
  wire       [4:0]    _zz_io_output_ar_payload_len_3;
  wire                when_BmbToAxi4Bridge_l243;

  assign _zz_io_output_ar_payload_len = _zz_io_output_ar_payload_len_1[13 : 5];
  assign _zz_io_output_ar_payload_len_1 = ({1'b0,contextRemover_io_output_cmd_payload_fragment_length} + _zz_io_output_ar_payload_len_2);
  assign _zz_io_output_ar_payload_len_3 = contextRemover_io_output_cmd_payload_fragment_address[4 : 0];
  assign _zz_io_output_ar_payload_len_2 = {9'd0, _zz_io_output_ar_payload_len_3};
  EfxDMA_BmbContextRemover contextRemover (
    .io_input_cmd_valid                     (io_input_cmd_valid                                         ), //i
    .io_input_cmd_ready                     (contextRemover_io_input_cmd_ready                          ), //o
    .io_input_cmd_payload_last              (io_input_cmd_payload_last                                  ), //i
    .io_input_cmd_payload_fragment_opcode   (io_input_cmd_payload_fragment_opcode                       ), //i
    .io_input_cmd_payload_fragment_address  (io_input_cmd_payload_fragment_address[31:0]                ), //i
    .io_input_cmd_payload_fragment_length   (io_input_cmd_payload_fragment_length[12:0]                 ), //i
    .io_input_cmd_payload_fragment_context  (io_input_cmd_payload_fragment_context[25:0]                ), //i
    .io_input_rsp_valid                     (contextRemover_io_input_rsp_valid                          ), //o
    .io_input_rsp_ready                     (io_input_rsp_ready                                         ), //i
    .io_input_rsp_payload_last              (contextRemover_io_input_rsp_payload_last                   ), //o
    .io_input_rsp_payload_fragment_opcode   (contextRemover_io_input_rsp_payload_fragment_opcode        ), //o
    .io_input_rsp_payload_fragment_data     (contextRemover_io_input_rsp_payload_fragment_data[255:0]   ), //o
    .io_input_rsp_payload_fragment_context  (contextRemover_io_input_rsp_payload_fragment_context[25:0] ), //o
    .io_output_cmd_valid                    (contextRemover_io_output_cmd_valid                         ), //o
    .io_output_cmd_ready                    (io_output_ar_ready                                         ), //i
    .io_output_cmd_payload_last             (contextRemover_io_output_cmd_payload_last                  ), //o
    .io_output_cmd_payload_fragment_opcode  (contextRemover_io_output_cmd_payload_fragment_opcode       ), //o
    .io_output_cmd_payload_fragment_address (contextRemover_io_output_cmd_payload_fragment_address[31:0]), //o
    .io_output_cmd_payload_fragment_length  (contextRemover_io_output_cmd_payload_fragment_length[12:0] ), //o
    .io_output_rsp_valid                    (io_output_r_valid                                          ), //i
    .io_output_rsp_ready                    (contextRemover_io_output_rsp_ready                         ), //o
    .io_output_rsp_payload_last             (io_output_r_payload_last                                   ), //i
    .io_output_rsp_payload_fragment_opcode  (contextRemover_io_output_rsp_payload_fragment_opcode       ), //i
    .io_output_rsp_payload_fragment_data    (io_output_r_payload_data[255:0]                            ), //i
    .clk                                    (clk                                                        ), //i
    .reset                                  (reset                                                      )  //i
  );
  assign io_input_cmd_ready = contextRemover_io_input_cmd_ready;
  assign io_input_rsp_valid = contextRemover_io_input_rsp_valid;
  assign io_input_rsp_payload_last = contextRemover_io_input_rsp_payload_last;
  assign io_input_rsp_payload_fragment_opcode = contextRemover_io_input_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = contextRemover_io_input_rsp_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = contextRemover_io_input_rsp_payload_fragment_context;
  assign io_output_ar_valid = contextRemover_io_output_cmd_valid;
  assign io_output_ar_payload_addr = contextRemover_io_output_cmd_payload_fragment_address;
  assign io_output_ar_payload_len = _zz_io_output_ar_payload_len[7:0];
  assign io_output_ar_payload_size = 3'b101;
  assign io_output_ar_payload_prot = 3'b010;
  assign io_output_ar_payload_cache = 4'b1111;
  assign io_output_r_ready = contextRemover_io_output_rsp_ready;
  assign when_BmbToAxi4Bridge_l243 = (io_output_r_payload_resp == 2'b00);
  always @(*) begin
    if(when_BmbToAxi4Bridge_l243) begin
      contextRemover_io_output_rsp_payload_fragment_opcode = 1'b0;
    end else begin
      contextRemover_io_output_rsp_payload_fragment_opcode = 1'b1;
    end
  end


endmodule

module EfxDMA_BmbSourceRemover (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [12:0]   io_input_cmd_payload_fragment_length,
  input  wire [24:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [255:0]  io_input_rsp_payload_fragment_data,
  output wire [24:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [12:0]   io_output_cmd_payload_fragment_length,
  output wire [25:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [255:0]  io_output_rsp_payload_fragment_data,
  input  wire [25:0]   io_output_rsp_payload_fragment_context
);

  wire       [0:0]    cmdContext_source;
  wire       [24:0]   cmdContext_context;
  wire       [0:0]    rspContext_source;
  wire       [24:0]   rspContext_context;
  wire       [25:0]   _zz_rspContext_source;

  assign cmdContext_source = io_input_cmd_payload_fragment_source;
  assign cmdContext_context = io_input_cmd_payload_fragment_context;
  assign io_output_cmd_valid = io_input_cmd_valid;
  assign io_input_cmd_ready = io_output_cmd_ready;
  assign io_output_cmd_payload_last = io_input_cmd_payload_last;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_output_cmd_payload_fragment_context = {cmdContext_context,cmdContext_source};
  assign _zz_rspContext_source = io_output_rsp_payload_fragment_context;
  assign rspContext_source = _zz_rspContext_source[0 : 0];
  assign rspContext_context = _zz_rspContext_source[25 : 1];
  assign io_input_rsp_valid = io_output_rsp_valid;
  assign io_output_rsp_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = io_output_rsp_payload_last;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_input_rsp_payload_fragment_source = rspContext_source;
  assign io_input_rsp_payload_fragment_context = rspContext_context;

endmodule

module EfxDMA_BufferCC_10 (
  input  wire [3:0]    io_dataIn,
  output wire [3:0]    io_dataOut,
  input  wire          ctrl_clk,
  input  wire          ctrl_reset
);

  (* async_reg = "true" *) reg        [3:0]    buffers_0;
  (* async_reg = "true" *) reg        [3:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge ctrl_clk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

module EfxDMA_Apb3CC (
  input  wire [13:0]   io_input_PADDR,
  input  wire [0:0]    io_input_PSEL,
  input  wire          io_input_PENABLE,
  output wire          io_input_PREADY,
  input  wire          io_input_PWRITE,
  input  wire [31:0]   io_input_PWDATA,
  output wire [31:0]   io_input_PRDATA,
  output wire          io_input_PSLVERROR,
  output wire [13:0]   io_output_PADDR,
  output reg  [0:0]    io_output_PSEL,
  output reg           io_output_PENABLE,
  input  wire          io_output_PREADY,
  output wire          io_output_PWRITE,
  output wire [31:0]   io_output_PWDATA,
  input  wire [31:0]   io_output_PRDATA,
  input  wire          io_output_PSLVERROR,
  input  wire          ctrl_clk,
  input  wire          ctrl_reset,
  input  wire          clk,
  input  wire          reset
);

  wire                flowCCUnsafeByToggle_io_output_valid;
  wire       [13:0]   flowCCUnsafeByToggle_io_output_payload_PADDR;
  wire                flowCCUnsafeByToggle_io_output_payload_PWRITE;
  wire       [31:0]   flowCCUnsafeByToggle_io_output_payload_PWDATA;
  wire                flowCCUnsafeByToggle_1_io_output_valid;
  wire       [31:0]   flowCCUnsafeByToggle_1_io_output_payload_PRDATA;
  wire                flowCCUnsafeByToggle_1_io_output_payload_PSLVERROR;
  wire                inputLogic_inputCmd_valid;
  wire       [13:0]   inputLogic_inputCmd_payload_PADDR;
  wire                inputLogic_inputCmd_payload_PWRITE;
  wire       [31:0]   inputLogic_inputCmd_payload_PWDATA;
  wire                inputLogic_inputRsp_valid;
  wire       [31:0]   inputLogic_inputRsp_payload_PRDATA;
  wire                inputLogic_inputRsp_payload_PSLVERROR;
  reg                 inputLogic_state;
  wire                flowCCUnsafeByToggle_io_output_toStream_valid;
  reg                 flowCCUnsafeByToggle_io_output_toStream_ready;
  wire       [13:0]   flowCCUnsafeByToggle_io_output_toStream_payload_PADDR;
  wire                flowCCUnsafeByToggle_io_output_toStream_payload_PWRITE;
  wire       [31:0]   flowCCUnsafeByToggle_io_output_toStream_payload_PWDATA;
  wire                outputLogic_outputCmd_valid;
  reg                 outputLogic_outputCmd_ready;
  wire       [13:0]   outputLogic_outputCmd_payload_PADDR;
  wire                outputLogic_outputCmd_payload_PWRITE;
  wire       [31:0]   outputLogic_outputCmd_payload_PWDATA;
  reg                 flowCCUnsafeByToggle_io_output_toStream_rValid;
  wire                flowCCUnsafeByToggle_io_output_toStream_fire;
  (* async_reg = "true" *) reg        [13:0]   flowCCUnsafeByToggle_io_output_toStream_rData_PADDR;
  (* async_reg = "true" *) reg                 flowCCUnsafeByToggle_io_output_toStream_rData_PWRITE;
  (* async_reg = "true" *) reg        [31:0]   flowCCUnsafeByToggle_io_output_toStream_rData_PWDATA;
  wire                when_Stream_l375;
  reg                 outputLogic_state;
  wire                when_Apb3CCToggle_l81;
  wire                outputLogic_outputRsp_valid;
  wire       [31:0]   outputLogic_outputRsp_payload_PRDATA;
  wire                outputLogic_outputRsp_payload_PSLVERROR;
  wire                outputLogic_outputCmd_fire;

  EfxDMA_FlowCCUnsafeByToggle flowCCUnsafeByToggle (
    .io_input_valid           (inputLogic_inputCmd_valid                          ), //i
    .io_input_payload_PADDR   (inputLogic_inputCmd_payload_PADDR[13:0]            ), //i
    .io_input_payload_PWRITE  (inputLogic_inputCmd_payload_PWRITE                 ), //i
    .io_input_payload_PWDATA  (inputLogic_inputCmd_payload_PWDATA[31:0]           ), //i
    .io_output_valid          (flowCCUnsafeByToggle_io_output_valid               ), //o
    .io_output_payload_PADDR  (flowCCUnsafeByToggle_io_output_payload_PADDR[13:0] ), //o
    .io_output_payload_PWRITE (flowCCUnsafeByToggle_io_output_payload_PWRITE      ), //o
    .io_output_payload_PWDATA (flowCCUnsafeByToggle_io_output_payload_PWDATA[31:0]), //o
    .ctrl_clk                 (ctrl_clk                                           ), //i
    .ctrl_reset               (ctrl_reset                                         ), //i
    .clk                      (clk                                                ), //i
    .reset                    (reset                                              )  //i
  );
  EfxDMA_FlowCCUnsafeByToggle_1 flowCCUnsafeByToggle_1 (
    .io_input_valid              (outputLogic_outputRsp_valid                          ), //i
    .io_input_payload_PRDATA     (outputLogic_outputRsp_payload_PRDATA[31:0]           ), //i
    .io_input_payload_PSLVERROR  (outputLogic_outputRsp_payload_PSLVERROR              ), //i
    .io_output_valid             (flowCCUnsafeByToggle_1_io_output_valid               ), //o
    .io_output_payload_PRDATA    (flowCCUnsafeByToggle_1_io_output_payload_PRDATA[31:0]), //o
    .io_output_payload_PSLVERROR (flowCCUnsafeByToggle_1_io_output_payload_PSLVERROR   ), //o
    .clk                         (clk                                                  ), //i
    .reset                       (reset                                                ), //i
    .ctrl_clk                    (ctrl_clk                                             ), //i
    .ctrl_reset                  (ctrl_reset                                           )  //i
  );
  assign inputLogic_inputCmd_valid = ((io_input_PSEL[0] && io_input_PENABLE) && (! inputLogic_state));
  assign inputLogic_inputCmd_payload_PADDR = io_input_PADDR;
  assign inputLogic_inputCmd_payload_PWRITE = io_input_PWRITE;
  assign inputLogic_inputCmd_payload_PWDATA = io_input_PWDATA;
  assign io_input_PREADY = inputLogic_inputRsp_valid;
  assign io_input_PRDATA = inputLogic_inputRsp_payload_PRDATA;
  assign io_input_PSLVERROR = inputLogic_inputRsp_payload_PSLVERROR;
  assign flowCCUnsafeByToggle_io_output_toStream_valid = flowCCUnsafeByToggle_io_output_valid;
  assign flowCCUnsafeByToggle_io_output_toStream_payload_PADDR = flowCCUnsafeByToggle_io_output_payload_PADDR;
  assign flowCCUnsafeByToggle_io_output_toStream_payload_PWRITE = flowCCUnsafeByToggle_io_output_payload_PWRITE;
  assign flowCCUnsafeByToggle_io_output_toStream_payload_PWDATA = flowCCUnsafeByToggle_io_output_payload_PWDATA;
  assign flowCCUnsafeByToggle_io_output_toStream_fire = (flowCCUnsafeByToggle_io_output_toStream_valid && flowCCUnsafeByToggle_io_output_toStream_ready);
  always @(*) begin
    flowCCUnsafeByToggle_io_output_toStream_ready = outputLogic_outputCmd_ready;
    if(when_Stream_l375) begin
      flowCCUnsafeByToggle_io_output_toStream_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! outputLogic_outputCmd_valid);
  assign outputLogic_outputCmd_valid = flowCCUnsafeByToggle_io_output_toStream_rValid;
  assign outputLogic_outputCmd_payload_PADDR = flowCCUnsafeByToggle_io_output_toStream_rData_PADDR;
  assign outputLogic_outputCmd_payload_PWRITE = flowCCUnsafeByToggle_io_output_toStream_rData_PWRITE;
  assign outputLogic_outputCmd_payload_PWDATA = flowCCUnsafeByToggle_io_output_toStream_rData_PWDATA;
  always @(*) begin
    io_output_PENABLE = 1'b0;
    if(outputLogic_outputCmd_valid) begin
      if(when_Apb3CCToggle_l81) begin
        io_output_PENABLE = 1'b0;
      end else begin
        io_output_PENABLE = 1'b1;
      end
    end
  end

  always @(*) begin
    io_output_PSEL = 1'b0;
    if(outputLogic_outputCmd_valid) begin
      io_output_PSEL = 1'b1;
    end
  end

  assign io_output_PADDR = outputLogic_outputCmd_payload_PADDR;
  assign io_output_PWDATA = outputLogic_outputCmd_payload_PWDATA;
  assign io_output_PWRITE = outputLogic_outputCmd_payload_PWRITE;
  always @(*) begin
    outputLogic_outputCmd_ready = 1'b0;
    if(outputLogic_outputCmd_valid) begin
      if(!when_Apb3CCToggle_l81) begin
        if(io_output_PREADY) begin
          outputLogic_outputCmd_ready = 1'b1;
        end
      end
    end
  end

  assign when_Apb3CCToggle_l81 = (! outputLogic_state);
  assign outputLogic_outputCmd_fire = (outputLogic_outputCmd_valid && outputLogic_outputCmd_ready);
  assign outputLogic_outputRsp_valid = outputLogic_outputCmd_fire;
  assign outputLogic_outputRsp_payload_PRDATA = io_output_PRDATA;
  assign outputLogic_outputRsp_payload_PSLVERROR = io_output_PSLVERROR;
  assign inputLogic_inputRsp_valid = flowCCUnsafeByToggle_1_io_output_valid;
  assign inputLogic_inputRsp_payload_PRDATA = flowCCUnsafeByToggle_1_io_output_payload_PRDATA;
  assign inputLogic_inputRsp_payload_PSLVERROR = flowCCUnsafeByToggle_1_io_output_payload_PSLVERROR;
  always @(posedge ctrl_clk) begin
    if(ctrl_reset) begin
      inputLogic_state <= 1'b0;
    end else begin
      if(inputLogic_inputCmd_valid) begin
        inputLogic_state <= 1'b1;
      end
      if(inputLogic_inputRsp_valid) begin
        inputLogic_state <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      flowCCUnsafeByToggle_io_output_toStream_rValid <= 1'b0;
      outputLogic_state <= 1'b0;
    end else begin
      if(flowCCUnsafeByToggle_io_output_toStream_ready) begin
        flowCCUnsafeByToggle_io_output_toStream_rValid <= flowCCUnsafeByToggle_io_output_toStream_valid;
      end
      if(outputLogic_outputCmd_valid) begin
        if(when_Apb3CCToggle_l81) begin
          outputLogic_state <= 1'b1;
        end else begin
          if(io_output_PREADY) begin
            outputLogic_state <= 1'b0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    if(flowCCUnsafeByToggle_io_output_toStream_fire) begin
      flowCCUnsafeByToggle_io_output_toStream_rData_PADDR <= flowCCUnsafeByToggle_io_output_toStream_payload_PADDR;
      flowCCUnsafeByToggle_io_output_toStream_rData_PWRITE <= flowCCUnsafeByToggle_io_output_toStream_payload_PWRITE;
      flowCCUnsafeByToggle_io_output_toStream_rData_PWDATA <= flowCCUnsafeByToggle_io_output_toStream_payload_PWDATA;
    end
  end


endmodule

module EfxDMA_Core (
  output reg           io_read_cmd_valid,
  input  wire          io_read_cmd_ready,
  output wire          io_read_cmd_payload_last,
  output wire [0:0]    io_read_cmd_payload_fragment_source,
  output wire [0:0]    io_read_cmd_payload_fragment_opcode,
  output wire [31:0]   io_read_cmd_payload_fragment_address,
  output wire [12:0]   io_read_cmd_payload_fragment_length,
  output wire [24:0]   io_read_cmd_payload_fragment_context,
  input  wire          io_read_rsp_valid,
  output wire          io_read_rsp_ready,
  input  wire          io_read_rsp_payload_last,
  input  wire [0:0]    io_read_rsp_payload_fragment_source,
  input  wire [0:0]    io_read_rsp_payload_fragment_opcode,
  input  wire [255:0]  io_read_rsp_payload_fragment_data,
  input  wire [24:0]   io_read_rsp_payload_fragment_context,
  output wire          io_write_cmd_valid,
  input  wire          io_write_cmd_ready,
  output wire          io_write_cmd_payload_last,
  output wire [0:0]    io_write_cmd_payload_fragment_source,
  output wire [0:0]    io_write_cmd_payload_fragment_opcode,
  output wire [31:0]   io_write_cmd_payload_fragment_address,
  output wire [12:0]   io_write_cmd_payload_fragment_length,
  output wire [255:0]  io_write_cmd_payload_fragment_data,
  output wire [31:0]   io_write_cmd_payload_fragment_mask,
  output wire [14:0]   io_write_cmd_payload_fragment_context,
  input  wire          io_write_rsp_valid,
  output wire          io_write_rsp_ready,
  input  wire          io_write_rsp_payload_last,
  input  wire [0:0]    io_write_rsp_payload_fragment_source,
  input  wire [0:0]    io_write_rsp_payload_fragment_opcode,
  input  wire [14:0]   io_write_rsp_payload_fragment_context,
  output wire          io_outputs_0_valid,
  input  wire          io_outputs_0_ready,
  output wire [127:0]  io_outputs_0_payload_data,
  output wire [15:0]   io_outputs_0_payload_mask,
  output wire [3:0]    io_outputs_0_payload_sink,
  output wire          io_outputs_0_payload_last,
  output wire          io_outputs_1_valid,
  input  wire          io_outputs_1_ready,
  output wire [127:0]  io_outputs_1_payload_data,
  output wire [15:0]   io_outputs_1_payload_mask,
  output wire [3:0]    io_outputs_1_payload_sink,
  output wire          io_outputs_1_payload_last,
  input  wire          io_inputs_0_valid,
  output reg           io_inputs_0_ready,
  input  wire [127:0]  io_inputs_0_payload_data,
  input  wire [15:0]   io_inputs_0_payload_mask,
  input  wire [3:0]    io_inputs_0_payload_sink,
  input  wire          io_inputs_0_payload_last,
  input  wire          io_inputs_1_valid,
  output reg           io_inputs_1_ready,
  input  wire [127:0]  io_inputs_1_payload_data,
  input  wire [15:0]   io_inputs_1_payload_mask,
  input  wire [3:0]    io_inputs_1_payload_sink,
  input  wire          io_inputs_1_payload_last,
  output reg  [3:0]    io_interrupts,
  input  wire [13:0]   io_ctrl_PADDR,
  input  wire [0:0]    io_ctrl_PSEL,
  input  wire          io_ctrl_PENABLE,
  output wire          io_ctrl_PREADY,
  input  wire          io_ctrl_PWRITE,
  input  wire [31:0]   io_ctrl_PWDATA,
  output reg  [31:0]   io_ctrl_PRDATA,
  output wire          io_ctrl_PSLVERROR,
  input  wire          clk,
  input  wire          reset
);

  wire       [12:0]   memory_core_io_writes_0_cmd_payload_address;
  wire       [7:0]    memory_core_io_writes_0_cmd_payload_context;
  wire       [12:0]   memory_core_io_writes_1_cmd_payload_address;
  wire       [7:0]    memory_core_io_writes_1_cmd_payload_context;
  wire       [12:0]   memory_core_io_writes_2_cmd_payload_address;
  reg        [31:0]   memory_core_io_writes_2_cmd_payload_mask;
  wire       [8:0]    memory_core_io_writes_2_cmd_payload_context;
  wire                memory_core_io_reads_0_cmd_valid;
  wire       [12:0]   memory_core_io_reads_0_cmd_payload_address;
  wire       [2:0]    memory_core_io_reads_0_cmd_payload_context;
  wire                memory_core_io_reads_1_cmd_valid;
  wire       [12:0]   memory_core_io_reads_1_cmd_payload_address;
  wire       [2:0]    memory_core_io_reads_1_cmd_payload_context;
  wire       [12:0]   memory_core_io_reads_2_cmd_payload_address;
  wire       [14:0]   memory_core_io_reads_2_cmd_payload_context;
  wire       [31:0]   b2m_fsm_aggregate_engine_io_input_payload_mask;
  wire                b2m_fsm_aggregate_engine_io_flush;
  wire       [4:0]    b2m_fsm_aggregate_engine_io_offset;
  wire                memory_core_io_writes_0_cmd_ready;
  wire                memory_core_io_writes_0_rsp_valid;
  wire       [7:0]    memory_core_io_writes_0_rsp_payload_context;
  wire                memory_core_io_writes_1_cmd_ready;
  wire                memory_core_io_writes_1_rsp_valid;
  wire       [7:0]    memory_core_io_writes_1_rsp_payload_context;
  wire                memory_core_io_writes_2_cmd_ready;
  wire                memory_core_io_writes_2_rsp_valid;
  wire       [8:0]    memory_core_io_writes_2_rsp_payload_context;
  wire                memory_core_io_reads_0_cmd_ready;
  wire                memory_core_io_reads_0_rsp_valid;
  wire       [127:0]  memory_core_io_reads_0_rsp_payload_data;
  wire       [15:0]   memory_core_io_reads_0_rsp_payload_mask;
  wire       [2:0]    memory_core_io_reads_0_rsp_payload_context;
  wire                memory_core_io_reads_1_cmd_ready;
  wire                memory_core_io_reads_1_rsp_valid;
  wire       [127:0]  memory_core_io_reads_1_rsp_payload_data;
  wire       [15:0]   memory_core_io_reads_1_rsp_payload_mask;
  wire       [2:0]    memory_core_io_reads_1_rsp_payload_context;
  wire                memory_core_io_reads_2_cmd_ready;
  wire                memory_core_io_reads_2_rsp_valid;
  wire       [255:0]  memory_core_io_reads_2_rsp_payload_data;
  wire       [31:0]   memory_core_io_reads_2_rsp_payload_mask;
  wire       [14:0]   memory_core_io_reads_2_rsp_payload_context;
  wire                b2m_fsm_aggregate_engine_io_input_ready;
  wire       [255:0]  b2m_fsm_aggregate_engine_io_output_data;
  wire       [31:0]   b2m_fsm_aggregate_engine_io_output_mask;
  wire                b2m_fsm_aggregate_engine_io_output_consumed;
  wire       [4:0]    b2m_fsm_aggregate_engine_io_output_usedUntil;
  wire       [17:0]   _zz_channels_0_fifo_pop_withOverride_backupNext;
  wire       [17:0]   _zz_channels_0_fifo_pop_withOverride_exposed;
  wire       [26:0]   _zz_channels_0_pop_b2m_selfFlush;
  wire       [17:0]   _zz_channels_0_pop_b2m_request;
  wire       [13:0]   _zz_channels_0_pop_b2m_request_1;
  wire       [12:0]   _zz_channels_0_pop_b2m_request_2;
  wire       [3:0]    _zz_channels_0_pop_b2m_memPending;
  wire       [3:0]    _zz_channels_0_pop_b2m_memPending_1;
  wire       [0:0]    _zz_channels_0_pop_b2m_memPending_2;
  wire       [3:0]    _zz_channels_0_pop_b2m_memPending_3;
  wire       [0:0]    _zz_channels_0_pop_b2m_memPending_4;
  wire       [31:0]   _zz_channels_0_pop_b2m_address;
  wire       [31:0]   _zz_channels_0_pop_b2m_address_1;
  wire       [13:0]   _zz_channels_0_fifo_push_available;
  wire       [17:0]   _zz_channels_1_fifo_pop_withoutOverride_exposed;
  wire       [3:0]    _zz_channels_1_push_m2b_memPending;
  wire       [3:0]    _zz_channels_1_push_m2b_memPending_1;
  wire       [0:0]    _zz_channels_1_push_m2b_memPending_2;
  wire       [3:0]    _zz_channels_1_push_m2b_memPending_3;
  wire       [0:0]    _zz_channels_1_push_m2b_memPending_4;
  wire       [13:0]   _zz_channels_1_push_m2b_loadRequest;
  wire       [8:0]    _zz_channels_1_push_m2b_loadRequest_1;
  wire       [25:0]   _zz_when_DmaSg_l486;
  wire       [31:0]   _zz_channels_1_push_m2b_address;
  wire       [31:0]   _zz_channels_1_push_m2b_address_1;
  wire       [13:0]   _zz_channels_1_fifo_push_available;
  wire       [17:0]   _zz_channels_2_fifo_pop_withOverride_backupNext;
  wire       [17:0]   _zz_channels_2_fifo_pop_withOverride_exposed;
  wire       [26:0]   _zz_channels_2_pop_b2m_selfFlush;
  wire       [17:0]   _zz_channels_2_pop_b2m_request;
  wire       [13:0]   _zz_channels_2_pop_b2m_request_1;
  wire       [12:0]   _zz_channels_2_pop_b2m_request_2;
  wire       [3:0]    _zz_channels_2_pop_b2m_memPending;
  wire       [3:0]    _zz_channels_2_pop_b2m_memPending_1;
  wire       [0:0]    _zz_channels_2_pop_b2m_memPending_2;
  wire       [3:0]    _zz_channels_2_pop_b2m_memPending_3;
  wire       [0:0]    _zz_channels_2_pop_b2m_memPending_4;
  wire       [31:0]   _zz_channels_2_pop_b2m_address;
  wire       [31:0]   _zz_channels_2_pop_b2m_address_1;
  wire       [13:0]   _zz_channels_2_fifo_push_available;
  wire       [17:0]   _zz_channels_3_fifo_pop_withoutOverride_exposed;
  wire       [3:0]    _zz_channels_3_push_m2b_memPending;
  wire       [3:0]    _zz_channels_3_push_m2b_memPending_1;
  wire       [0:0]    _zz_channels_3_push_m2b_memPending_2;
  wire       [3:0]    _zz_channels_3_push_m2b_memPending_3;
  wire       [0:0]    _zz_channels_3_push_m2b_memPending_4;
  wire       [13:0]   _zz_channels_3_push_m2b_loadRequest;
  wire       [8:0]    _zz_channels_3_push_m2b_loadRequest_1;
  wire       [25:0]   _zz_when_DmaSg_l486_1;
  wire       [31:0]   _zz_channels_3_push_m2b_address;
  wire       [31:0]   _zz_channels_3_push_m2b_address_1;
  wire       [13:0]   _zz_channels_3_fifo_push_available;
  wire       [0:0]    _zz_s2b_0_cmd_firsts;
  wire       [4:0]    _zz_s2b_0_cmd_firsts_1;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_8;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_9;
  reg        [4:0]    _zz_s2b_0_cmd_byteCount_10;
  wire       [2:0]    _zz_s2b_0_cmd_byteCount_11;
  reg        [4:0]    _zz_s2b_0_cmd_byteCount_12;
  wire       [2:0]    _zz_s2b_0_cmd_byteCount_13;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_14;
  reg        [4:0]    _zz_s2b_0_cmd_byteCount_15;
  wire       [2:0]    _zz_s2b_0_cmd_byteCount_16;
  reg        [4:0]    _zz_s2b_0_cmd_byteCount_17;
  wire       [2:0]    _zz_s2b_0_cmd_byteCount_18;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_19;
  reg        [4:0]    _zz_s2b_0_cmd_byteCount_20;
  wire       [2:0]    _zz_s2b_0_cmd_byteCount_21;
  reg        [4:0]    _zz_s2b_0_cmd_byteCount_22;
  wire       [2:0]    _zz_s2b_0_cmd_byteCount_23;
  wire       [0:0]    _zz_s2b_0_cmd_byteCount_24;
  wire       [0:0]    _zz_s2b_1_cmd_firsts;
  wire       [4:0]    _zz_s2b_1_cmd_firsts_1;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_8;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_9;
  reg        [4:0]    _zz_s2b_1_cmd_byteCount_10;
  wire       [2:0]    _zz_s2b_1_cmd_byteCount_11;
  reg        [4:0]    _zz_s2b_1_cmd_byteCount_12;
  wire       [2:0]    _zz_s2b_1_cmd_byteCount_13;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_14;
  reg        [4:0]    _zz_s2b_1_cmd_byteCount_15;
  wire       [2:0]    _zz_s2b_1_cmd_byteCount_16;
  reg        [4:0]    _zz_s2b_1_cmd_byteCount_17;
  wire       [2:0]    _zz_s2b_1_cmd_byteCount_18;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_19;
  reg        [4:0]    _zz_s2b_1_cmd_byteCount_20;
  wire       [2:0]    _zz_s2b_1_cmd_byteCount_21;
  reg        [4:0]    _zz_s2b_1_cmd_byteCount_22;
  wire       [2:0]    _zz_s2b_1_cmd_byteCount_23;
  wire       [0:0]    _zz_s2b_1_cmd_byteCount_24;
  wire       [3:0]    _zz__zz_m2b_cmd_s0_priority_chosenOh_2;
  wire       [3:0]    _zz__zz_m2b_cmd_s0_priority_chosenOh_2_1;
  wire       [1:0]    _zz__zz_m2b_cmd_s0_priority_chosenOh_2_2;
  reg        [1:0]    _zz__zz_m2b_cmd_s0_priority_chosenOh_2_3;
  reg                 _zz_m2b_cmd_s0_priority_weightLast;
  reg        [31:0]   _zz_m2b_cmd_s0_address;
  reg        [25:0]   _zz_m2b_cmd_s0_bytesLeft;
  reg        [12:0]   _zz_m2b_cmd_s0_lengthHead;
  wire       [25:0]   _zz_m2b_cmd_s0_length;
  wire       [25:0]   _zz_m2b_cmd_s0_length_1;
  wire       [25:0]   _zz_m2b_cmd_s0_length_2;
  wire       [25:0]   _zz_m2b_cmd_s0_lastBurst;
  wire       [31:0]   _zz_m2b_cmd_s1_context_stop;
  wire       [31:0]   _zz_m2b_cmd_s1_context_stop_1;
  wire       [31:0]   _zz_m2b_cmd_s1_addressNext;
  wire       [31:0]   _zz_m2b_cmd_s1_addressNext_1;
  wire       [25:0]   _zz_m2b_cmd_s1_byteLeftNext;
  wire       [25:0]   _zz_m2b_cmd_s1_byteLeftNext_1;
  wire       [13:0]   _zz_m2b_cmd_s1_fifoPushDecr;
  wire       [12:0]   _zz_m2b_cmd_s1_fifoPushDecr_1;
  wire       [12:0]   _zz_m2b_cmd_s1_fifoPushDecr_2;
  wire       [4:0]    _zz_m2b_cmd_s1_fifoPushDecr_3;
  wire       [13:0]   _zz_m2b_cmd_s1_fifoPushDecr_4;
  wire       [1:0]    _zz_m2b_cmd_s1_fifoPushDecr_5;
  reg        [13:0]   _zz_io_writes_2_cmd_payload_address;
  wire       [3:0]    _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2;
  wire       [3:0]    _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_1;
  wire       [1:0]    _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_2;
  reg        [1:0]    _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_3;
  reg                 _zz_b2m_fsm_arbiter_logic_priority_weightLast;
  reg        [31:0]   _zz_b2m_fsm_sel_address;
  reg        [13:0]   _zz_b2m_fsm_sel_ptr;
  reg        [13:0]   _zz_b2m_fsm_sel_ptrMask;
  reg        [12:0]   _zz_b2m_fsm_sel_bytePerBurst;
  reg        [17:0]   _zz_b2m_fsm_sel_bytesInFifo;
  reg                 _zz_b2m_fsm_sel_flush;
  reg                 _zz_b2m_fsm_sel_packet;
  reg        [26:0]   _zz_b2m_fsm_sel_bytesLeft;
  wire       [13:0]   _zz_b2m_fsm_bytesInBurstP1;
  wire       [1:0]    _zz_b2m_fsm_bytesInBurstP1_1;
  wire       [31:0]   _zz_b2m_fsm_addressNext;
  wire       [26:0]   _zz_b2m_fsm_bytesLeftNext;
  wire       [14:0]   _zz_b2m_fsm_bytesLeftNext_1;
  wire       [25:0]   _zz__zz_b2m_fsm_sel_bytesInBurst_1;
  wire       [25:0]   _zz__zz_b2m_fsm_sel_bytesInBurst_1_1;
  wire       [12:0]   _zz__zz_b2m_fsm_sel_bytesInBurst_2;
  wire       [25:0]   _zz_b2m_fsm_sel_bytesInBurst_3;
  wire       [25:0]   _zz_b2m_fsm_sel_bytesInBurst_4;
  wire       [25:0]   _zz_b2m_fsm_sel_bytesInBurst_5;
  wire       [17:0]   _zz_b2m_fsm_fifoCompletion;
  wire       [17:0]   _zz_b2m_fsm_fifoCompletion_1;
  wire       [12:0]   _zz_b2m_fsm_beatCounter;
  wire       [12:0]   _zz_b2m_fsm_beatCounter_1;
  wire       [4:0]    _zz_b2m_fsm_beatCounter_2;
  reg        [13:0]   _zz_b2m_fsm_fetch_context_ptr;
  wire       [13:0]   _zz_b2m_fsm_sel_ptr_1;
  reg        [4:0]    _zz_b2m_fsm_aggregate_bytesToSkip;
  wire       [4:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_1;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_2;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_3;
  wire       [0:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_4;
  wire       [25:0]   _zz_b2m_fsm_aggregate_bytesToSkipMask_5;
  wire       [4:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_6;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_7;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_8;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_9;
  wire       [0:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_10;
  wire       [19:0]   _zz_b2m_fsm_aggregate_bytesToSkipMask_11;
  wire       [4:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_12;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_13;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_14;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_15;
  wire       [0:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_16;
  wire       [13:0]   _zz_b2m_fsm_aggregate_bytesToSkipMask_17;
  wire       [4:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_18;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_19;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_20;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_21;
  wire       [0:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_22;
  wire       [7:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_23;
  wire       [4:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_24;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_25;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_26;
  wire                _zz_b2m_fsm_aggregate_bytesToSkipMask_27;
  wire       [0:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_28;
  wire       [1:0]    _zz_b2m_fsm_aggregate_bytesToSkipMask_29;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskLastTriggerComb;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskLast;
  wire                _zz_b2m_fsm_cmd_maskLast_1;
  wire       [0:0]    _zz_b2m_fsm_cmd_maskLast_2;
  wire       [23:0]   _zz_b2m_fsm_cmd_maskLast_3;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskLast_4;
  wire                _zz_b2m_fsm_cmd_maskLast_5;
  wire       [0:0]    _zz_b2m_fsm_cmd_maskLast_6;
  wire       [15:0]   _zz_b2m_fsm_cmd_maskLast_7;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskLast_8;
  wire                _zz_b2m_fsm_cmd_maskLast_9;
  wire       [0:0]    _zz_b2m_fsm_cmd_maskLast_10;
  wire       [7:0]    _zz_b2m_fsm_cmd_maskLast_11;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskLast_12;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskLast_13;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskFirst;
  wire                _zz_b2m_fsm_cmd_maskFirst_1;
  wire       [0:0]    _zz_b2m_fsm_cmd_maskFirst_2;
  wire       [23:0]   _zz_b2m_fsm_cmd_maskFirst_3;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskFirst_4;
  wire                _zz_b2m_fsm_cmd_maskFirst_5;
  wire       [0:0]    _zz_b2m_fsm_cmd_maskFirst_6;
  wire       [15:0]   _zz_b2m_fsm_cmd_maskFirst_7;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskFirst_8;
  wire                _zz_b2m_fsm_cmd_maskFirst_9;
  wire       [0:0]    _zz_b2m_fsm_cmd_maskFirst_10;
  wire       [7:0]    _zz_b2m_fsm_cmd_maskFirst_11;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskFirst_12;
  wire       [4:0]    _zz_b2m_fsm_cmd_maskFirst_13;
  wire       [0:0]    _zz_channels_0_channelStart;
  wire       [0:0]    _zz_channels_0_ctrl_kick;
  wire       [0:0]    _zz_channels_0_interrupts_completion_valid;
  wire       [0:0]    _zz_channels_0_interrupts_onChannelCompletion_valid;
  wire       [0:0]    _zz_channels_0_interrupts_s2mPacket_valid;
  wire       [0:0]    _zz_channels_1_channelStart;
  wire       [0:0]    _zz_channels_1_ctrl_kick;
  wire       [0:0]    _zz_channels_1_interrupts_completion_valid;
  wire       [0:0]    _zz_channels_1_interrupts_onChannelCompletion_valid;
  wire       [0:0]    _zz_channels_2_channelStart;
  wire       [0:0]    _zz_channels_2_ctrl_kick;
  wire       [0:0]    _zz_channels_2_interrupts_completion_valid;
  wire       [0:0]    _zz_channels_2_interrupts_onChannelCompletion_valid;
  wire       [0:0]    _zz_channels_2_interrupts_s2mPacket_valid;
  wire       [0:0]    _zz_channels_3_channelStart;
  wire       [0:0]    _zz_channels_3_ctrl_kick;
  wire       [0:0]    _zz_channels_3_interrupts_completion_valid;
  wire       [0:0]    _zz_channels_3_interrupts_onChannelCompletion_valid;
  wire       [13:0]   _zz_channels_0_fifo_push_ptrIncr_value;
  wire       [0:0]    _zz_channels_0_fifo_push_ptrIncr_value_1;
  wire       [17:0]   _zz_channels_0_fifo_pop_bytesIncr_value_1;
  wire       [4:0]    _zz_channels_0_fifo_pop_bytesIncr_value_2;
  wire       [13:0]   _zz_channels_0_fifo_pop_ptrIncr_value;
  wire       [1:0]    _zz_channels_0_fifo_pop_ptrIncr_value_1;
  wire       [13:0]   _zz_channels_1_fifo_push_ptrIncr_value;
  wire       [1:0]    _zz_channels_1_fifo_push_ptrIncr_value_1;
  wire       [17:0]   _zz_channels_1_fifo_pop_bytesIncr_value_1;
  wire       [5:0]    _zz_channels_1_fifo_pop_bytesIncr_value_2;
  wire       [5:0]    _zz_channels_1_fifo_pop_bytesIncr_value_3;
  wire       [13:0]   _zz_channels_1_fifo_pop_ptrIncr_value;
  wire       [0:0]    _zz_channels_1_fifo_pop_ptrIncr_value_1;
  wire       [13:0]   _zz_channels_2_fifo_push_ptrIncr_value;
  wire       [0:0]    _zz_channels_2_fifo_push_ptrIncr_value_1;
  wire       [17:0]   _zz_channels_2_fifo_pop_bytesIncr_value_1;
  wire       [4:0]    _zz_channels_2_fifo_pop_bytesIncr_value_2;
  wire       [13:0]   _zz_channels_2_fifo_pop_ptrIncr_value;
  wire       [1:0]    _zz_channels_2_fifo_pop_ptrIncr_value_1;
  wire       [13:0]   _zz_channels_3_fifo_push_ptrIncr_value;
  wire       [1:0]    _zz_channels_3_fifo_push_ptrIncr_value_1;
  wire       [17:0]   _zz_channels_3_fifo_pop_bytesIncr_value_1;
  wire       [5:0]    _zz_channels_3_fifo_pop_bytesIncr_value_2;
  wire       [5:0]    _zz_channels_3_fifo_pop_bytesIncr_value_3;
  wire       [13:0]   _zz_channels_3_fifo_pop_ptrIncr_value;
  wire       [0:0]    _zz_channels_3_fifo_pop_ptrIncr_value_1;
  wire                ctrl_readErrorFlag;
  wire                ctrl_writeErrorFlag;
  wire                ctrl_askWrite;
  wire                ctrl_askRead;
  wire                ctrl_doWrite;
  wire                ctrl_doRead;
  reg                 channels_0_channelStart;
  reg                 channels_0_channelStop;
  reg                 channels_0_channelCompletion;
  reg                 channels_0_channelValid;
  reg                 channels_0_descriptorStart;
  reg                 channels_0_descriptorCompletion;
  reg                 channels_0_descriptorValid;
  reg        [25:0]   channels_0_bytes;
  reg        [1:0]    channels_0_priority;
  reg        [1:0]    channels_0_weight;
  reg                 channels_0_selfRestart;
  reg                 channels_0_readyToStop;
  reg                 channels_0_ctrl_kick;
  wire       [13:0]   channels_0_fifo_base;
  wire       [13:0]   channels_0_fifo_words;
  reg        [13:0]   channels_0_fifo_push_available;
  wire       [13:0]   channels_0_fifo_push_availableDecr;
  reg        [13:0]   channels_0_fifo_push_ptr;
  wire       [13:0]   channels_0_fifo_push_ptrWithBase;
  wire       [13:0]   channels_0_fifo_push_ptrIncr_value;
  reg        [13:0]   channels_0_fifo_pop_ptr;
  wire       [17:0]   channels_0_fifo_pop_bytes;
  wire       [13:0]   channels_0_fifo_pop_ptrWithBase;
  wire       [17:0]   channels_0_fifo_pop_bytesIncr_value;
  wire       [17:0]   channels_0_fifo_pop_bytesDecr_value;
  wire                channels_0_fifo_pop_empty;
  wire       [13:0]   channels_0_fifo_pop_ptrIncr_value;
  reg        [17:0]   channels_0_fifo_pop_withOverride_backup;
  wire       [17:0]   channels_0_fifo_pop_withOverride_backupNext;
  reg                 channels_0_fifo_pop_withOverride_load;
  reg                 channels_0_fifo_pop_withOverride_unload;
  reg        [17:0]   channels_0_fifo_pop_withOverride_exposed;
  reg                 channels_0_fifo_pop_withOverride_valid;
  wire                when_DmaSg_l409;
  wire                channels_0_fifo_empty;
  reg                 channels_0_push_memory;
  reg                 channels_0_push_s2b_completionOnLast;
  reg                 channels_0_push_s2b_packetEvent;
  reg                 channels_0_push_s2b_packetLock;
  reg                 channels_0_push_s2b_waitFirst;
  wire                when_DmaSg_l457;
  reg                 channels_0_pop_memory;
  wire       [12:0]   channels_0_pop_b2m_bytePerBurst;
  reg                 channels_0_pop_b2m_fire;
  reg                 channels_0_pop_b2m_waitFinalRsp;
  reg                 channels_0_pop_b2m_flush;
  reg                 channels_0_pop_b2m_packetSync;
  reg                 channels_0_pop_b2m_packet;
  wire                when_DmaSg_l505;
  reg                 channels_0_pop_b2m_memRsp;
  reg        [3:0]    channels_0_pop_b2m_memPending;
  reg        [31:0]   channels_0_pop_b2m_address;
  reg        [26:0]   channels_0_pop_b2m_bytesLeft;
  wire                channels_0_pop_b2m_selfFlush;
  wire                channels_0_pop_b2m_request;
  reg        [4:0]    channels_0_pop_b2m_bytesToSkip;
  reg        [17:0]   channels_0_pop_b2m_decrBytes;
  reg                 channels_0_pop_b2m_memPendingInc;
  wire                when_DmaSg_l523;
  wire                when_DmaSg_l532;
  wire                when_DmaSg_l547;
  wire                when_DmaSg_l563;
  wire                channels_0_readyForChannelCompletion;
  wire                when_DmaSg_l575;
  reg                 _zz_when_DmaSg_l593;
  wire                when_DmaSg_l578;
  wire                when_DmaSg_l593;
  wire                channels_0_s2b_full;
  reg        [13:0]   channels_0_fifo_pop_ptrIncr_value_regNext;
  wire                when_DmaSg_l255;
  reg                 channels_0_interrupts_completion_enable;
  reg                 channels_0_interrupts_completion_valid;
  wire                when_DmaSg_l255_1;
  wire                when_DmaSg_l255_2;
  reg                 channels_0_interrupts_onChannelCompletion_enable;
  reg                 channels_0_interrupts_onChannelCompletion_valid;
  wire                when_DmaSg_l255_3;
  reg                 channels_0_interrupts_s2mPacket_enable;
  reg                 channels_0_interrupts_s2mPacket_valid;
  wire                when_DmaSg_l255_4;
  reg                 channels_1_channelStart;
  reg                 channels_1_channelStop;
  reg                 channels_1_channelCompletion;
  reg                 channels_1_channelValid;
  reg                 channels_1_descriptorStart;
  reg                 channels_1_descriptorCompletion;
  reg                 channels_1_descriptorValid;
  reg        [25:0]   channels_1_bytes;
  reg        [1:0]    channels_1_priority;
  reg        [1:0]    channels_1_weight;
  reg                 channels_1_selfRestart;
  reg                 channels_1_readyToStop;
  reg                 channels_1_ctrl_kick;
  wire       [13:0]   channels_1_fifo_base;
  wire       [13:0]   channels_1_fifo_words;
  reg        [13:0]   channels_1_fifo_push_available;
  reg        [13:0]   channels_1_fifo_push_availableDecr;
  reg        [13:0]   channels_1_fifo_push_ptr;
  wire       [13:0]   channels_1_fifo_push_ptrWithBase;
  wire       [13:0]   channels_1_fifo_push_ptrIncr_value;
  reg        [13:0]   channels_1_fifo_pop_ptr;
  wire       [17:0]   channels_1_fifo_pop_bytes;
  wire       [13:0]   channels_1_fifo_pop_ptrWithBase;
  wire       [17:0]   channels_1_fifo_pop_bytesIncr_value;
  wire       [17:0]   channels_1_fifo_pop_bytesDecr_value;
  wire                channels_1_fifo_pop_empty;
  wire       [13:0]   channels_1_fifo_pop_ptrIncr_value;
  reg        [17:0]   channels_1_fifo_pop_withoutOverride_exposed;
  wire                channels_1_fifo_empty;
  reg                 channels_1_push_memory;
  reg        [31:0]   channels_1_push_m2b_address;
  wire       [12:0]   channels_1_push_m2b_bytePerBurst;
  reg                 channels_1_push_m2b_loadDone;
  reg        [25:0]   channels_1_push_m2b_bytesLeft;
  reg        [3:0]    channels_1_push_m2b_memPending;
  reg                 channels_1_push_m2b_memPendingIncr;
  reg                 channels_1_push_m2b_memPendingDecr;
  reg                 channels_1_push_m2b_loadRequest;
  reg                 channels_1_pop_memory;
  reg                 channels_1_pop_b2s_last;
  reg        [0:0]    channels_1_pop_b2s_portId;
  reg        [3:0]    channels_1_pop_b2s_sinkId;
  reg                 channels_1_pop_b2s_veryLastTrigger;
  reg                 channels_1_pop_b2s_veryLastValid;
  wire                when_DmaSg_l474;
  reg        [13:0]   channels_1_pop_b2s_veryLastPtr;
  reg                 channels_1_pop_b2s_veryLastEndPacket;
  wire                when_DmaSg_l483;
  wire                when_DmaSg_l486;
  wire                when_DmaSg_l562;
  reg                 channels_1_readyForChannelCompletion;
  wire                when_DmaSg_l566;
  wire                when_DmaSg_l575_1;
  reg                 _zz_when_DmaSg_l593_1;
  wire                when_DmaSg_l578_1;
  wire                when_DmaSg_l593_1;
  wire                channels_1_s2b_full;
  reg        [13:0]   channels_1_fifo_pop_ptrIncr_value_regNext;
  wire                when_DmaSg_l255_5;
  reg                 channels_1_interrupts_completion_enable;
  reg                 channels_1_interrupts_completion_valid;
  wire                when_DmaSg_l255_6;
  wire                when_DmaSg_l255_7;
  reg                 channels_1_interrupts_onChannelCompletion_enable;
  reg                 channels_1_interrupts_onChannelCompletion_valid;
  wire                when_DmaSg_l255_8;
  reg                 channels_2_channelStart;
  reg                 channels_2_channelStop;
  reg                 channels_2_channelCompletion;
  reg                 channels_2_channelValid;
  reg                 channels_2_descriptorStart;
  reg                 channels_2_descriptorCompletion;
  reg                 channels_2_descriptorValid;
  reg        [25:0]   channels_2_bytes;
  reg        [1:0]    channels_2_priority;
  reg        [1:0]    channels_2_weight;
  reg                 channels_2_selfRestart;
  reg                 channels_2_readyToStop;
  reg                 channels_2_ctrl_kick;
  wire       [13:0]   channels_2_fifo_base;
  wire       [13:0]   channels_2_fifo_words;
  reg        [13:0]   channels_2_fifo_push_available;
  wire       [13:0]   channels_2_fifo_push_availableDecr;
  reg        [13:0]   channels_2_fifo_push_ptr;
  wire       [13:0]   channels_2_fifo_push_ptrWithBase;
  wire       [13:0]   channels_2_fifo_push_ptrIncr_value;
  reg        [13:0]   channels_2_fifo_pop_ptr;
  wire       [17:0]   channels_2_fifo_pop_bytes;
  wire       [13:0]   channels_2_fifo_pop_ptrWithBase;
  wire       [17:0]   channels_2_fifo_pop_bytesIncr_value;
  wire       [17:0]   channels_2_fifo_pop_bytesDecr_value;
  wire                channels_2_fifo_pop_empty;
  wire       [13:0]   channels_2_fifo_pop_ptrIncr_value;
  reg        [17:0]   channels_2_fifo_pop_withOverride_backup;
  wire       [17:0]   channels_2_fifo_pop_withOverride_backupNext;
  reg                 channels_2_fifo_pop_withOverride_load;
  reg                 channels_2_fifo_pop_withOverride_unload;
  reg        [17:0]   channels_2_fifo_pop_withOverride_exposed;
  reg                 channels_2_fifo_pop_withOverride_valid;
  wire                when_DmaSg_l409_1;
  wire                channels_2_fifo_empty;
  reg                 channels_2_push_memory;
  reg                 channels_2_push_s2b_completionOnLast;
  reg                 channels_2_push_s2b_packetEvent;
  reg                 channels_2_push_s2b_packetLock;
  reg                 channels_2_push_s2b_waitFirst;
  wire                when_DmaSg_l457_1;
  reg                 channels_2_pop_memory;
  wire       [12:0]   channels_2_pop_b2m_bytePerBurst;
  reg                 channels_2_pop_b2m_fire;
  reg                 channels_2_pop_b2m_waitFinalRsp;
  reg                 channels_2_pop_b2m_flush;
  reg                 channels_2_pop_b2m_packetSync;
  reg                 channels_2_pop_b2m_packet;
  wire                when_DmaSg_l505_1;
  reg                 channels_2_pop_b2m_memRsp;
  reg        [3:0]    channels_2_pop_b2m_memPending;
  reg        [31:0]   channels_2_pop_b2m_address;
  reg        [26:0]   channels_2_pop_b2m_bytesLeft;
  wire                channels_2_pop_b2m_selfFlush;
  wire                channels_2_pop_b2m_request;
  reg        [4:0]    channels_2_pop_b2m_bytesToSkip;
  reg        [17:0]   channels_2_pop_b2m_decrBytes;
  reg                 channels_2_pop_b2m_memPendingInc;
  wire                when_DmaSg_l523_1;
  wire                when_DmaSg_l532_1;
  wire                when_DmaSg_l547_1;
  wire                when_DmaSg_l563_1;
  wire                channels_2_readyForChannelCompletion;
  wire                when_DmaSg_l575_2;
  reg                 _zz_when_DmaSg_l593_2;
  wire                when_DmaSg_l578_2;
  wire                when_DmaSg_l593_2;
  wire                channels_2_s2b_full;
  reg        [13:0]   channels_2_fifo_pop_ptrIncr_value_regNext;
  wire                when_DmaSg_l255_9;
  reg                 channels_2_interrupts_completion_enable;
  reg                 channels_2_interrupts_completion_valid;
  wire                when_DmaSg_l255_10;
  wire                when_DmaSg_l255_11;
  reg                 channels_2_interrupts_onChannelCompletion_enable;
  reg                 channels_2_interrupts_onChannelCompletion_valid;
  wire                when_DmaSg_l255_12;
  reg                 channels_2_interrupts_s2mPacket_enable;
  reg                 channels_2_interrupts_s2mPacket_valid;
  wire                when_DmaSg_l255_13;
  reg                 channels_3_channelStart;
  reg                 channels_3_channelStop;
  reg                 channels_3_channelCompletion;
  reg                 channels_3_channelValid;
  reg                 channels_3_descriptorStart;
  reg                 channels_3_descriptorCompletion;
  reg                 channels_3_descriptorValid;
  reg        [25:0]   channels_3_bytes;
  reg        [1:0]    channels_3_priority;
  reg        [1:0]    channels_3_weight;
  reg                 channels_3_selfRestart;
  reg                 channels_3_readyToStop;
  reg                 channels_3_ctrl_kick;
  wire       [13:0]   channels_3_fifo_base;
  wire       [13:0]   channels_3_fifo_words;
  reg        [13:0]   channels_3_fifo_push_available;
  reg        [13:0]   channels_3_fifo_push_availableDecr;
  reg        [13:0]   channels_3_fifo_push_ptr;
  wire       [13:0]   channels_3_fifo_push_ptrWithBase;
  wire       [13:0]   channels_3_fifo_push_ptrIncr_value;
  reg        [13:0]   channels_3_fifo_pop_ptr;
  wire       [17:0]   channels_3_fifo_pop_bytes;
  wire       [13:0]   channels_3_fifo_pop_ptrWithBase;
  wire       [17:0]   channels_3_fifo_pop_bytesIncr_value;
  wire       [17:0]   channels_3_fifo_pop_bytesDecr_value;
  wire                channels_3_fifo_pop_empty;
  wire       [13:0]   channels_3_fifo_pop_ptrIncr_value;
  reg        [17:0]   channels_3_fifo_pop_withoutOverride_exposed;
  wire                channels_3_fifo_empty;
  reg                 channels_3_push_memory;
  reg        [31:0]   channels_3_push_m2b_address;
  wire       [12:0]   channels_3_push_m2b_bytePerBurst;
  reg                 channels_3_push_m2b_loadDone;
  reg        [25:0]   channels_3_push_m2b_bytesLeft;
  reg        [3:0]    channels_3_push_m2b_memPending;
  reg                 channels_3_push_m2b_memPendingIncr;
  reg                 channels_3_push_m2b_memPendingDecr;
  reg                 channels_3_push_m2b_loadRequest;
  reg                 channels_3_pop_memory;
  reg                 channels_3_pop_b2s_last;
  reg        [0:0]    channels_3_pop_b2s_portId;
  reg        [3:0]    channels_3_pop_b2s_sinkId;
  reg                 channels_3_pop_b2s_veryLastTrigger;
  reg                 channels_3_pop_b2s_veryLastValid;
  wire                when_DmaSg_l474_1;
  reg        [13:0]   channels_3_pop_b2s_veryLastPtr;
  reg                 channels_3_pop_b2s_veryLastEndPacket;
  wire                when_DmaSg_l483_1;
  wire                when_DmaSg_l486_1;
  wire                when_DmaSg_l562_1;
  reg                 channels_3_readyForChannelCompletion;
  wire                when_DmaSg_l566_1;
  wire                when_DmaSg_l575_3;
  reg                 _zz_when_DmaSg_l593_3;
  wire                when_DmaSg_l578_3;
  wire                when_DmaSg_l593_3;
  wire                channels_3_s2b_full;
  reg        [13:0]   channels_3_fifo_pop_ptrIncr_value_regNext;
  wire                when_DmaSg_l255_14;
  reg                 channels_3_interrupts_completion_enable;
  reg                 channels_3_interrupts_completion_valid;
  wire                when_DmaSg_l255_15;
  wire                when_DmaSg_l255_16;
  reg                 channels_3_interrupts_onChannelCompletion_enable;
  reg                 channels_3_interrupts_onChannelCompletion_valid;
  wire                when_DmaSg_l255_17;
  wire                io_inputs_0_fire;
  wire                when_package_l12;
  reg                 io_inputs_0_payload_last_regNextWhen;
  wire                when_package_l12_1;
  reg                 io_inputs_0_payload_last_regNextWhen_1;
  wire                when_package_l12_2;
  reg                 io_inputs_0_payload_last_regNextWhen_2;
  wire                when_package_l12_3;
  reg                 io_inputs_0_payload_last_regNextWhen_3;
  wire                when_package_l12_4;
  reg                 io_inputs_0_payload_last_regNextWhen_4;
  wire                when_package_l12_5;
  reg                 io_inputs_0_payload_last_regNextWhen_5;
  wire                when_package_l12_6;
  reg                 io_inputs_0_payload_last_regNextWhen_6;
  wire                when_package_l12_7;
  reg                 io_inputs_0_payload_last_regNextWhen_7;
  wire                when_package_l12_8;
  reg                 io_inputs_0_payload_last_regNextWhen_8;
  wire                when_package_l12_9;
  reg                 io_inputs_0_payload_last_regNextWhen_9;
  wire                when_package_l12_10;
  reg                 io_inputs_0_payload_last_regNextWhen_10;
  wire                when_package_l12_11;
  reg                 io_inputs_0_payload_last_regNextWhen_11;
  wire                when_package_l12_12;
  reg                 io_inputs_0_payload_last_regNextWhen_12;
  wire                when_package_l12_13;
  reg                 io_inputs_0_payload_last_regNextWhen_13;
  wire                when_package_l12_14;
  reg                 io_inputs_0_payload_last_regNextWhen_14;
  wire                when_package_l12_15;
  reg                 io_inputs_0_payload_last_regNextWhen_15;
  wire       [15:0]   s2b_0_cmd_firsts;
  wire                s2b_0_cmd_first;
  wire       [0:0]    s2b_0_cmd_channelsOh;
  wire                s2b_0_cmd_noHit;
  wire       [0:0]    s2b_0_cmd_channelsFull;
  reg                 io_inputs_0_thrown_valid;
  wire                io_inputs_0_thrown_ready;
  wire       [127:0]  io_inputs_0_thrown_payload_data;
  wire       [15:0]   io_inputs_0_thrown_payload_mask;
  wire       [3:0]    io_inputs_0_thrown_payload_sink;
  wire                io_inputs_0_thrown_payload_last;
  wire                _zz_io_inputs_0_thrown_ready;
  wire                s2b_0_cmd_sinkHalted_valid;
  wire                s2b_0_cmd_sinkHalted_ready;
  wire       [127:0]  s2b_0_cmd_sinkHalted_payload_data;
  wire       [15:0]   s2b_0_cmd_sinkHalted_payload_mask;
  wire       [3:0]    s2b_0_cmd_sinkHalted_payload_sink;
  wire                s2b_0_cmd_sinkHalted_payload_last;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_1;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_2;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_3;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_4;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_5;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_6;
  wire       [4:0]    _zz_s2b_0_cmd_byteCount_7;
  wire       [4:0]    s2b_0_cmd_byteCount;
  wire       [0:0]    s2b_0_cmd_context_channel;
  wire       [4:0]    s2b_0_cmd_context_bytes;
  wire                s2b_0_cmd_context_flush;
  wire                s2b_0_cmd_context_packet;
  wire                memory_core_io_writes_0_cmd_fire;
  wire                when_DmaSg_l665;
  wire       [0:0]    s2b_0_rsp_context_channel;
  wire       [4:0]    s2b_0_rsp_context_bytes;
  wire                s2b_0_rsp_context_flush;
  wire                s2b_0_rsp_context_packet;
  wire       [7:0]    _zz_s2b_0_rsp_context_channel;
  wire                _zz_channels_0_fifo_pop_bytesIncr_value;
  wire                when_DmaSg_l679;
  wire                when_DmaSg_l681;
  wire                when_DmaSg_l682;
  wire                io_inputs_1_fire;
  wire                when_package_l12_16;
  reg                 io_inputs_1_payload_last_regNextWhen;
  wire                when_package_l12_17;
  reg                 io_inputs_1_payload_last_regNextWhen_1;
  wire                when_package_l12_18;
  reg                 io_inputs_1_payload_last_regNextWhen_2;
  wire                when_package_l12_19;
  reg                 io_inputs_1_payload_last_regNextWhen_3;
  wire                when_package_l12_20;
  reg                 io_inputs_1_payload_last_regNextWhen_4;
  wire                when_package_l12_21;
  reg                 io_inputs_1_payload_last_regNextWhen_5;
  wire                when_package_l12_22;
  reg                 io_inputs_1_payload_last_regNextWhen_6;
  wire                when_package_l12_23;
  reg                 io_inputs_1_payload_last_regNextWhen_7;
  wire                when_package_l12_24;
  reg                 io_inputs_1_payload_last_regNextWhen_8;
  wire                when_package_l12_25;
  reg                 io_inputs_1_payload_last_regNextWhen_9;
  wire                when_package_l12_26;
  reg                 io_inputs_1_payload_last_regNextWhen_10;
  wire                when_package_l12_27;
  reg                 io_inputs_1_payload_last_regNextWhen_11;
  wire                when_package_l12_28;
  reg                 io_inputs_1_payload_last_regNextWhen_12;
  wire                when_package_l12_29;
  reg                 io_inputs_1_payload_last_regNextWhen_13;
  wire                when_package_l12_30;
  reg                 io_inputs_1_payload_last_regNextWhen_14;
  wire                when_package_l12_31;
  reg                 io_inputs_1_payload_last_regNextWhen_15;
  wire       [15:0]   s2b_1_cmd_firsts;
  wire                s2b_1_cmd_first;
  wire       [0:0]    s2b_1_cmd_channelsOh;
  wire                s2b_1_cmd_noHit;
  wire       [0:0]    s2b_1_cmd_channelsFull;
  reg                 io_inputs_1_thrown_valid;
  wire                io_inputs_1_thrown_ready;
  wire       [127:0]  io_inputs_1_thrown_payload_data;
  wire       [15:0]   io_inputs_1_thrown_payload_mask;
  wire       [3:0]    io_inputs_1_thrown_payload_sink;
  wire                io_inputs_1_thrown_payload_last;
  wire                _zz_io_inputs_1_thrown_ready;
  wire                s2b_1_cmd_sinkHalted_valid;
  wire                s2b_1_cmd_sinkHalted_ready;
  wire       [127:0]  s2b_1_cmd_sinkHalted_payload_data;
  wire       [15:0]   s2b_1_cmd_sinkHalted_payload_mask;
  wire       [3:0]    s2b_1_cmd_sinkHalted_payload_sink;
  wire                s2b_1_cmd_sinkHalted_payload_last;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_1;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_2;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_3;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_4;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_5;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_6;
  wire       [4:0]    _zz_s2b_1_cmd_byteCount_7;
  wire       [4:0]    s2b_1_cmd_byteCount;
  wire       [0:0]    s2b_1_cmd_context_channel;
  wire       [4:0]    s2b_1_cmd_context_bytes;
  wire                s2b_1_cmd_context_flush;
  wire                s2b_1_cmd_context_packet;
  wire                memory_core_io_writes_1_cmd_fire;
  wire                when_DmaSg_l665_1;
  wire       [0:0]    s2b_1_rsp_context_channel;
  wire       [4:0]    s2b_1_rsp_context_bytes;
  wire                s2b_1_rsp_context_flush;
  wire                s2b_1_rsp_context_packet;
  wire       [7:0]    _zz_s2b_1_rsp_context_channel;
  wire                _zz_channels_2_fifo_pop_bytesIncr_value;
  wire                when_DmaSg_l679_1;
  wire                when_DmaSg_l681_1;
  wire                when_DmaSg_l682_1;
  wire       [0:0]    b2s_0_cmd_channelsOh;
  wire       [0:0]    b2s_0_cmd_context_channel;
  wire                b2s_0_cmd_context_veryLast;
  wire                b2s_0_cmd_context_endPacket;
  wire       [13:0]   b2s_0_cmd_veryLastPtr;
  wire       [13:0]   b2s_0_cmd_address;
  wire       [0:0]    b2s_0_rsp_context_channel;
  wire                b2s_0_rsp_context_veryLast;
  wire                b2s_0_rsp_context_endPacket;
  wire       [2:0]    _zz_b2s_0_rsp_context_channel;
  wire                io_outputs_0_fire;
  wire                when_DmaSg_l725;
  wire                when_DmaSg_l726;
  wire       [0:0]    b2s_1_cmd_channelsOh;
  wire       [0:0]    b2s_1_cmd_context_channel;
  wire                b2s_1_cmd_context_veryLast;
  wire                b2s_1_cmd_context_endPacket;
  wire       [13:0]   b2s_1_cmd_veryLastPtr;
  wire       [13:0]   b2s_1_cmd_address;
  wire       [0:0]    b2s_1_rsp_context_channel;
  wire                b2s_1_rsp_context_veryLast;
  wire                b2s_1_rsp_context_endPacket;
  wire       [2:0]    _zz_b2s_1_rsp_context_channel;
  wire                io_outputs_1_fire;
  wire                when_DmaSg_l725_1;
  wire                when_DmaSg_l726_1;
  reg                 m2b_cmd_s0_valid;
  reg        [0:0]    m2b_cmd_s0_chosen;
  wire       [1:0]    _zz_m2b_cmd_s0_priority_masked;
  wire       [1:0]    _zz_m2b_cmd_s0_priority_masked_1;
  wire       [1:0]    _zz_m2b_cmd_s0_priority_masked_2;
  wire       [1:0]    m2b_cmd_s0_priority_masked;
  reg        [1:0]    m2b_cmd_s0_priority_roundRobins_0;
  reg        [1:0]    m2b_cmd_s0_priority_roundRobins_1;
  reg        [1:0]    m2b_cmd_s0_priority_roundRobins_2;
  reg        [1:0]    m2b_cmd_s0_priority_roundRobins_3;
  reg        [1:0]    m2b_cmd_s0_priority_counter;
  wire       [1:0]    _zz_m2b_cmd_s0_priority_chosenOh;
  wire       [3:0]    _zz_m2b_cmd_s0_priority_chosenOh_1;
  wire       [3:0]    _zz_m2b_cmd_s0_priority_chosenOh_2;
  wire       [1:0]    m2b_cmd_s0_priority_chosenOh;
  wire                _zz_m2b_cmd_s0_priority_chosen;
  wire       [0:0]    m2b_cmd_s0_priority_chosen;
  wire                m2b_cmd_s0_priority_weightLast;
  wire       [1:0]    m2b_cmd_s0_priority_contextNext;
  wire                when_DmaSg_l758;
  wire                when_DmaSg_l760;
  wire                when_DmaSg_l763;
  wire                when_DmaSg_l763_1;
  wire                when_DmaSg_l763_2;
  wire                when_DmaSg_l763_3;
  wire                when_DmaSg_l773;
  wire                when_DmaSg_l773_1;
  wire       [31:0]   m2b_cmd_s0_address;
  wire       [25:0]   m2b_cmd_s0_bytesLeft;
  wire       [12:0]   m2b_cmd_s0_readAddressBurstRange;
  wire       [12:0]   m2b_cmd_s0_lengthHead;
  wire       [12:0]   m2b_cmd_s0_length;
  wire                m2b_cmd_s0_lastBurst;
  reg                 m2b_cmd_s1_valid;
  reg        [31:0]   m2b_cmd_s1_address;
  reg        [12:0]   m2b_cmd_s1_length;
  reg                 m2b_cmd_s1_lastBurst;
  reg        [25:0]   m2b_cmd_s1_bytesLeft;
  wire       [0:0]    m2b_cmd_s1_context_channel;
  wire       [4:0]    m2b_cmd_s1_context_start;
  wire       [4:0]    m2b_cmd_s1_context_stop;
  wire       [12:0]   m2b_cmd_s1_context_length;
  wire                m2b_cmd_s1_context_last;
  wire       [31:0]   m2b_cmd_s1_addressNext;
  wire       [25:0]   m2b_cmd_s1_byteLeftNext;
  wire       [9:0]    m2b_cmd_s1_fifoPushDecr;
  wire                when_DmaSg_l828;
  wire                when_DmaSg_l828_1;
  wire       [0:0]    m2b_rsp_context_channel;
  wire       [4:0]    m2b_rsp_context_start;
  wire       [4:0]    m2b_rsp_context_stop;
  wire       [12:0]   m2b_rsp_context_length;
  wire                m2b_rsp_context_last;
  wire       [24:0]   _zz_m2b_rsp_context_channel;
  wire                m2b_rsp_veryLast;
  wire                io_read_rsp_fire;
  wire                when_DmaSg_l847;
  wire                when_DmaSg_l848;
  wire                when_DmaSg_l848_1;
  reg                 m2b_rsp_first;
  wire                m2b_rsp_writeContext_last;
  wire                m2b_rsp_writeContext_lastOfBurst;
  wire       [0:0]    m2b_rsp_writeContext_channel;
  wire       [5:0]    m2b_rsp_writeContext_loadByteInNextBeat;
  wire                memory_core_io_writes_2_cmd_fire;
  wire                m2b_writeRsp_context_last;
  wire                m2b_writeRsp_context_lastOfBurst;
  wire       [0:0]    m2b_writeRsp_context_channel;
  wire       [5:0]    m2b_writeRsp_context_loadByteInNextBeat;
  wire       [8:0]    _zz_m2b_writeRsp_context_last;
  wire                _zz_channels_1_fifo_pop_bytesIncr_value;
  wire                when_DmaSg_l893;
  wire                _zz_channels_3_fifo_pop_bytesIncr_value;
  wire                when_DmaSg_l893_1;
  reg                 b2m_fsm_sel_valid;
  reg                 b2m_fsm_sel_ready;
  reg        [0:0]    b2m_fsm_sel_channel;
  reg        [12:0]   b2m_fsm_sel_bytePerBurst;
  reg        [12:0]   b2m_fsm_sel_bytesInBurst;
  reg        [17:0]   b2m_fsm_sel_bytesInFifo;
  reg        [31:0]   b2m_fsm_sel_address;
  reg        [13:0]   b2m_fsm_sel_ptr;
  reg        [13:0]   b2m_fsm_sel_ptrMask;
  reg                 b2m_fsm_sel_flush;
  reg                 b2m_fsm_sel_packet;
  reg        [25:0]   b2m_fsm_sel_bytesLeft;
  reg                 b2m_fsm_arbiter_logic_valid;
  reg        [0:0]    b2m_fsm_arbiter_logic_chosen;
  wire       [1:0]    _zz_b2m_fsm_arbiter_logic_priority_masked;
  wire       [1:0]    _zz_b2m_fsm_arbiter_logic_priority_masked_1;
  wire       [1:0]    _zz_b2m_fsm_arbiter_logic_priority_masked_2;
  wire       [1:0]    b2m_fsm_arbiter_logic_priority_masked;
  reg        [1:0]    b2m_fsm_arbiter_logic_priority_roundRobins_0;
  reg        [1:0]    b2m_fsm_arbiter_logic_priority_roundRobins_1;
  reg        [1:0]    b2m_fsm_arbiter_logic_priority_roundRobins_2;
  reg        [1:0]    b2m_fsm_arbiter_logic_priority_roundRobins_3;
  reg        [1:0]    b2m_fsm_arbiter_logic_priority_counter;
  wire       [1:0]    _zz_b2m_fsm_arbiter_logic_priority_chosenOh;
  wire       [3:0]    _zz_b2m_fsm_arbiter_logic_priority_chosenOh_1;
  wire       [3:0]    _zz_b2m_fsm_arbiter_logic_priority_chosenOh_2;
  wire       [1:0]    b2m_fsm_arbiter_logic_priority_chosenOh;
  wire                _zz_b2m_fsm_arbiter_logic_priority_chosen;
  wire       [0:0]    b2m_fsm_arbiter_logic_priority_chosen;
  wire                b2m_fsm_arbiter_logic_priority_weightLast;
  wire       [1:0]    b2m_fsm_arbiter_logic_priority_contextNext;
  wire                when_DmaSg_l758_1;
  wire                when_DmaSg_l760_1;
  wire                when_DmaSg_l763_4;
  wire                when_DmaSg_l763_5;
  wire                when_DmaSg_l763_6;
  wire                when_DmaSg_l763_7;
  wire                when_DmaSg_l773_2;
  wire                when_DmaSg_l773_3;
  wire                when_DmaSg_l935;
  wire       [1:0]    _zz_1;
  wire       [13:0]   b2m_fsm_bytesInBurstP1;
  wire       [31:0]   b2m_fsm_addressNext;
  wire       [26:0]   b2m_fsm_bytesLeftNext;
  wire                b2m_fsm_isFinalCmd;
  reg        [7:0]    b2m_fsm_beatCounter;
  reg                 b2m_fsm_sel_valid_regNext;
  wire                b2m_fsm_s0;
  reg                 b2m_fsm_s1;
  reg                 b2m_fsm_s2;
  wire                when_DmaSg_l986;
  wire       [17:0]   _zz_b2m_fsm_sel_bytesInBurst;
  wire       [25:0]   _zz_b2m_fsm_sel_bytesInBurst_1;
  wire       [12:0]   _zz_b2m_fsm_sel_bytesInBurst_2;
  wire                b2m_fsm_fifoCompletion;
  wire                when_DmaSg_l996;
  wire                when_DmaSg_l1001;
  wire                when_DmaSg_l996_1;
  wire                when_DmaSg_l1001_1;
  reg                 b2m_fsm_toggle;
  wire                when_DmaSg_l1013;
  wire       [13:0]   b2m_fsm_fetch_context_ptr;
  wire                b2m_fsm_fetch_context_toggle;
  wire                when_DmaSg_l1033;
  wire       [13:0]   b2m_fsm_aggregate_context_ptr;
  wire                b2m_fsm_aggregate_context_toggle;
  wire       [14:0]   _zz_b2m_fsm_aggregate_context_ptr;
  wire                memory_core_io_reads_2_rsp_s2mPipe_valid;
  reg                 memory_core_io_reads_2_rsp_s2mPipe_ready;
  wire       [255:0]  memory_core_io_reads_2_rsp_s2mPipe_payload_data;
  wire       [31:0]   memory_core_io_reads_2_rsp_s2mPipe_payload_mask;
  wire       [14:0]   memory_core_io_reads_2_rsp_s2mPipe_payload_context;
  reg                 memory_core_io_reads_2_rsp_rValidN;
  reg        [255:0]  memory_core_io_reads_2_rsp_rData_data;
  reg        [31:0]   memory_core_io_reads_2_rsp_rData_mask;
  reg        [14:0]   memory_core_io_reads_2_rsp_rData_context;
  wire                when_Stream_l445;
  reg                 b2m_fsm_aggregate_memoryPort_valid;
  wire                b2m_fsm_aggregate_memoryPort_ready;
  wire       [255:0]  b2m_fsm_aggregate_memoryPort_payload_data;
  wire       [31:0]   b2m_fsm_aggregate_memoryPort_payload_mask;
  wire       [14:0]   b2m_fsm_aggregate_memoryPort_payload_context;
  reg                 b2m_fsm_aggregate_first;
  wire                b2m_fsm_aggregate_memoryPort_fire;
  wire                when_DmaSg_l1050;
  wire       [4:0]    b2m_fsm_aggregate_bytesToSkip;
  wire       [31:0]   b2m_fsm_aggregate_bytesToSkipMask;
  reg                 _zz_io_flush;
  wire       [4:0]    b2m_fsm_cmd_maskFirstTrigger;
  wire       [4:0]    b2m_fsm_cmd_maskLastTriggerComb;
  reg        [4:0]    b2m_fsm_cmd_maskLastTriggerReg;
  reg        [31:0]   b2m_fsm_cmd_maskLast;
  wire       [31:0]   b2m_fsm_cmd_maskFirst;
  wire                b2m_fsm_cmd_enoughAggregation;
  wire                io_write_cmd_fire;
  reg                 io_write_cmd_payload_first;
  wire                b2m_fsm_cmd_doPtrIncr;
  wire       [0:0]    b2m_fsm_cmd_context_channel;
  wire       [12:0]   b2m_fsm_cmd_context_length;
  wire                b2m_fsm_cmd_context_doPacketSync;
  wire                when_DmaSg_l1102;
  wire       [1:0]    _zz_2;
  wire       [4:0]    _zz_channels_0_pop_b2m_bytesToSkip;
  wire       [0:0]    b2m_rsp_context_channel;
  wire       [12:0]   b2m_rsp_context_length;
  wire                b2m_rsp_context_doPacketSync;
  wire       [14:0]   _zz_b2m_rsp_context_channel;
  wire                io_write_rsp_fire;
  wire       [1:0]    _zz_3;
  wire                when_DmaSg_l1116;
  wire                when_DmaSg_l1116_1;
  reg                 when_BusSlaveFactory_l377;
  wire                when_BusSlaveFactory_l379;
  reg                 when_BusSlaveFactory_l377_1;
  wire                when_BusSlaveFactory_l379_1;
  reg                 when_BusSlaveFactory_l341;
  wire                when_BusSlaveFactory_l347;
  reg                 when_BusSlaveFactory_l341_1;
  wire                when_BusSlaveFactory_l347_1;
  reg                 when_BusSlaveFactory_l341_2;
  wire                when_BusSlaveFactory_l347_2;
  reg                 when_BusSlaveFactory_l377_2;
  wire                when_BusSlaveFactory_l379_2;
  reg                 when_BusSlaveFactory_l377_3;
  wire                when_BusSlaveFactory_l379_3;
  reg                 when_BusSlaveFactory_l341_3;
  wire                when_BusSlaveFactory_l347_3;
  reg                 when_BusSlaveFactory_l341_4;
  wire                when_BusSlaveFactory_l347_4;
  reg                 when_BusSlaveFactory_l377_4;
  wire                when_BusSlaveFactory_l379_4;
  reg                 when_BusSlaveFactory_l377_5;
  wire                when_BusSlaveFactory_l379_5;
  reg                 when_BusSlaveFactory_l341_5;
  wire                when_BusSlaveFactory_l347_5;
  reg                 when_BusSlaveFactory_l341_6;
  wire                when_BusSlaveFactory_l347_6;
  reg                 when_BusSlaveFactory_l341_7;
  wire                when_BusSlaveFactory_l347_7;
  reg                 when_BusSlaveFactory_l377_6;
  wire                when_BusSlaveFactory_l379_6;
  reg                 when_BusSlaveFactory_l377_7;
  wire                when_BusSlaveFactory_l379_7;
  reg                 when_BusSlaveFactory_l341_8;
  wire                when_BusSlaveFactory_l347_8;
  reg                 when_BusSlaveFactory_l341_9;
  wire                when_BusSlaveFactory_l347_9;
  wire                when_Apb3SlaveFactory_l81;
  wire                when_Apb3SlaveFactory_l81_1;
  wire                when_Apb3SlaveFactory_l81_2;
  wire                when_Apb3SlaveFactory_l81_3;

  assign _zz_channels_0_fifo_pop_withOverride_backupNext = (channels_0_fifo_pop_withOverride_backup + channels_0_fifo_pop_bytesIncr_value);
  assign _zz_channels_0_fifo_pop_withOverride_exposed = (channels_0_fifo_pop_withOverride_exposed - channels_0_fifo_pop_bytesDecr_value);
  assign _zz_channels_0_pop_b2m_selfFlush = {9'd0, channels_0_fifo_pop_bytes};
  assign _zz_channels_0_pop_b2m_request = {5'd0, channels_0_pop_b2m_bytePerBurst};
  assign _zz_channels_0_pop_b2m_request_2 = (channels_0_fifo_words >>> 1'd1);
  assign _zz_channels_0_pop_b2m_request_1 = {1'd0, _zz_channels_0_pop_b2m_request_2};
  assign _zz_channels_0_pop_b2m_memPending = (channels_0_pop_b2m_memPending + _zz_channels_0_pop_b2m_memPending_1);
  assign _zz_channels_0_pop_b2m_memPending_2 = channels_0_pop_b2m_memPendingInc;
  assign _zz_channels_0_pop_b2m_memPending_1 = {3'd0, _zz_channels_0_pop_b2m_memPending_2};
  assign _zz_channels_0_pop_b2m_memPending_4 = channels_0_pop_b2m_memRsp;
  assign _zz_channels_0_pop_b2m_memPending_3 = {3'd0, _zz_channels_0_pop_b2m_memPending_4};
  assign _zz_channels_0_pop_b2m_address = (channels_0_pop_b2m_address - _zz_channels_0_pop_b2m_address_1);
  assign _zz_channels_0_pop_b2m_address_1 = {6'd0, channels_0_bytes};
  assign _zz_channels_0_fifo_push_available = (channels_0_fifo_push_available + channels_0_fifo_pop_ptrIncr_value_regNext);
  assign _zz_channels_1_fifo_pop_withoutOverride_exposed = (channels_1_fifo_pop_withoutOverride_exposed + channels_1_fifo_pop_bytesIncr_value);
  assign _zz_channels_1_push_m2b_memPending = (channels_1_push_m2b_memPending + _zz_channels_1_push_m2b_memPending_1);
  assign _zz_channels_1_push_m2b_memPending_2 = channels_1_push_m2b_memPendingIncr;
  assign _zz_channels_1_push_m2b_memPending_1 = {3'd0, _zz_channels_1_push_m2b_memPending_2};
  assign _zz_channels_1_push_m2b_memPending_4 = channels_1_push_m2b_memPendingDecr;
  assign _zz_channels_1_push_m2b_memPending_3 = {3'd0, _zz_channels_1_push_m2b_memPending_4};
  assign _zz_channels_1_push_m2b_loadRequest_1 = (channels_1_push_m2b_bytePerBurst >>> 3'd4);
  assign _zz_channels_1_push_m2b_loadRequest = {5'd0, _zz_channels_1_push_m2b_loadRequest_1};
  assign _zz_when_DmaSg_l486 = {13'd0, channels_1_push_m2b_bytePerBurst};
  assign _zz_channels_1_push_m2b_address = (channels_1_push_m2b_address - _zz_channels_1_push_m2b_address_1);
  assign _zz_channels_1_push_m2b_address_1 = {6'd0, channels_1_bytes};
  assign _zz_channels_1_fifo_push_available = (channels_1_fifo_push_available + channels_1_fifo_pop_ptrIncr_value_regNext);
  assign _zz_channels_2_fifo_pop_withOverride_backupNext = (channels_2_fifo_pop_withOverride_backup + channels_2_fifo_pop_bytesIncr_value);
  assign _zz_channels_2_fifo_pop_withOverride_exposed = (channels_2_fifo_pop_withOverride_exposed - channels_2_fifo_pop_bytesDecr_value);
  assign _zz_channels_2_pop_b2m_selfFlush = {9'd0, channels_2_fifo_pop_bytes};
  assign _zz_channels_2_pop_b2m_request = {5'd0, channels_2_pop_b2m_bytePerBurst};
  assign _zz_channels_2_pop_b2m_request_2 = (channels_2_fifo_words >>> 1'd1);
  assign _zz_channels_2_pop_b2m_request_1 = {1'd0, _zz_channels_2_pop_b2m_request_2};
  assign _zz_channels_2_pop_b2m_memPending = (channels_2_pop_b2m_memPending + _zz_channels_2_pop_b2m_memPending_1);
  assign _zz_channels_2_pop_b2m_memPending_2 = channels_2_pop_b2m_memPendingInc;
  assign _zz_channels_2_pop_b2m_memPending_1 = {3'd0, _zz_channels_2_pop_b2m_memPending_2};
  assign _zz_channels_2_pop_b2m_memPending_4 = channels_2_pop_b2m_memRsp;
  assign _zz_channels_2_pop_b2m_memPending_3 = {3'd0, _zz_channels_2_pop_b2m_memPending_4};
  assign _zz_channels_2_pop_b2m_address = (channels_2_pop_b2m_address - _zz_channels_2_pop_b2m_address_1);
  assign _zz_channels_2_pop_b2m_address_1 = {6'd0, channels_2_bytes};
  assign _zz_channels_2_fifo_push_available = (channels_2_fifo_push_available + channels_2_fifo_pop_ptrIncr_value_regNext);
  assign _zz_channels_3_fifo_pop_withoutOverride_exposed = (channels_3_fifo_pop_withoutOverride_exposed + channels_3_fifo_pop_bytesIncr_value);
  assign _zz_channels_3_push_m2b_memPending = (channels_3_push_m2b_memPending + _zz_channels_3_push_m2b_memPending_1);
  assign _zz_channels_3_push_m2b_memPending_2 = channels_3_push_m2b_memPendingIncr;
  assign _zz_channels_3_push_m2b_memPending_1 = {3'd0, _zz_channels_3_push_m2b_memPending_2};
  assign _zz_channels_3_push_m2b_memPending_4 = channels_3_push_m2b_memPendingDecr;
  assign _zz_channels_3_push_m2b_memPending_3 = {3'd0, _zz_channels_3_push_m2b_memPending_4};
  assign _zz_channels_3_push_m2b_loadRequest_1 = (channels_3_push_m2b_bytePerBurst >>> 3'd4);
  assign _zz_channels_3_push_m2b_loadRequest = {5'd0, _zz_channels_3_push_m2b_loadRequest_1};
  assign _zz_when_DmaSg_l486_1 = {13'd0, channels_3_push_m2b_bytePerBurst};
  assign _zz_channels_3_push_m2b_address = (channels_3_push_m2b_address - _zz_channels_3_push_m2b_address_1);
  assign _zz_channels_3_push_m2b_address_1 = {6'd0, channels_3_bytes};
  assign _zz_channels_3_fifo_push_available = (channels_3_fifo_push_available + channels_3_fifo_pop_ptrIncr_value_regNext);
  assign _zz_s2b_0_cmd_byteCount_8 = (_zz_s2b_0_cmd_byteCount_9 + _zz_s2b_0_cmd_byteCount_14);
  assign _zz_s2b_0_cmd_byteCount_9 = (_zz_s2b_0_cmd_byteCount_10 + _zz_s2b_0_cmd_byteCount_12);
  assign _zz_s2b_0_cmd_byteCount_14 = (_zz_s2b_0_cmd_byteCount_15 + _zz_s2b_0_cmd_byteCount_17);
  assign _zz_s2b_0_cmd_byteCount_19 = (_zz_s2b_0_cmd_byteCount_20 + _zz_s2b_0_cmd_byteCount_22);
  assign _zz_s2b_0_cmd_byteCount_24 = s2b_0_cmd_sinkHalted_payload_mask[15];
  assign _zz_s2b_0_cmd_byteCount_23 = {2'd0, _zz_s2b_0_cmd_byteCount_24};
  assign _zz_s2b_1_cmd_byteCount_8 = (_zz_s2b_1_cmd_byteCount_9 + _zz_s2b_1_cmd_byteCount_14);
  assign _zz_s2b_1_cmd_byteCount_9 = (_zz_s2b_1_cmd_byteCount_10 + _zz_s2b_1_cmd_byteCount_12);
  assign _zz_s2b_1_cmd_byteCount_14 = (_zz_s2b_1_cmd_byteCount_15 + _zz_s2b_1_cmd_byteCount_17);
  assign _zz_s2b_1_cmd_byteCount_19 = (_zz_s2b_1_cmd_byteCount_20 + _zz_s2b_1_cmd_byteCount_22);
  assign _zz_s2b_1_cmd_byteCount_24 = s2b_1_cmd_sinkHalted_payload_mask[15];
  assign _zz_s2b_1_cmd_byteCount_23 = {2'd0, _zz_s2b_1_cmd_byteCount_24};
  assign _zz__zz_m2b_cmd_s0_priority_chosenOh_2 = (_zz_m2b_cmd_s0_priority_chosenOh_1 - _zz__zz_m2b_cmd_s0_priority_chosenOh_2_1);
  assign _zz__zz_m2b_cmd_s0_priority_chosenOh_2_2 = _zz__zz_m2b_cmd_s0_priority_chosenOh_2_3;
  assign _zz__zz_m2b_cmd_s0_priority_chosenOh_2_1 = {2'd0, _zz__zz_m2b_cmd_s0_priority_chosenOh_2_2};
  assign _zz_m2b_cmd_s0_length = ((_zz_m2b_cmd_s0_length_1 < m2b_cmd_s0_bytesLeft) ? _zz_m2b_cmd_s0_length_2 : m2b_cmd_s0_bytesLeft);
  assign _zz_m2b_cmd_s0_length_1 = {13'd0, m2b_cmd_s0_lengthHead};
  assign _zz_m2b_cmd_s0_length_2 = {13'd0, m2b_cmd_s0_lengthHead};
  assign _zz_m2b_cmd_s0_lastBurst = {13'd0, m2b_cmd_s0_length};
  assign _zz_m2b_cmd_s1_context_stop = (m2b_cmd_s1_address + _zz_m2b_cmd_s1_context_stop_1);
  assign _zz_m2b_cmd_s1_context_stop_1 = {19'd0, m2b_cmd_s1_length};
  assign _zz_m2b_cmd_s1_addressNext = (m2b_cmd_s1_address + _zz_m2b_cmd_s1_addressNext_1);
  assign _zz_m2b_cmd_s1_addressNext_1 = {19'd0, m2b_cmd_s1_length};
  assign _zz_m2b_cmd_s1_byteLeftNext = (m2b_cmd_s1_bytesLeft - _zz_m2b_cmd_s1_byteLeftNext_1);
  assign _zz_m2b_cmd_s1_byteLeftNext_1 = {13'd0, m2b_cmd_s1_length};
  assign _zz_m2b_cmd_s1_fifoPushDecr = ({1'b0,(_zz_m2b_cmd_s1_fifoPushDecr_1 | 13'h001f)} + _zz_m2b_cmd_s1_fifoPushDecr_4);
  assign _zz_m2b_cmd_s1_fifoPushDecr_1 = (_zz_m2b_cmd_s1_fifoPushDecr_2 + io_read_cmd_payload_fragment_length);
  assign _zz_m2b_cmd_s1_fifoPushDecr_3 = m2b_cmd_s1_address[4 : 0];
  assign _zz_m2b_cmd_s1_fifoPushDecr_2 = {8'd0, _zz_m2b_cmd_s1_fifoPushDecr_3};
  assign _zz_m2b_cmd_s1_fifoPushDecr_5 = {1'b0,1'b1};
  assign _zz_m2b_cmd_s1_fifoPushDecr_4 = {12'd0, _zz_m2b_cmd_s1_fifoPushDecr_5};
  assign _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2 = (_zz_b2m_fsm_arbiter_logic_priority_chosenOh_1 - _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_1);
  assign _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_2 = _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_3;
  assign _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_1 = {2'd0, _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_2};
  assign _zz_b2m_fsm_bytesInBurstP1_1 = {1'b0,1'b1};
  assign _zz_b2m_fsm_bytesInBurstP1 = {12'd0, _zz_b2m_fsm_bytesInBurstP1_1};
  assign _zz_b2m_fsm_addressNext = {18'd0, b2m_fsm_bytesInBurstP1};
  assign _zz_b2m_fsm_bytesLeftNext_1 = {1'b0,b2m_fsm_bytesInBurstP1};
  assign _zz_b2m_fsm_bytesLeftNext = {12'd0, _zz_b2m_fsm_bytesLeftNext_1};
  assign _zz__zz_b2m_fsm_sel_bytesInBurst_1 = {8'd0, _zz_b2m_fsm_sel_bytesInBurst};
  assign _zz__zz_b2m_fsm_sel_bytesInBurst_1_1 = {8'd0, _zz_b2m_fsm_sel_bytesInBurst};
  assign _zz__zz_b2m_fsm_sel_bytesInBurst_2 = b2m_fsm_sel_address[12:0];
  assign _zz_b2m_fsm_sel_bytesInBurst_3 = ((_zz_b2m_fsm_sel_bytesInBurst_1 < _zz_b2m_fsm_sel_bytesInBurst_4) ? _zz_b2m_fsm_sel_bytesInBurst_1 : _zz_b2m_fsm_sel_bytesInBurst_5);
  assign _zz_b2m_fsm_sel_bytesInBurst_4 = {13'd0, _zz_b2m_fsm_sel_bytesInBurst_2};
  assign _zz_b2m_fsm_sel_bytesInBurst_5 = {13'd0, _zz_b2m_fsm_sel_bytesInBurst_2};
  assign _zz_b2m_fsm_fifoCompletion = {5'd0, b2m_fsm_sel_bytesInBurst};
  assign _zz_b2m_fsm_fifoCompletion_1 = (b2m_fsm_sel_bytesInFifo - 18'h00001);
  assign _zz_b2m_fsm_beatCounter = (_zz_b2m_fsm_beatCounter_1 + b2m_fsm_sel_bytesInBurst);
  assign _zz_b2m_fsm_beatCounter_2 = b2m_fsm_sel_address[4 : 0];
  assign _zz_b2m_fsm_beatCounter_1 = {8'd0, _zz_b2m_fsm_beatCounter_2};
  assign _zz_b2m_fsm_sel_ptr_1 = (b2m_fsm_sel_ptr + 14'h0002);
  assign _zz_b2m_fsm_cmd_maskLastTriggerComb = b2m_fsm_sel_bytesInBurst[4:0];
  assign _zz_channels_0_channelStart = 1'b1;
  assign _zz_channels_0_ctrl_kick = 1'b1;
  assign _zz_channels_0_interrupts_completion_valid = 1'b0;
  assign _zz_channels_0_interrupts_onChannelCompletion_valid = 1'b0;
  assign _zz_channels_0_interrupts_s2mPacket_valid = 1'b0;
  assign _zz_channels_1_channelStart = 1'b1;
  assign _zz_channels_1_ctrl_kick = 1'b1;
  assign _zz_channels_1_interrupts_completion_valid = 1'b0;
  assign _zz_channels_1_interrupts_onChannelCompletion_valid = 1'b0;
  assign _zz_channels_2_channelStart = 1'b1;
  assign _zz_channels_2_ctrl_kick = 1'b1;
  assign _zz_channels_2_interrupts_completion_valid = 1'b0;
  assign _zz_channels_2_interrupts_onChannelCompletion_valid = 1'b0;
  assign _zz_channels_2_interrupts_s2mPacket_valid = 1'b0;
  assign _zz_channels_3_channelStart = 1'b1;
  assign _zz_channels_3_ctrl_kick = 1'b1;
  assign _zz_channels_3_interrupts_completion_valid = 1'b0;
  assign _zz_channels_3_interrupts_onChannelCompletion_valid = 1'b0;
  assign _zz_channels_0_fifo_push_ptrIncr_value_1 = ((when_DmaSg_l665 && (|s2b_0_cmd_sinkHalted_payload_mask)) ? 1'b1 : 1'b0);
  assign _zz_channels_0_fifo_push_ptrIncr_value = {13'd0, _zz_channels_0_fifo_push_ptrIncr_value_1};
  assign _zz_channels_0_fifo_pop_bytesIncr_value_2 = (_zz_channels_0_fifo_pop_bytesIncr_value ? s2b_0_rsp_context_bytes : 5'h0);
  assign _zz_channels_0_fifo_pop_bytesIncr_value_1 = {13'd0, _zz_channels_0_fifo_pop_bytesIncr_value_2};
  assign _zz_channels_0_fifo_pop_ptrIncr_value_1 = ((b2m_fsm_cmd_doPtrIncr && (b2m_fsm_sel_channel == 1'b0)) ? 2'b10 : 2'b00);
  assign _zz_channels_0_fifo_pop_ptrIncr_value = {12'd0, _zz_channels_0_fifo_pop_ptrIncr_value_1};
  assign _zz_channels_1_fifo_push_ptrIncr_value_1 = ((memory_core_io_writes_2_cmd_fire && (m2b_rsp_context_channel == 1'b0)) ? 2'b10 : 2'b00);
  assign _zz_channels_1_fifo_push_ptrIncr_value = {12'd0, _zz_channels_1_fifo_push_ptrIncr_value_1};
  assign _zz_channels_1_fifo_pop_bytesIncr_value_2 = (_zz_channels_1_fifo_pop_bytesIncr_value ? _zz_channels_1_fifo_pop_bytesIncr_value_3 : 6'h0);
  assign _zz_channels_1_fifo_pop_bytesIncr_value_1 = {12'd0, _zz_channels_1_fifo_pop_bytesIncr_value_2};
  assign _zz_channels_1_fifo_pop_bytesIncr_value_3 = (m2b_writeRsp_context_loadByteInNextBeat + 6'h01);
  assign _zz_channels_1_fifo_pop_ptrIncr_value_1 = ((b2s_0_cmd_channelsOh[0] && memory_core_io_reads_0_cmd_ready) ? 1'b1 : 1'b0);
  assign _zz_channels_1_fifo_pop_ptrIncr_value = {13'd0, _zz_channels_1_fifo_pop_ptrIncr_value_1};
  assign _zz_channels_2_fifo_push_ptrIncr_value_1 = ((when_DmaSg_l665_1 && (|s2b_1_cmd_sinkHalted_payload_mask)) ? 1'b1 : 1'b0);
  assign _zz_channels_2_fifo_push_ptrIncr_value = {13'd0, _zz_channels_2_fifo_push_ptrIncr_value_1};
  assign _zz_channels_2_fifo_pop_bytesIncr_value_2 = (_zz_channels_2_fifo_pop_bytesIncr_value ? s2b_1_rsp_context_bytes : 5'h0);
  assign _zz_channels_2_fifo_pop_bytesIncr_value_1 = {13'd0, _zz_channels_2_fifo_pop_bytesIncr_value_2};
  assign _zz_channels_2_fifo_pop_ptrIncr_value_1 = ((b2m_fsm_cmd_doPtrIncr && (b2m_fsm_sel_channel == 1'b1)) ? 2'b10 : 2'b00);
  assign _zz_channels_2_fifo_pop_ptrIncr_value = {12'd0, _zz_channels_2_fifo_pop_ptrIncr_value_1};
  assign _zz_channels_3_fifo_push_ptrIncr_value_1 = ((memory_core_io_writes_2_cmd_fire && (m2b_rsp_context_channel == 1'b1)) ? 2'b10 : 2'b00);
  assign _zz_channels_3_fifo_push_ptrIncr_value = {12'd0, _zz_channels_3_fifo_push_ptrIncr_value_1};
  assign _zz_channels_3_fifo_pop_bytesIncr_value_2 = (_zz_channels_3_fifo_pop_bytesIncr_value ? _zz_channels_3_fifo_pop_bytesIncr_value_3 : 6'h0);
  assign _zz_channels_3_fifo_pop_bytesIncr_value_1 = {12'd0, _zz_channels_3_fifo_pop_bytesIncr_value_2};
  assign _zz_channels_3_fifo_pop_bytesIncr_value_3 = (m2b_writeRsp_context_loadByteInNextBeat + 6'h01);
  assign _zz_channels_3_fifo_pop_ptrIncr_value_1 = ((b2s_1_cmd_channelsOh[0] && memory_core_io_reads_1_cmd_ready) ? 1'b1 : 1'b0);
  assign _zz_channels_3_fifo_pop_ptrIncr_value = {13'd0, _zz_channels_3_fifo_pop_ptrIncr_value_1};
  assign _zz_s2b_0_cmd_byteCount_11 = {s2b_0_cmd_sinkHalted_payload_mask[2],{s2b_0_cmd_sinkHalted_payload_mask[1],s2b_0_cmd_sinkHalted_payload_mask[0]}};
  assign _zz_s2b_0_cmd_byteCount_13 = {s2b_0_cmd_sinkHalted_payload_mask[5],{s2b_0_cmd_sinkHalted_payload_mask[4],s2b_0_cmd_sinkHalted_payload_mask[3]}};
  assign _zz_s2b_0_cmd_byteCount_16 = {s2b_0_cmd_sinkHalted_payload_mask[8],{s2b_0_cmd_sinkHalted_payload_mask[7],s2b_0_cmd_sinkHalted_payload_mask[6]}};
  assign _zz_s2b_0_cmd_byteCount_18 = {s2b_0_cmd_sinkHalted_payload_mask[11],{s2b_0_cmd_sinkHalted_payload_mask[10],s2b_0_cmd_sinkHalted_payload_mask[9]}};
  assign _zz_s2b_0_cmd_byteCount_21 = {s2b_0_cmd_sinkHalted_payload_mask[14],{s2b_0_cmd_sinkHalted_payload_mask[13],s2b_0_cmd_sinkHalted_payload_mask[12]}};
  assign _zz_s2b_1_cmd_byteCount_11 = {s2b_1_cmd_sinkHalted_payload_mask[2],{s2b_1_cmd_sinkHalted_payload_mask[1],s2b_1_cmd_sinkHalted_payload_mask[0]}};
  assign _zz_s2b_1_cmd_byteCount_13 = {s2b_1_cmd_sinkHalted_payload_mask[5],{s2b_1_cmd_sinkHalted_payload_mask[4],s2b_1_cmd_sinkHalted_payload_mask[3]}};
  assign _zz_s2b_1_cmd_byteCount_16 = {s2b_1_cmd_sinkHalted_payload_mask[8],{s2b_1_cmd_sinkHalted_payload_mask[7],s2b_1_cmd_sinkHalted_payload_mask[6]}};
  assign _zz_s2b_1_cmd_byteCount_18 = {s2b_1_cmd_sinkHalted_payload_mask[11],{s2b_1_cmd_sinkHalted_payload_mask[10],s2b_1_cmd_sinkHalted_payload_mask[9]}};
  assign _zz_s2b_1_cmd_byteCount_21 = {s2b_1_cmd_sinkHalted_payload_mask[14],{s2b_1_cmd_sinkHalted_payload_mask[13],s2b_1_cmd_sinkHalted_payload_mask[12]}};
  assign _zz_s2b_0_cmd_firsts = io_inputs_0_payload_last_regNextWhen_5;
  assign _zz_s2b_0_cmd_firsts_1 = {io_inputs_0_payload_last_regNextWhen_4,{io_inputs_0_payload_last_regNextWhen_3,{io_inputs_0_payload_last_regNextWhen_2,{io_inputs_0_payload_last_regNextWhen_1,io_inputs_0_payload_last_regNextWhen}}}};
  assign _zz_s2b_1_cmd_firsts = io_inputs_1_payload_last_regNextWhen_5;
  assign _zz_s2b_1_cmd_firsts_1 = {io_inputs_1_payload_last_regNextWhen_4,{io_inputs_1_payload_last_regNextWhen_3,{io_inputs_1_payload_last_regNextWhen_2,{io_inputs_1_payload_last_regNextWhen_1,io_inputs_1_payload_last_regNextWhen}}}};
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask = 5'h1d;
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_1 = (! b2m_fsm_aggregate_first);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_2 = (b2m_fsm_aggregate_bytesToSkip <= 5'h1c);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_3 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h1b));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_4 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h1a));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_5 = {((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h19)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h18)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= _zz_b2m_fsm_aggregate_bytesToSkipMask_6)),{(_zz_b2m_fsm_aggregate_bytesToSkipMask_7 || _zz_b2m_fsm_aggregate_bytesToSkipMask_8),{_zz_b2m_fsm_aggregate_bytesToSkipMask_9,{_zz_b2m_fsm_aggregate_bytesToSkipMask_10,_zz_b2m_fsm_aggregate_bytesToSkipMask_11}}}}}};
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_6 = 5'h17;
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_7 = (! b2m_fsm_aggregate_first);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_8 = (b2m_fsm_aggregate_bytesToSkip <= 5'h16);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_9 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h15));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_10 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h14));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_11 = {((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h13)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h12)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= _zz_b2m_fsm_aggregate_bytesToSkipMask_12)),{(_zz_b2m_fsm_aggregate_bytesToSkipMask_13 || _zz_b2m_fsm_aggregate_bytesToSkipMask_14),{_zz_b2m_fsm_aggregate_bytesToSkipMask_15,{_zz_b2m_fsm_aggregate_bytesToSkipMask_16,_zz_b2m_fsm_aggregate_bytesToSkipMask_17}}}}}};
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_12 = 5'h11;
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_13 = (! b2m_fsm_aggregate_first);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_14 = (b2m_fsm_aggregate_bytesToSkip <= 5'h10);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_15 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h0f));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_16 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h0e));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_17 = {((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h0d)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h0c)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= _zz_b2m_fsm_aggregate_bytesToSkipMask_18)),{(_zz_b2m_fsm_aggregate_bytesToSkipMask_19 || _zz_b2m_fsm_aggregate_bytesToSkipMask_20),{_zz_b2m_fsm_aggregate_bytesToSkipMask_21,{_zz_b2m_fsm_aggregate_bytesToSkipMask_22,_zz_b2m_fsm_aggregate_bytesToSkipMask_23}}}}}};
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_18 = 5'h0b;
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_19 = (! b2m_fsm_aggregate_first);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_20 = (b2m_fsm_aggregate_bytesToSkip <= 5'h0a);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_21 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h09));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_22 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h08));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_23 = {((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h07)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h06)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= _zz_b2m_fsm_aggregate_bytesToSkipMask_24)),{(_zz_b2m_fsm_aggregate_bytesToSkipMask_25 || _zz_b2m_fsm_aggregate_bytesToSkipMask_26),{_zz_b2m_fsm_aggregate_bytesToSkipMask_27,{_zz_b2m_fsm_aggregate_bytesToSkipMask_28,_zz_b2m_fsm_aggregate_bytesToSkipMask_29}}}}}};
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_24 = 5'h05;
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_25 = (! b2m_fsm_aggregate_first);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_26 = (b2m_fsm_aggregate_bytesToSkip <= 5'h04);
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_27 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h03));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_28 = ((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h02));
  assign _zz_b2m_fsm_aggregate_bytesToSkipMask_29 = {((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h01)),((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h0))};
  assign _zz_b2m_fsm_cmd_maskLast = 5'h1a;
  assign _zz_b2m_fsm_cmd_maskLast_1 = (5'h19 <= b2m_fsm_cmd_maskLastTriggerComb);
  assign _zz_b2m_fsm_cmd_maskLast_2 = (5'h18 <= b2m_fsm_cmd_maskLastTriggerComb);
  assign _zz_b2m_fsm_cmd_maskLast_3 = {(5'h17 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h16 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h15 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h14 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h13 <= b2m_fsm_cmd_maskLastTriggerComb),{(_zz_b2m_fsm_cmd_maskLast_4 <= b2m_fsm_cmd_maskLastTriggerComb),{_zz_b2m_fsm_cmd_maskLast_5,{_zz_b2m_fsm_cmd_maskLast_6,_zz_b2m_fsm_cmd_maskLast_7}}}}}}}};
  assign _zz_b2m_fsm_cmd_maskLast_4 = 5'h12;
  assign _zz_b2m_fsm_cmd_maskLast_5 = (5'h11 <= b2m_fsm_cmd_maskLastTriggerComb);
  assign _zz_b2m_fsm_cmd_maskLast_6 = (5'h10 <= b2m_fsm_cmd_maskLastTriggerComb);
  assign _zz_b2m_fsm_cmd_maskLast_7 = {(5'h0f <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h0e <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h0d <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h0c <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h0b <= b2m_fsm_cmd_maskLastTriggerComb),{(_zz_b2m_fsm_cmd_maskLast_8 <= b2m_fsm_cmd_maskLastTriggerComb),{_zz_b2m_fsm_cmd_maskLast_9,{_zz_b2m_fsm_cmd_maskLast_10,_zz_b2m_fsm_cmd_maskLast_11}}}}}}}};
  assign _zz_b2m_fsm_cmd_maskLast_8 = 5'h0a;
  assign _zz_b2m_fsm_cmd_maskLast_9 = (5'h09 <= b2m_fsm_cmd_maskLastTriggerComb);
  assign _zz_b2m_fsm_cmd_maskLast_10 = (5'h08 <= b2m_fsm_cmd_maskLastTriggerComb);
  assign _zz_b2m_fsm_cmd_maskLast_11 = {(5'h07 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h06 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h05 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h04 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h03 <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h02 <= b2m_fsm_cmd_maskLastTriggerComb),{(_zz_b2m_fsm_cmd_maskLast_12 <= b2m_fsm_cmd_maskLastTriggerComb),(_zz_b2m_fsm_cmd_maskLast_13 <= b2m_fsm_cmd_maskLastTriggerComb)}}}}}}};
  assign _zz_b2m_fsm_cmd_maskLast_12 = 5'h01;
  assign _zz_b2m_fsm_cmd_maskLast_13 = 5'h0;
  assign _zz_b2m_fsm_cmd_maskFirst = 5'h1a;
  assign _zz_b2m_fsm_cmd_maskFirst_1 = (b2m_fsm_cmd_maskFirstTrigger <= 5'h19);
  assign _zz_b2m_fsm_cmd_maskFirst_2 = (b2m_fsm_cmd_maskFirstTrigger <= 5'h18);
  assign _zz_b2m_fsm_cmd_maskFirst_3 = {(b2m_fsm_cmd_maskFirstTrigger <= 5'h17),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h16),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h15),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h14),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h13),{(b2m_fsm_cmd_maskFirstTrigger <= _zz_b2m_fsm_cmd_maskFirst_4),{_zz_b2m_fsm_cmd_maskFirst_5,{_zz_b2m_fsm_cmd_maskFirst_6,_zz_b2m_fsm_cmd_maskFirst_7}}}}}}}};
  assign _zz_b2m_fsm_cmd_maskFirst_4 = 5'h12;
  assign _zz_b2m_fsm_cmd_maskFirst_5 = (b2m_fsm_cmd_maskFirstTrigger <= 5'h11);
  assign _zz_b2m_fsm_cmd_maskFirst_6 = (b2m_fsm_cmd_maskFirstTrigger <= 5'h10);
  assign _zz_b2m_fsm_cmd_maskFirst_7 = {(b2m_fsm_cmd_maskFirstTrigger <= 5'h0f),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h0e),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h0d),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h0c),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h0b),{(b2m_fsm_cmd_maskFirstTrigger <= _zz_b2m_fsm_cmd_maskFirst_8),{_zz_b2m_fsm_cmd_maskFirst_9,{_zz_b2m_fsm_cmd_maskFirst_10,_zz_b2m_fsm_cmd_maskFirst_11}}}}}}}};
  assign _zz_b2m_fsm_cmd_maskFirst_8 = 5'h0a;
  assign _zz_b2m_fsm_cmd_maskFirst_9 = (b2m_fsm_cmd_maskFirstTrigger <= 5'h09);
  assign _zz_b2m_fsm_cmd_maskFirst_10 = (b2m_fsm_cmd_maskFirstTrigger <= 5'h08);
  assign _zz_b2m_fsm_cmd_maskFirst_11 = {(b2m_fsm_cmd_maskFirstTrigger <= 5'h07),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h06),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h05),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h04),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h03),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h02),{(b2m_fsm_cmd_maskFirstTrigger <= _zz_b2m_fsm_cmd_maskFirst_12),(b2m_fsm_cmd_maskFirstTrigger <= _zz_b2m_fsm_cmd_maskFirst_13)}}}}}}};
  assign _zz_b2m_fsm_cmd_maskFirst_12 = 5'h01;
  assign _zz_b2m_fsm_cmd_maskFirst_13 = 5'h0;
  EfxDMA_DmaMemoryCore memory_core (
    .io_writes_0_cmd_valid            (s2b_0_cmd_sinkHalted_valid                       ), //i
    .io_writes_0_cmd_ready            (memory_core_io_writes_0_cmd_ready                ), //o
    .io_writes_0_cmd_payload_address  (memory_core_io_writes_0_cmd_payload_address[12:0]), //i
    .io_writes_0_cmd_payload_data     (s2b_0_cmd_sinkHalted_payload_data[127:0]         ), //i
    .io_writes_0_cmd_payload_mask     (s2b_0_cmd_sinkHalted_payload_mask[15:0]          ), //i
    .io_writes_0_cmd_payload_priority (channels_0_priority[1:0]                         ), //i
    .io_writes_0_cmd_payload_context  (memory_core_io_writes_0_cmd_payload_context[7:0] ), //i
    .io_writes_0_rsp_valid            (memory_core_io_writes_0_rsp_valid                ), //o
    .io_writes_0_rsp_payload_context  (memory_core_io_writes_0_rsp_payload_context[7:0] ), //o
    .io_writes_1_cmd_valid            (s2b_1_cmd_sinkHalted_valid                       ), //i
    .io_writes_1_cmd_ready            (memory_core_io_writes_1_cmd_ready                ), //o
    .io_writes_1_cmd_payload_address  (memory_core_io_writes_1_cmd_payload_address[12:0]), //i
    .io_writes_1_cmd_payload_data     (s2b_1_cmd_sinkHalted_payload_data[127:0]         ), //i
    .io_writes_1_cmd_payload_mask     (s2b_1_cmd_sinkHalted_payload_mask[15:0]          ), //i
    .io_writes_1_cmd_payload_priority (channels_2_priority[1:0]                         ), //i
    .io_writes_1_cmd_payload_context  (memory_core_io_writes_1_cmd_payload_context[7:0] ), //i
    .io_writes_1_rsp_valid            (memory_core_io_writes_1_rsp_valid                ), //o
    .io_writes_1_rsp_payload_context  (memory_core_io_writes_1_rsp_payload_context[7:0] ), //o
    .io_writes_2_cmd_valid            (io_read_rsp_valid                                ), //i
    .io_writes_2_cmd_ready            (memory_core_io_writes_2_cmd_ready                ), //o
    .io_writes_2_cmd_payload_address  (memory_core_io_writes_2_cmd_payload_address[12:0]), //i
    .io_writes_2_cmd_payload_data     (io_read_rsp_payload_fragment_data[255:0]         ), //i
    .io_writes_2_cmd_payload_mask     (memory_core_io_writes_2_cmd_payload_mask[31:0]   ), //i
    .io_writes_2_cmd_payload_context  (memory_core_io_writes_2_cmd_payload_context[8:0] ), //i
    .io_writes_2_rsp_valid            (memory_core_io_writes_2_rsp_valid                ), //o
    .io_writes_2_rsp_payload_context  (memory_core_io_writes_2_rsp_payload_context[8:0] ), //o
    .io_reads_0_cmd_valid             (memory_core_io_reads_0_cmd_valid                 ), //i
    .io_reads_0_cmd_ready             (memory_core_io_reads_0_cmd_ready                 ), //o
    .io_reads_0_cmd_payload_address   (memory_core_io_reads_0_cmd_payload_address[12:0] ), //i
    .io_reads_0_cmd_payload_priority  (channels_1_priority[1:0]                         ), //i
    .io_reads_0_cmd_payload_context   (memory_core_io_reads_0_cmd_payload_context[2:0]  ), //i
    .io_reads_0_rsp_valid             (memory_core_io_reads_0_rsp_valid                 ), //o
    .io_reads_0_rsp_ready             (io_outputs_0_ready                               ), //i
    .io_reads_0_rsp_payload_data      (memory_core_io_reads_0_rsp_payload_data[127:0]   ), //o
    .io_reads_0_rsp_payload_mask      (memory_core_io_reads_0_rsp_payload_mask[15:0]    ), //o
    .io_reads_0_rsp_payload_context   (memory_core_io_reads_0_rsp_payload_context[2:0]  ), //o
    .io_reads_1_cmd_valid             (memory_core_io_reads_1_cmd_valid                 ), //i
    .io_reads_1_cmd_ready             (memory_core_io_reads_1_cmd_ready                 ), //o
    .io_reads_1_cmd_payload_address   (memory_core_io_reads_1_cmd_payload_address[12:0] ), //i
    .io_reads_1_cmd_payload_priority  (channels_3_priority[1:0]                         ), //i
    .io_reads_1_cmd_payload_context   (memory_core_io_reads_1_cmd_payload_context[2:0]  ), //i
    .io_reads_1_rsp_valid             (memory_core_io_reads_1_rsp_valid                 ), //o
    .io_reads_1_rsp_ready             (io_outputs_1_ready                               ), //i
    .io_reads_1_rsp_payload_data      (memory_core_io_reads_1_rsp_payload_data[127:0]   ), //o
    .io_reads_1_rsp_payload_mask      (memory_core_io_reads_1_rsp_payload_mask[15:0]    ), //o
    .io_reads_1_rsp_payload_context   (memory_core_io_reads_1_rsp_payload_context[2:0]  ), //o
    .io_reads_2_cmd_valid             (b2m_fsm_sel_valid                                ), //i
    .io_reads_2_cmd_ready             (memory_core_io_reads_2_cmd_ready                 ), //o
    .io_reads_2_cmd_payload_address   (memory_core_io_reads_2_cmd_payload_address[12:0] ), //i
    .io_reads_2_cmd_payload_context   (memory_core_io_reads_2_cmd_payload_context[14:0] ), //i
    .io_reads_2_rsp_valid             (memory_core_io_reads_2_rsp_valid                 ), //o
    .io_reads_2_rsp_ready             (memory_core_io_reads_2_rsp_rValidN               ), //i
    .io_reads_2_rsp_payload_data      (memory_core_io_reads_2_rsp_payload_data[255:0]   ), //o
    .io_reads_2_rsp_payload_mask      (memory_core_io_reads_2_rsp_payload_mask[31:0]    ), //o
    .io_reads_2_rsp_payload_context   (memory_core_io_reads_2_rsp_payload_context[14:0] ), //o
    .clk                              (clk                                              ), //i
    .reset                            (reset                                            )  //i
  );
  EfxDMA_Aggregator b2m_fsm_aggregate_engine (
    .io_input_valid         (b2m_fsm_aggregate_memoryPort_valid                  ), //i
    .io_input_ready         (b2m_fsm_aggregate_engine_io_input_ready             ), //o
    .io_input_payload_data  (b2m_fsm_aggregate_memoryPort_payload_data[255:0]    ), //i
    .io_input_payload_mask  (b2m_fsm_aggregate_engine_io_input_payload_mask[31:0]), //i
    .io_output_data         (b2m_fsm_aggregate_engine_io_output_data[255:0]      ), //o
    .io_output_mask         (b2m_fsm_aggregate_engine_io_output_mask[31:0]       ), //o
    .io_output_enough       (b2m_fsm_cmd_enoughAggregation                       ), //i
    .io_output_consume      (io_write_cmd_fire                                   ), //i
    .io_output_consumed     (b2m_fsm_aggregate_engine_io_output_consumed         ), //o
    .io_output_lastByteUsed (b2m_fsm_cmd_maskLastTriggerReg[4:0]                 ), //i
    .io_output_usedUntil    (b2m_fsm_aggregate_engine_io_output_usedUntil[4:0]   ), //o
    .io_flush               (b2m_fsm_aggregate_engine_io_flush                   ), //i
    .io_offset              (b2m_fsm_aggregate_engine_io_offset[4:0]             ), //i
    .io_burstLength         (b2m_fsm_sel_bytesInBurst[12:0]                      ), //i
    .clk                    (clk                                                 ), //i
    .reset                  (reset                                               )  //i
  );
  always @(*) begin
    case(_zz_s2b_0_cmd_byteCount_11)
      3'b000 : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount;
      3'b001 : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount_1;
      3'b010 : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount_2;
      3'b011 : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount_3;
      3'b100 : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount_4;
      3'b101 : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount_5;
      3'b110 : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount_6;
      default : _zz_s2b_0_cmd_byteCount_10 = _zz_s2b_0_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_0_cmd_byteCount_13)
      3'b000 : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount;
      3'b001 : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount_1;
      3'b010 : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount_2;
      3'b011 : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount_3;
      3'b100 : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount_4;
      3'b101 : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount_5;
      3'b110 : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount_6;
      default : _zz_s2b_0_cmd_byteCount_12 = _zz_s2b_0_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_0_cmd_byteCount_16)
      3'b000 : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount;
      3'b001 : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount_1;
      3'b010 : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount_2;
      3'b011 : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount_3;
      3'b100 : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount_4;
      3'b101 : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount_5;
      3'b110 : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount_6;
      default : _zz_s2b_0_cmd_byteCount_15 = _zz_s2b_0_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_0_cmd_byteCount_18)
      3'b000 : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount;
      3'b001 : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount_1;
      3'b010 : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount_2;
      3'b011 : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount_3;
      3'b100 : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount_4;
      3'b101 : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount_5;
      3'b110 : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount_6;
      default : _zz_s2b_0_cmd_byteCount_17 = _zz_s2b_0_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_0_cmd_byteCount_21)
      3'b000 : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount;
      3'b001 : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount_1;
      3'b010 : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount_2;
      3'b011 : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount_3;
      3'b100 : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount_4;
      3'b101 : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount_5;
      3'b110 : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount_6;
      default : _zz_s2b_0_cmd_byteCount_20 = _zz_s2b_0_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_0_cmd_byteCount_23)
      3'b000 : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount;
      3'b001 : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount_1;
      3'b010 : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount_2;
      3'b011 : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount_3;
      3'b100 : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount_4;
      3'b101 : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount_5;
      3'b110 : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount_6;
      default : _zz_s2b_0_cmd_byteCount_22 = _zz_s2b_0_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_1_cmd_byteCount_11)
      3'b000 : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount;
      3'b001 : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount_1;
      3'b010 : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount_2;
      3'b011 : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount_3;
      3'b100 : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount_4;
      3'b101 : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount_5;
      3'b110 : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount_6;
      default : _zz_s2b_1_cmd_byteCount_10 = _zz_s2b_1_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_1_cmd_byteCount_13)
      3'b000 : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount;
      3'b001 : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount_1;
      3'b010 : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount_2;
      3'b011 : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount_3;
      3'b100 : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount_4;
      3'b101 : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount_5;
      3'b110 : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount_6;
      default : _zz_s2b_1_cmd_byteCount_12 = _zz_s2b_1_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_1_cmd_byteCount_16)
      3'b000 : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount;
      3'b001 : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount_1;
      3'b010 : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount_2;
      3'b011 : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount_3;
      3'b100 : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount_4;
      3'b101 : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount_5;
      3'b110 : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount_6;
      default : _zz_s2b_1_cmd_byteCount_15 = _zz_s2b_1_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_1_cmd_byteCount_18)
      3'b000 : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount;
      3'b001 : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount_1;
      3'b010 : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount_2;
      3'b011 : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount_3;
      3'b100 : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount_4;
      3'b101 : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount_5;
      3'b110 : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount_6;
      default : _zz_s2b_1_cmd_byteCount_17 = _zz_s2b_1_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_1_cmd_byteCount_21)
      3'b000 : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount;
      3'b001 : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount_1;
      3'b010 : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount_2;
      3'b011 : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount_3;
      3'b100 : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount_4;
      3'b101 : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount_5;
      3'b110 : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount_6;
      default : _zz_s2b_1_cmd_byteCount_20 = _zz_s2b_1_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_s2b_1_cmd_byteCount_23)
      3'b000 : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount;
      3'b001 : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount_1;
      3'b010 : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount_2;
      3'b011 : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount_3;
      3'b100 : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount_4;
      3'b101 : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount_5;
      3'b110 : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount_6;
      default : _zz_s2b_1_cmd_byteCount_22 = _zz_s2b_1_cmd_byteCount_7;
    endcase
  end

  always @(*) begin
    case(_zz_m2b_cmd_s0_priority_masked_2)
      2'b00 : _zz__zz_m2b_cmd_s0_priority_chosenOh_2_3 = m2b_cmd_s0_priority_roundRobins_0;
      2'b01 : _zz__zz_m2b_cmd_s0_priority_chosenOh_2_3 = m2b_cmd_s0_priority_roundRobins_1;
      2'b10 : _zz__zz_m2b_cmd_s0_priority_chosenOh_2_3 = m2b_cmd_s0_priority_roundRobins_2;
      default : _zz__zz_m2b_cmd_s0_priority_chosenOh_2_3 = m2b_cmd_s0_priority_roundRobins_3;
    endcase
  end

  always @(*) begin
    case(m2b_cmd_s0_priority_chosen)
      1'b0 : _zz_m2b_cmd_s0_priority_weightLast = (channels_1_weight == m2b_cmd_s0_priority_counter);
      default : _zz_m2b_cmd_s0_priority_weightLast = (channels_3_weight == m2b_cmd_s0_priority_counter);
    endcase
  end

  always @(*) begin
    case(m2b_cmd_s0_chosen)
      1'b0 : begin
        _zz_m2b_cmd_s0_address = channels_1_push_m2b_address;
        _zz_m2b_cmd_s0_bytesLeft = channels_1_push_m2b_bytesLeft;
        _zz_m2b_cmd_s0_lengthHead = channels_1_push_m2b_bytePerBurst;
      end
      default : begin
        _zz_m2b_cmd_s0_address = channels_3_push_m2b_address;
        _zz_m2b_cmd_s0_bytesLeft = channels_3_push_m2b_bytesLeft;
        _zz_m2b_cmd_s0_lengthHead = channels_3_push_m2b_bytePerBurst;
      end
    endcase
  end

  always @(*) begin
    case(m2b_rsp_context_channel)
      1'b0 : _zz_io_writes_2_cmd_payload_address = channels_1_fifo_push_ptrWithBase;
      default : _zz_io_writes_2_cmd_payload_address = channels_3_fifo_push_ptrWithBase;
    endcase
  end

  always @(*) begin
    case(_zz_b2m_fsm_arbiter_logic_priority_masked_2)
      2'b00 : _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_3 = b2m_fsm_arbiter_logic_priority_roundRobins_0;
      2'b01 : _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_3 = b2m_fsm_arbiter_logic_priority_roundRobins_1;
      2'b10 : _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_3 = b2m_fsm_arbiter_logic_priority_roundRobins_2;
      default : _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2_3 = b2m_fsm_arbiter_logic_priority_roundRobins_3;
    endcase
  end

  always @(*) begin
    case(b2m_fsm_arbiter_logic_priority_chosen)
      1'b0 : _zz_b2m_fsm_arbiter_logic_priority_weightLast = (channels_0_weight == b2m_fsm_arbiter_logic_priority_counter);
      default : _zz_b2m_fsm_arbiter_logic_priority_weightLast = (channels_2_weight == b2m_fsm_arbiter_logic_priority_counter);
    endcase
  end

  always @(*) begin
    case(b2m_fsm_arbiter_logic_chosen)
      1'b0 : begin
        _zz_b2m_fsm_sel_address = channels_0_pop_b2m_address;
        _zz_b2m_fsm_sel_ptr = channels_0_fifo_pop_ptrWithBase;
        _zz_b2m_fsm_sel_ptrMask = channels_0_fifo_words;
        _zz_b2m_fsm_sel_bytePerBurst = channels_0_pop_b2m_bytePerBurst;
        _zz_b2m_fsm_sel_bytesInFifo = channels_0_fifo_pop_bytes;
        _zz_b2m_fsm_sel_flush = channels_0_pop_b2m_flush;
        _zz_b2m_fsm_sel_packet = channels_0_pop_b2m_packet;
        _zz_b2m_fsm_sel_bytesLeft = channels_0_pop_b2m_bytesLeft;
      end
      default : begin
        _zz_b2m_fsm_sel_address = channels_2_pop_b2m_address;
        _zz_b2m_fsm_sel_ptr = channels_2_fifo_pop_ptrWithBase;
        _zz_b2m_fsm_sel_ptrMask = channels_2_fifo_words;
        _zz_b2m_fsm_sel_bytePerBurst = channels_2_pop_b2m_bytePerBurst;
        _zz_b2m_fsm_sel_bytesInFifo = channels_2_fifo_pop_bytes;
        _zz_b2m_fsm_sel_flush = channels_2_pop_b2m_flush;
        _zz_b2m_fsm_sel_packet = channels_2_pop_b2m_packet;
        _zz_b2m_fsm_sel_bytesLeft = channels_2_pop_b2m_bytesLeft;
      end
    endcase
  end

  always @(*) begin
    case(b2m_fsm_sel_channel)
      1'b0 : begin
        _zz_b2m_fsm_fetch_context_ptr = channels_0_fifo_pop_ptr;
        _zz_b2m_fsm_aggregate_bytesToSkip = channels_0_pop_b2m_bytesToSkip;
      end
      default : begin
        _zz_b2m_fsm_fetch_context_ptr = channels_2_fifo_pop_ptr;
        _zz_b2m_fsm_aggregate_bytesToSkip = channels_2_pop_b2m_bytesToSkip;
      end
    endcase
  end

  assign ctrl_readErrorFlag = 1'b0;
  assign ctrl_writeErrorFlag = 1'b0;
  assign io_ctrl_PREADY = 1'b1;
  always @(*) begin
    io_ctrl_PRDATA = 32'h0;
    case(io_ctrl_PADDR)
      14'h002c : begin
        io_ctrl_PRDATA[0 : 0] = channels_0_channelValid;
      end
      14'h0054 : begin
        io_ctrl_PRDATA[0 : 0] = channels_0_interrupts_completion_valid;
        io_ctrl_PRDATA[2 : 2] = channels_0_interrupts_onChannelCompletion_valid;
        io_ctrl_PRDATA[4 : 4] = channels_0_interrupts_s2mPacket_valid;
      end
      14'h00ac : begin
        io_ctrl_PRDATA[0 : 0] = channels_1_channelValid;
      end
      14'h00d4 : begin
        io_ctrl_PRDATA[0 : 0] = channels_1_interrupts_completion_valid;
        io_ctrl_PRDATA[2 : 2] = channels_1_interrupts_onChannelCompletion_valid;
      end
      14'h012c : begin
        io_ctrl_PRDATA[0 : 0] = channels_2_channelValid;
      end
      14'h0154 : begin
        io_ctrl_PRDATA[0 : 0] = channels_2_interrupts_completion_valid;
        io_ctrl_PRDATA[2 : 2] = channels_2_interrupts_onChannelCompletion_valid;
        io_ctrl_PRDATA[4 : 4] = channels_2_interrupts_s2mPacket_valid;
      end
      14'h01ac : begin
        io_ctrl_PRDATA[0 : 0] = channels_3_channelValid;
      end
      14'h01d4 : begin
        io_ctrl_PRDATA[0 : 0] = channels_3_interrupts_completion_valid;
        io_ctrl_PRDATA[2 : 2] = channels_3_interrupts_onChannelCompletion_valid;
      end
      default : begin
      end
    endcase
  end

  assign ctrl_askWrite = ((io_ctrl_PSEL[0] && io_ctrl_PENABLE) && io_ctrl_PWRITE);
  assign ctrl_askRead = ((io_ctrl_PSEL[0] && io_ctrl_PENABLE) && (! io_ctrl_PWRITE));
  assign ctrl_doWrite = (((io_ctrl_PSEL[0] && io_ctrl_PENABLE) && io_ctrl_PREADY) && io_ctrl_PWRITE);
  assign ctrl_doRead = (((io_ctrl_PSEL[0] && io_ctrl_PENABLE) && io_ctrl_PREADY) && (! io_ctrl_PWRITE));
  assign io_ctrl_PSLVERROR = ((ctrl_doWrite && ctrl_writeErrorFlag) || (ctrl_doRead && ctrl_readErrorFlag));
  always @(*) begin
    channels_0_channelStart = 1'b0;
    if(when_BusSlaveFactory_l377) begin
      if(when_BusSlaveFactory_l379) begin
        channels_0_channelStart = _zz_channels_0_channelStart[0];
      end
    end
  end

  always @(*) begin
    channels_0_channelCompletion = 1'b0;
    if(channels_0_channelValid) begin
      if(channels_0_channelStop) begin
        if(channels_0_readyToStop) begin
          channels_0_channelCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_0_descriptorStart = 1'b0;
    if(channels_0_ctrl_kick) begin
      channels_0_descriptorStart = 1'b1;
    end
    if(channels_0_channelValid) begin
      if(!channels_0_channelStop) begin
        if(when_DmaSg_l575) begin
          if(when_DmaSg_l578) begin
            channels_0_descriptorStart = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    channels_0_descriptorCompletion = 1'b0;
    if(channels_0_pop_b2m_packetSync) begin
      if(when_DmaSg_l532) begin
        if(channels_0_push_s2b_completionOnLast) begin
          channels_0_descriptorCompletion = 1'b1;
        end
      end
    end
    if(when_DmaSg_l547) begin
      channels_0_descriptorCompletion = 1'b1;
    end
    if(channels_0_channelValid) begin
      if(channels_0_channelStop) begin
        if(channels_0_readyToStop) begin
          channels_0_descriptorCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_0_readyToStop = 1'b1;
    if(when_DmaSg_l563) begin
      channels_0_readyToStop = 1'b0;
    end
  end

  assign channels_0_fifo_base = 14'h0;
  assign channels_0_fifo_words = 14'h007f;
  assign channels_0_fifo_push_availableDecr = 14'h0;
  assign channels_0_fifo_push_ptrWithBase = ((channels_0_fifo_base & (~ channels_0_fifo_words)) | (channels_0_fifo_push_ptr & channels_0_fifo_words));
  assign channels_0_fifo_pop_ptrWithBase = ((channels_0_fifo_base & (~ channels_0_fifo_words)) | (channels_0_fifo_pop_ptr & channels_0_fifo_words));
  assign channels_0_fifo_pop_empty = (channels_0_fifo_pop_ptr == channels_0_fifo_push_ptr);
  assign channels_0_fifo_pop_withOverride_backupNext = (_zz_channels_0_fifo_pop_withOverride_backupNext - channels_0_fifo_pop_bytesDecr_value);
  always @(*) begin
    channels_0_fifo_pop_withOverride_load = 1'b0;
    if(when_DmaSg_l457) begin
      channels_0_fifo_pop_withOverride_load = 1'b1;
    end
  end

  always @(*) begin
    channels_0_fifo_pop_withOverride_unload = 1'b0;
    if(channels_0_pop_b2m_packetSync) begin
      channels_0_fifo_pop_withOverride_unload = 1'b1;
    end
  end

  assign when_DmaSg_l409 = (channels_0_channelStart || channels_0_fifo_pop_withOverride_unload);
  assign channels_0_fifo_pop_bytes = channels_0_fifo_pop_withOverride_exposed;
  assign channels_0_fifo_empty = (channels_0_fifo_push_ptr == channels_0_fifo_pop_ptr);
  always @(*) begin
    channels_0_push_s2b_packetEvent = 1'b0;
    if(when_DmaSg_l679) begin
      channels_0_push_s2b_packetEvent = 1'b1;
    end
  end

  assign when_DmaSg_l457 = (channels_0_push_s2b_packetEvent && channels_0_push_s2b_completionOnLast);
  assign channels_0_pop_b2m_bytePerBurst = 13'h01ff;
  always @(*) begin
    channels_0_pop_b2m_fire = 1'b0;
    if(when_DmaSg_l935) begin
      if(_zz_1[0]) begin
        channels_0_pop_b2m_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    channels_0_pop_b2m_packetSync = 1'b0;
    if(when_DmaSg_l523) begin
      if(channels_0_pop_b2m_packet) begin
        channels_0_pop_b2m_packetSync = 1'b1;
      end
    end
    if(io_write_rsp_fire) begin
      if(when_DmaSg_l1116) begin
        if(b2m_rsp_context_doPacketSync) begin
          channels_0_pop_b2m_packetSync = 1'b1;
        end
      end
    end
  end

  assign when_DmaSg_l505 = (channels_0_channelStart || channels_0_pop_b2m_fire);
  always @(*) begin
    channels_0_pop_b2m_memRsp = 1'b0;
    if(io_write_rsp_fire) begin
      if(_zz_3[0]) begin
        channels_0_pop_b2m_memRsp = 1'b1;
      end
    end
  end

  assign channels_0_pop_b2m_selfFlush = (channels_0_pop_b2m_bytesLeft < _zz_channels_0_pop_b2m_selfFlush);
  assign channels_0_pop_b2m_request = ((((((channels_0_descriptorValid && (! channels_0_channelStop)) && (! channels_0_pop_b2m_waitFinalRsp)) && channels_0_pop_memory) && ((_zz_channels_0_pop_b2m_request < channels_0_fifo_pop_bytes) || (((channels_0_fifo_push_available < _zz_channels_0_pop_b2m_request_1) || channels_0_pop_b2m_flush) || channels_0_pop_b2m_selfFlush))) && (channels_0_fifo_pop_bytes != 18'h0)) && (channels_0_pop_b2m_memPending != 4'b1111));
  always @(*) begin
    channels_0_pop_b2m_memPendingInc = 1'b0;
    if(when_DmaSg_l758_1) begin
      if(when_DmaSg_l773_2) begin
        channels_0_pop_b2m_memPendingInc = 1'b1;
      end
    end
  end

  always @(*) begin
    channels_0_pop_b2m_decrBytes = 18'h0;
    if(b2m_fsm_s1) begin
      if(when_DmaSg_l996) begin
        channels_0_pop_b2m_decrBytes = {4'd0, b2m_fsm_bytesInBurstP1};
      end
    end
  end

  assign when_DmaSg_l523 = ((channels_0_pop_b2m_memPending == 4'b0000) && (channels_0_fifo_pop_bytes == 18'h0));
  assign when_DmaSg_l532 = (channels_0_descriptorValid && (! channels_0_push_memory));
  assign when_DmaSg_l547 = ((channels_0_descriptorValid && (channels_0_pop_b2m_memPending == 4'b0000)) && channels_0_pop_b2m_waitFinalRsp);
  assign when_DmaSg_l563 = (channels_0_pop_b2m_memPending != 4'b0000);
  assign channels_0_readyForChannelCompletion = 1'b1;
  assign when_DmaSg_l575 = (! channels_0_descriptorValid);
  always @(*) begin
    _zz_when_DmaSg_l593 = 1'b1;
    if(when_DmaSg_l578) begin
      _zz_when_DmaSg_l593 = 1'b0;
    end
    if(channels_0_ctrl_kick) begin
      _zz_when_DmaSg_l593 = 1'b0;
    end
  end

  assign when_DmaSg_l578 = (channels_0_selfRestart && (! channels_0_ctrl_kick));
  assign when_DmaSg_l593 = (_zz_when_DmaSg_l593 && channels_0_readyForChannelCompletion);
  assign channels_0_s2b_full = (channels_0_fifo_push_available < 14'h0002);
  assign when_DmaSg_l255 = (channels_0_descriptorValid && channels_0_descriptorCompletion);
  assign when_DmaSg_l255_1 = (! channels_0_interrupts_completion_enable);
  assign when_DmaSg_l255_2 = (channels_0_channelValid && channels_0_channelCompletion);
  assign when_DmaSg_l255_3 = (! channels_0_interrupts_onChannelCompletion_enable);
  assign when_DmaSg_l255_4 = (! channels_0_interrupts_s2mPacket_enable);
  always @(*) begin
    channels_1_channelStart = 1'b0;
    if(when_BusSlaveFactory_l377_2) begin
      if(when_BusSlaveFactory_l379_2) begin
        channels_1_channelStart = _zz_channels_1_channelStart[0];
      end
    end
  end

  always @(*) begin
    channels_1_channelCompletion = 1'b0;
    if(channels_1_channelValid) begin
      if(channels_1_channelStop) begin
        if(channels_1_readyToStop) begin
          channels_1_channelCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_1_descriptorStart = 1'b0;
    if(channels_1_ctrl_kick) begin
      channels_1_descriptorStart = 1'b1;
    end
    if(channels_1_channelValid) begin
      if(!channels_1_channelStop) begin
        if(when_DmaSg_l575_1) begin
          if(when_DmaSg_l578_1) begin
            channels_1_descriptorStart = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    channels_1_descriptorCompletion = 1'b0;
    if(when_DmaSg_l483) begin
      channels_1_descriptorCompletion = 1'b1;
    end
    if(channels_1_channelValid) begin
      if(channels_1_channelStop) begin
        if(channels_1_readyToStop) begin
          channels_1_descriptorCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_1_readyToStop = 1'b1;
    if(when_DmaSg_l562) begin
      channels_1_readyToStop = 1'b0;
    end
  end

  assign channels_1_fifo_base = 14'h0080;
  assign channels_1_fifo_words = 14'h007f;
  always @(*) begin
    channels_1_fifo_push_availableDecr = 14'h0;
    if(m2b_cmd_s1_valid) begin
      if(io_read_cmd_ready) begin
        if(when_DmaSg_l828) begin
          channels_1_fifo_push_availableDecr = {4'd0, m2b_cmd_s1_fifoPushDecr};
        end
      end
    end
  end

  assign channels_1_fifo_push_ptrWithBase = ((channels_1_fifo_base & (~ channels_1_fifo_words)) | (channels_1_fifo_push_ptr & channels_1_fifo_words));
  assign channels_1_fifo_pop_ptrWithBase = ((channels_1_fifo_base & (~ channels_1_fifo_words)) | (channels_1_fifo_pop_ptr & channels_1_fifo_words));
  assign channels_1_fifo_pop_empty = (channels_1_fifo_pop_ptr == channels_1_fifo_push_ptr);
  assign channels_1_fifo_pop_bytes = channels_1_fifo_pop_withoutOverride_exposed;
  assign channels_1_fifo_empty = (channels_1_fifo_push_ptr == channels_1_fifo_pop_ptr);
  assign channels_1_push_m2b_bytePerBurst = 13'h03ff;
  always @(*) begin
    channels_1_push_m2b_memPendingIncr = 1'b0;
    if(when_DmaSg_l758) begin
      if(when_DmaSg_l773) begin
        channels_1_push_m2b_memPendingIncr = 1'b1;
      end
    end
  end

  always @(*) begin
    channels_1_push_m2b_memPendingDecr = 1'b0;
    if(when_DmaSg_l893) begin
      channels_1_push_m2b_memPendingDecr = 1'b1;
    end
  end

  always @(*) begin
    channels_1_push_m2b_loadRequest = (((((channels_1_descriptorValid && (! channels_1_channelStop)) && (! channels_1_push_m2b_loadDone)) && channels_1_push_memory) && (_zz_channels_1_push_m2b_loadRequest < channels_1_fifo_push_available)) && (channels_1_push_m2b_memPending != 4'b1111));
    if(when_DmaSg_l486) begin
      channels_1_push_m2b_loadRequest = 1'b0;
    end
  end

  always @(*) begin
    channels_1_pop_b2s_veryLastTrigger = 1'b0;
    if(when_DmaSg_l847) begin
      if(when_DmaSg_l848) begin
        channels_1_pop_b2s_veryLastTrigger = 1'b1;
      end
    end
  end

  assign when_DmaSg_l474 = (channels_1_pop_b2s_veryLastTrigger && channels_1_pop_b2s_last);
  assign when_DmaSg_l483 = ((((channels_1_descriptorValid && (! channels_1_pop_memory)) && channels_1_push_memory) && channels_1_push_m2b_loadDone) && (channels_1_push_m2b_memPending == 4'b0000));
  assign when_DmaSg_l486 = (((! channels_1_pop_memory) && channels_1_pop_b2s_veryLastValid) && (channels_1_push_m2b_bytesLeft <= _zz_when_DmaSg_l486));
  assign when_DmaSg_l562 = (channels_1_push_m2b_memPending != 4'b0000);
  always @(*) begin
    channels_1_readyForChannelCompletion = 1'b1;
    if(when_DmaSg_l566) begin
      channels_1_readyForChannelCompletion = 1'b0;
    end
  end

  assign when_DmaSg_l566 = ((! channels_1_pop_memory) && (! channels_1_fifo_pop_empty));
  assign when_DmaSg_l575_1 = (! channels_1_descriptorValid);
  always @(*) begin
    _zz_when_DmaSg_l593_1 = 1'b1;
    if(when_DmaSg_l578_1) begin
      _zz_when_DmaSg_l593_1 = 1'b0;
    end
    if(channels_1_ctrl_kick) begin
      _zz_when_DmaSg_l593_1 = 1'b0;
    end
  end

  assign when_DmaSg_l578_1 = (channels_1_selfRestart && (! channels_1_ctrl_kick));
  assign when_DmaSg_l593_1 = (_zz_when_DmaSg_l593_1 && channels_1_readyForChannelCompletion);
  assign channels_1_s2b_full = (channels_1_fifo_push_available < 14'h0002);
  assign when_DmaSg_l255_5 = (channels_1_descriptorValid && channels_1_descriptorCompletion);
  assign when_DmaSg_l255_6 = (! channels_1_interrupts_completion_enable);
  assign when_DmaSg_l255_7 = (channels_1_channelValid && channels_1_channelCompletion);
  assign when_DmaSg_l255_8 = (! channels_1_interrupts_onChannelCompletion_enable);
  always @(*) begin
    channels_2_channelStart = 1'b0;
    if(when_BusSlaveFactory_l377_4) begin
      if(when_BusSlaveFactory_l379_4) begin
        channels_2_channelStart = _zz_channels_2_channelStart[0];
      end
    end
  end

  always @(*) begin
    channels_2_channelCompletion = 1'b0;
    if(channels_2_channelValid) begin
      if(channels_2_channelStop) begin
        if(channels_2_readyToStop) begin
          channels_2_channelCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_2_descriptorStart = 1'b0;
    if(channels_2_ctrl_kick) begin
      channels_2_descriptorStart = 1'b1;
    end
    if(channels_2_channelValid) begin
      if(!channels_2_channelStop) begin
        if(when_DmaSg_l575_2) begin
          if(when_DmaSg_l578_2) begin
            channels_2_descriptorStart = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    channels_2_descriptorCompletion = 1'b0;
    if(channels_2_pop_b2m_packetSync) begin
      if(when_DmaSg_l532_1) begin
        if(channels_2_push_s2b_completionOnLast) begin
          channels_2_descriptorCompletion = 1'b1;
        end
      end
    end
    if(when_DmaSg_l547_1) begin
      channels_2_descriptorCompletion = 1'b1;
    end
    if(channels_2_channelValid) begin
      if(channels_2_channelStop) begin
        if(channels_2_readyToStop) begin
          channels_2_descriptorCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_2_readyToStop = 1'b1;
    if(when_DmaSg_l563_1) begin
      channels_2_readyToStop = 1'b0;
    end
  end

  assign channels_2_fifo_base = 14'h0100;
  assign channels_2_fifo_words = 14'h007f;
  assign channels_2_fifo_push_availableDecr = 14'h0;
  assign channels_2_fifo_push_ptrWithBase = ((channels_2_fifo_base & (~ channels_2_fifo_words)) | (channels_2_fifo_push_ptr & channels_2_fifo_words));
  assign channels_2_fifo_pop_ptrWithBase = ((channels_2_fifo_base & (~ channels_2_fifo_words)) | (channels_2_fifo_pop_ptr & channels_2_fifo_words));
  assign channels_2_fifo_pop_empty = (channels_2_fifo_pop_ptr == channels_2_fifo_push_ptr);
  assign channels_2_fifo_pop_withOverride_backupNext = (_zz_channels_2_fifo_pop_withOverride_backupNext - channels_2_fifo_pop_bytesDecr_value);
  always @(*) begin
    channels_2_fifo_pop_withOverride_load = 1'b0;
    if(when_DmaSg_l457_1) begin
      channels_2_fifo_pop_withOverride_load = 1'b1;
    end
  end

  always @(*) begin
    channels_2_fifo_pop_withOverride_unload = 1'b0;
    if(channels_2_pop_b2m_packetSync) begin
      channels_2_fifo_pop_withOverride_unload = 1'b1;
    end
  end

  assign when_DmaSg_l409_1 = (channels_2_channelStart || channels_2_fifo_pop_withOverride_unload);
  assign channels_2_fifo_pop_bytes = channels_2_fifo_pop_withOverride_exposed;
  assign channels_2_fifo_empty = (channels_2_fifo_push_ptr == channels_2_fifo_pop_ptr);
  always @(*) begin
    channels_2_push_s2b_packetEvent = 1'b0;
    if(when_DmaSg_l679_1) begin
      channels_2_push_s2b_packetEvent = 1'b1;
    end
  end

  assign when_DmaSg_l457_1 = (channels_2_push_s2b_packetEvent && channels_2_push_s2b_completionOnLast);
  assign channels_2_pop_b2m_bytePerBurst = 13'h01ff;
  always @(*) begin
    channels_2_pop_b2m_fire = 1'b0;
    if(when_DmaSg_l935) begin
      if(_zz_1[1]) begin
        channels_2_pop_b2m_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    channels_2_pop_b2m_packetSync = 1'b0;
    if(when_DmaSg_l523_1) begin
      if(channels_2_pop_b2m_packet) begin
        channels_2_pop_b2m_packetSync = 1'b1;
      end
    end
    if(io_write_rsp_fire) begin
      if(when_DmaSg_l1116_1) begin
        if(b2m_rsp_context_doPacketSync) begin
          channels_2_pop_b2m_packetSync = 1'b1;
        end
      end
    end
  end

  assign when_DmaSg_l505_1 = (channels_2_channelStart || channels_2_pop_b2m_fire);
  always @(*) begin
    channels_2_pop_b2m_memRsp = 1'b0;
    if(io_write_rsp_fire) begin
      if(_zz_3[1]) begin
        channels_2_pop_b2m_memRsp = 1'b1;
      end
    end
  end

  assign channels_2_pop_b2m_selfFlush = (channels_2_pop_b2m_bytesLeft < _zz_channels_2_pop_b2m_selfFlush);
  assign channels_2_pop_b2m_request = ((((((channels_2_descriptorValid && (! channels_2_channelStop)) && (! channels_2_pop_b2m_waitFinalRsp)) && channels_2_pop_memory) && ((_zz_channels_2_pop_b2m_request < channels_2_fifo_pop_bytes) || (((channels_2_fifo_push_available < _zz_channels_2_pop_b2m_request_1) || channels_2_pop_b2m_flush) || channels_2_pop_b2m_selfFlush))) && (channels_2_fifo_pop_bytes != 18'h0)) && (channels_2_pop_b2m_memPending != 4'b1111));
  always @(*) begin
    channels_2_pop_b2m_memPendingInc = 1'b0;
    if(when_DmaSg_l758_1) begin
      if(when_DmaSg_l773_3) begin
        channels_2_pop_b2m_memPendingInc = 1'b1;
      end
    end
  end

  always @(*) begin
    channels_2_pop_b2m_decrBytes = 18'h0;
    if(b2m_fsm_s1) begin
      if(when_DmaSg_l996_1) begin
        channels_2_pop_b2m_decrBytes = {4'd0, b2m_fsm_bytesInBurstP1};
      end
    end
  end

  assign when_DmaSg_l523_1 = ((channels_2_pop_b2m_memPending == 4'b0000) && (channels_2_fifo_pop_bytes == 18'h0));
  assign when_DmaSg_l532_1 = (channels_2_descriptorValid && (! channels_2_push_memory));
  assign when_DmaSg_l547_1 = ((channels_2_descriptorValid && (channels_2_pop_b2m_memPending == 4'b0000)) && channels_2_pop_b2m_waitFinalRsp);
  assign when_DmaSg_l563_1 = (channels_2_pop_b2m_memPending != 4'b0000);
  assign channels_2_readyForChannelCompletion = 1'b1;
  assign when_DmaSg_l575_2 = (! channels_2_descriptorValid);
  always @(*) begin
    _zz_when_DmaSg_l593_2 = 1'b1;
    if(when_DmaSg_l578_2) begin
      _zz_when_DmaSg_l593_2 = 1'b0;
    end
    if(channels_2_ctrl_kick) begin
      _zz_when_DmaSg_l593_2 = 1'b0;
    end
  end

  assign when_DmaSg_l578_2 = (channels_2_selfRestart && (! channels_2_ctrl_kick));
  assign when_DmaSg_l593_2 = (_zz_when_DmaSg_l593_2 && channels_2_readyForChannelCompletion);
  assign channels_2_s2b_full = (channels_2_fifo_push_available < 14'h0002);
  assign when_DmaSg_l255_9 = (channels_2_descriptorValid && channels_2_descriptorCompletion);
  assign when_DmaSg_l255_10 = (! channels_2_interrupts_completion_enable);
  assign when_DmaSg_l255_11 = (channels_2_channelValid && channels_2_channelCompletion);
  assign when_DmaSg_l255_12 = (! channels_2_interrupts_onChannelCompletion_enable);
  assign when_DmaSg_l255_13 = (! channels_2_interrupts_s2mPacket_enable);
  always @(*) begin
    channels_3_channelStart = 1'b0;
    if(when_BusSlaveFactory_l377_6) begin
      if(when_BusSlaveFactory_l379_6) begin
        channels_3_channelStart = _zz_channels_3_channelStart[0];
      end
    end
  end

  always @(*) begin
    channels_3_channelCompletion = 1'b0;
    if(channels_3_channelValid) begin
      if(channels_3_channelStop) begin
        if(channels_3_readyToStop) begin
          channels_3_channelCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_3_descriptorStart = 1'b0;
    if(channels_3_ctrl_kick) begin
      channels_3_descriptorStart = 1'b1;
    end
    if(channels_3_channelValid) begin
      if(!channels_3_channelStop) begin
        if(when_DmaSg_l575_3) begin
          if(when_DmaSg_l578_3) begin
            channels_3_descriptorStart = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    channels_3_descriptorCompletion = 1'b0;
    if(when_DmaSg_l483_1) begin
      channels_3_descriptorCompletion = 1'b1;
    end
    if(channels_3_channelValid) begin
      if(channels_3_channelStop) begin
        if(channels_3_readyToStop) begin
          channels_3_descriptorCompletion = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    channels_3_readyToStop = 1'b1;
    if(when_DmaSg_l562_1) begin
      channels_3_readyToStop = 1'b0;
    end
  end

  assign channels_3_fifo_base = 14'h0180;
  assign channels_3_fifo_words = 14'h007f;
  always @(*) begin
    channels_3_fifo_push_availableDecr = 14'h0;
    if(m2b_cmd_s1_valid) begin
      if(io_read_cmd_ready) begin
        if(when_DmaSg_l828_1) begin
          channels_3_fifo_push_availableDecr = {4'd0, m2b_cmd_s1_fifoPushDecr};
        end
      end
    end
  end

  assign channels_3_fifo_push_ptrWithBase = ((channels_3_fifo_base & (~ channels_3_fifo_words)) | (channels_3_fifo_push_ptr & channels_3_fifo_words));
  assign channels_3_fifo_pop_ptrWithBase = ((channels_3_fifo_base & (~ channels_3_fifo_words)) | (channels_3_fifo_pop_ptr & channels_3_fifo_words));
  assign channels_3_fifo_pop_empty = (channels_3_fifo_pop_ptr == channels_3_fifo_push_ptr);
  assign channels_3_fifo_pop_bytes = channels_3_fifo_pop_withoutOverride_exposed;
  assign channels_3_fifo_empty = (channels_3_fifo_push_ptr == channels_3_fifo_pop_ptr);
  assign channels_3_push_m2b_bytePerBurst = 13'h01ff;
  always @(*) begin
    channels_3_push_m2b_memPendingIncr = 1'b0;
    if(when_DmaSg_l758) begin
      if(when_DmaSg_l773_1) begin
        channels_3_push_m2b_memPendingIncr = 1'b1;
      end
    end
  end

  always @(*) begin
    channels_3_push_m2b_memPendingDecr = 1'b0;
    if(when_DmaSg_l893_1) begin
      channels_3_push_m2b_memPendingDecr = 1'b1;
    end
  end

  always @(*) begin
    channels_3_push_m2b_loadRequest = (((((channels_3_descriptorValid && (! channels_3_channelStop)) && (! channels_3_push_m2b_loadDone)) && channels_3_push_memory) && (_zz_channels_3_push_m2b_loadRequest < channels_3_fifo_push_available)) && (channels_3_push_m2b_memPending != 4'b1111));
    if(when_DmaSg_l486_1) begin
      channels_3_push_m2b_loadRequest = 1'b0;
    end
  end

  always @(*) begin
    channels_3_pop_b2s_veryLastTrigger = 1'b0;
    if(when_DmaSg_l847) begin
      if(when_DmaSg_l848_1) begin
        channels_3_pop_b2s_veryLastTrigger = 1'b1;
      end
    end
  end

  assign when_DmaSg_l474_1 = (channels_3_pop_b2s_veryLastTrigger && channels_3_pop_b2s_last);
  assign when_DmaSg_l483_1 = ((((channels_3_descriptorValid && (! channels_3_pop_memory)) && channels_3_push_memory) && channels_3_push_m2b_loadDone) && (channels_3_push_m2b_memPending == 4'b0000));
  assign when_DmaSg_l486_1 = (((! channels_3_pop_memory) && channels_3_pop_b2s_veryLastValid) && (channels_3_push_m2b_bytesLeft <= _zz_when_DmaSg_l486_1));
  assign when_DmaSg_l562_1 = (channels_3_push_m2b_memPending != 4'b0000);
  always @(*) begin
    channels_3_readyForChannelCompletion = 1'b1;
    if(when_DmaSg_l566_1) begin
      channels_3_readyForChannelCompletion = 1'b0;
    end
  end

  assign when_DmaSg_l566_1 = ((! channels_3_pop_memory) && (! channels_3_fifo_pop_empty));
  assign when_DmaSg_l575_3 = (! channels_3_descriptorValid);
  always @(*) begin
    _zz_when_DmaSg_l593_3 = 1'b1;
    if(when_DmaSg_l578_3) begin
      _zz_when_DmaSg_l593_3 = 1'b0;
    end
    if(channels_3_ctrl_kick) begin
      _zz_when_DmaSg_l593_3 = 1'b0;
    end
  end

  assign when_DmaSg_l578_3 = (channels_3_selfRestart && (! channels_3_ctrl_kick));
  assign when_DmaSg_l593_3 = (_zz_when_DmaSg_l593_3 && channels_3_readyForChannelCompletion);
  assign channels_3_s2b_full = (channels_3_fifo_push_available < 14'h0002);
  assign when_DmaSg_l255_14 = (channels_3_descriptorValid && channels_3_descriptorCompletion);
  assign when_DmaSg_l255_15 = (! channels_3_interrupts_completion_enable);
  assign when_DmaSg_l255_16 = (channels_3_channelValid && channels_3_channelCompletion);
  assign when_DmaSg_l255_17 = (! channels_3_interrupts_onChannelCompletion_enable);
  assign io_inputs_0_fire = (io_inputs_0_valid && io_inputs_0_ready);
  assign when_package_l12 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0000));
  assign when_package_l12_1 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0001));
  assign when_package_l12_2 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0010));
  assign when_package_l12_3 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0011));
  assign when_package_l12_4 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0100));
  assign when_package_l12_5 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0101));
  assign when_package_l12_6 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0110));
  assign when_package_l12_7 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b0111));
  assign when_package_l12_8 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1000));
  assign when_package_l12_9 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1001));
  assign when_package_l12_10 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1010));
  assign when_package_l12_11 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1011));
  assign when_package_l12_12 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1100));
  assign when_package_l12_13 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1101));
  assign when_package_l12_14 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1110));
  assign when_package_l12_15 = (io_inputs_0_fire && (io_inputs_0_payload_sink == 4'b1111));
  assign s2b_0_cmd_firsts = {io_inputs_0_payload_last_regNextWhen_15,{io_inputs_0_payload_last_regNextWhen_14,{io_inputs_0_payload_last_regNextWhen_13,{io_inputs_0_payload_last_regNextWhen_12,{io_inputs_0_payload_last_regNextWhen_11,{io_inputs_0_payload_last_regNextWhen_10,{io_inputs_0_payload_last_regNextWhen_9,{io_inputs_0_payload_last_regNextWhen_8,{io_inputs_0_payload_last_regNextWhen_7,{io_inputs_0_payload_last_regNextWhen_6,{_zz_s2b_0_cmd_firsts,_zz_s2b_0_cmd_firsts_1}}}}}}}}}}};
  assign s2b_0_cmd_first = s2b_0_cmd_firsts[io_inputs_0_payload_sink];
  assign s2b_0_cmd_channelsOh = ((((channels_0_channelValid && (s2b_0_cmd_first || (! channels_0_push_s2b_waitFirst))) && (! channels_0_push_memory)) && 1'b1) && (io_inputs_0_payload_sink == 4'b0000));
  assign s2b_0_cmd_noHit = (! (|s2b_0_cmd_channelsOh));
  assign s2b_0_cmd_channelsFull = (channels_0_s2b_full || (channels_0_push_s2b_packetLock && io_inputs_0_payload_last));
  always @(*) begin
    io_inputs_0_thrown_valid = io_inputs_0_valid;
    if(s2b_0_cmd_noHit) begin
      io_inputs_0_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    io_inputs_0_ready = io_inputs_0_thrown_ready;
    if(s2b_0_cmd_noHit) begin
      io_inputs_0_ready = 1'b1;
    end
  end

  assign io_inputs_0_thrown_payload_data = io_inputs_0_payload_data;
  assign io_inputs_0_thrown_payload_mask = io_inputs_0_payload_mask;
  assign io_inputs_0_thrown_payload_sink = io_inputs_0_payload_sink;
  assign io_inputs_0_thrown_payload_last = io_inputs_0_payload_last;
  assign _zz_io_inputs_0_thrown_ready = (! (|(s2b_0_cmd_channelsOh & s2b_0_cmd_channelsFull)));
  assign s2b_0_cmd_sinkHalted_valid = (io_inputs_0_thrown_valid && _zz_io_inputs_0_thrown_ready);
  assign io_inputs_0_thrown_ready = (s2b_0_cmd_sinkHalted_ready && _zz_io_inputs_0_thrown_ready);
  assign s2b_0_cmd_sinkHalted_payload_data = io_inputs_0_thrown_payload_data;
  assign s2b_0_cmd_sinkHalted_payload_mask = io_inputs_0_thrown_payload_mask;
  assign s2b_0_cmd_sinkHalted_payload_sink = io_inputs_0_thrown_payload_sink;
  assign s2b_0_cmd_sinkHalted_payload_last = io_inputs_0_thrown_payload_last;
  assign _zz_s2b_0_cmd_byteCount = 5'h0;
  assign _zz_s2b_0_cmd_byteCount_1 = 5'h01;
  assign _zz_s2b_0_cmd_byteCount_2 = 5'h01;
  assign _zz_s2b_0_cmd_byteCount_3 = 5'h02;
  assign _zz_s2b_0_cmd_byteCount_4 = 5'h01;
  assign _zz_s2b_0_cmd_byteCount_5 = 5'h02;
  assign _zz_s2b_0_cmd_byteCount_6 = 5'h02;
  assign _zz_s2b_0_cmd_byteCount_7 = 5'h03;
  assign s2b_0_cmd_byteCount = (_zz_s2b_0_cmd_byteCount_8 + _zz_s2b_0_cmd_byteCount_19);
  assign s2b_0_cmd_context_channel = s2b_0_cmd_channelsOh;
  assign s2b_0_cmd_context_bytes = s2b_0_cmd_byteCount;
  assign s2b_0_cmd_context_flush = io_inputs_0_payload_last;
  assign s2b_0_cmd_context_packet = io_inputs_0_payload_last;
  assign s2b_0_cmd_sinkHalted_ready = memory_core_io_writes_0_cmd_ready;
  assign memory_core_io_writes_0_cmd_payload_address = channels_0_fifo_push_ptrWithBase[12:0];
  assign memory_core_io_writes_0_cmd_payload_context = {s2b_0_cmd_context_packet,{s2b_0_cmd_context_flush,{s2b_0_cmd_context_bytes,s2b_0_cmd_context_channel}}};
  assign memory_core_io_writes_0_cmd_fire = (s2b_0_cmd_sinkHalted_valid && memory_core_io_writes_0_cmd_ready);
  assign when_DmaSg_l665 = (s2b_0_cmd_channelsOh[0] && memory_core_io_writes_0_cmd_fire);
  assign _zz_s2b_0_rsp_context_channel = memory_core_io_writes_0_rsp_payload_context;
  assign s2b_0_rsp_context_channel = _zz_s2b_0_rsp_context_channel[0 : 0];
  assign s2b_0_rsp_context_bytes = _zz_s2b_0_rsp_context_channel[5 : 1];
  assign s2b_0_rsp_context_flush = _zz_s2b_0_rsp_context_channel[6];
  assign s2b_0_rsp_context_packet = _zz_s2b_0_rsp_context_channel[7];
  assign _zz_channels_0_fifo_pop_bytesIncr_value = (memory_core_io_writes_0_rsp_valid && s2b_0_rsp_context_channel[0]);
  assign when_DmaSg_l679 = (_zz_channels_0_fifo_pop_bytesIncr_value && s2b_0_rsp_context_packet);
  assign when_DmaSg_l681 = (_zz_channels_0_fifo_pop_bytesIncr_value && s2b_0_rsp_context_flush);
  assign when_DmaSg_l682 = (_zz_channels_0_fifo_pop_bytesIncr_value && s2b_0_rsp_context_packet);
  assign io_inputs_1_fire = (io_inputs_1_valid && io_inputs_1_ready);
  assign when_package_l12_16 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0000));
  assign when_package_l12_17 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0001));
  assign when_package_l12_18 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0010));
  assign when_package_l12_19 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0011));
  assign when_package_l12_20 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0100));
  assign when_package_l12_21 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0101));
  assign when_package_l12_22 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0110));
  assign when_package_l12_23 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b0111));
  assign when_package_l12_24 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1000));
  assign when_package_l12_25 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1001));
  assign when_package_l12_26 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1010));
  assign when_package_l12_27 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1011));
  assign when_package_l12_28 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1100));
  assign when_package_l12_29 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1101));
  assign when_package_l12_30 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1110));
  assign when_package_l12_31 = (io_inputs_1_fire && (io_inputs_1_payload_sink == 4'b1111));
  assign s2b_1_cmd_firsts = {io_inputs_1_payload_last_regNextWhen_15,{io_inputs_1_payload_last_regNextWhen_14,{io_inputs_1_payload_last_regNextWhen_13,{io_inputs_1_payload_last_regNextWhen_12,{io_inputs_1_payload_last_regNextWhen_11,{io_inputs_1_payload_last_regNextWhen_10,{io_inputs_1_payload_last_regNextWhen_9,{io_inputs_1_payload_last_regNextWhen_8,{io_inputs_1_payload_last_regNextWhen_7,{io_inputs_1_payload_last_regNextWhen_6,{_zz_s2b_1_cmd_firsts,_zz_s2b_1_cmd_firsts_1}}}}}}}}}}};
  assign s2b_1_cmd_first = s2b_1_cmd_firsts[io_inputs_1_payload_sink];
  assign s2b_1_cmd_channelsOh = ((((channels_2_channelValid && (s2b_1_cmd_first || (! channels_2_push_s2b_waitFirst))) && (! channels_2_push_memory)) && 1'b1) && (io_inputs_1_payload_sink == 4'b0000));
  assign s2b_1_cmd_noHit = (! (|s2b_1_cmd_channelsOh));
  assign s2b_1_cmd_channelsFull = (channels_2_s2b_full || (channels_2_push_s2b_packetLock && io_inputs_1_payload_last));
  always @(*) begin
    io_inputs_1_thrown_valid = io_inputs_1_valid;
    if(s2b_1_cmd_noHit) begin
      io_inputs_1_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    io_inputs_1_ready = io_inputs_1_thrown_ready;
    if(s2b_1_cmd_noHit) begin
      io_inputs_1_ready = 1'b1;
    end
  end

  assign io_inputs_1_thrown_payload_data = io_inputs_1_payload_data;
  assign io_inputs_1_thrown_payload_mask = io_inputs_1_payload_mask;
  assign io_inputs_1_thrown_payload_sink = io_inputs_1_payload_sink;
  assign io_inputs_1_thrown_payload_last = io_inputs_1_payload_last;
  assign _zz_io_inputs_1_thrown_ready = (! (|(s2b_1_cmd_channelsOh & s2b_1_cmd_channelsFull)));
  assign s2b_1_cmd_sinkHalted_valid = (io_inputs_1_thrown_valid && _zz_io_inputs_1_thrown_ready);
  assign io_inputs_1_thrown_ready = (s2b_1_cmd_sinkHalted_ready && _zz_io_inputs_1_thrown_ready);
  assign s2b_1_cmd_sinkHalted_payload_data = io_inputs_1_thrown_payload_data;
  assign s2b_1_cmd_sinkHalted_payload_mask = io_inputs_1_thrown_payload_mask;
  assign s2b_1_cmd_sinkHalted_payload_sink = io_inputs_1_thrown_payload_sink;
  assign s2b_1_cmd_sinkHalted_payload_last = io_inputs_1_thrown_payload_last;
  assign _zz_s2b_1_cmd_byteCount = 5'h0;
  assign _zz_s2b_1_cmd_byteCount_1 = 5'h01;
  assign _zz_s2b_1_cmd_byteCount_2 = 5'h01;
  assign _zz_s2b_1_cmd_byteCount_3 = 5'h02;
  assign _zz_s2b_1_cmd_byteCount_4 = 5'h01;
  assign _zz_s2b_1_cmd_byteCount_5 = 5'h02;
  assign _zz_s2b_1_cmd_byteCount_6 = 5'h02;
  assign _zz_s2b_1_cmd_byteCount_7 = 5'h03;
  assign s2b_1_cmd_byteCount = (_zz_s2b_1_cmd_byteCount_8 + _zz_s2b_1_cmd_byteCount_19);
  assign s2b_1_cmd_context_channel = s2b_1_cmd_channelsOh;
  assign s2b_1_cmd_context_bytes = s2b_1_cmd_byteCount;
  assign s2b_1_cmd_context_flush = io_inputs_1_payload_last;
  assign s2b_1_cmd_context_packet = io_inputs_1_payload_last;
  assign s2b_1_cmd_sinkHalted_ready = memory_core_io_writes_1_cmd_ready;
  assign memory_core_io_writes_1_cmd_payload_address = channels_2_fifo_push_ptrWithBase[12:0];
  assign memory_core_io_writes_1_cmd_payload_context = {s2b_1_cmd_context_packet,{s2b_1_cmd_context_flush,{s2b_1_cmd_context_bytes,s2b_1_cmd_context_channel}}};
  assign memory_core_io_writes_1_cmd_fire = (s2b_1_cmd_sinkHalted_valid && memory_core_io_writes_1_cmd_ready);
  assign when_DmaSg_l665_1 = (s2b_1_cmd_channelsOh[0] && memory_core_io_writes_1_cmd_fire);
  assign _zz_s2b_1_rsp_context_channel = memory_core_io_writes_1_rsp_payload_context;
  assign s2b_1_rsp_context_channel = _zz_s2b_1_rsp_context_channel[0 : 0];
  assign s2b_1_rsp_context_bytes = _zz_s2b_1_rsp_context_channel[5 : 1];
  assign s2b_1_rsp_context_flush = _zz_s2b_1_rsp_context_channel[6];
  assign s2b_1_rsp_context_packet = _zz_s2b_1_rsp_context_channel[7];
  assign _zz_channels_2_fifo_pop_bytesIncr_value = (memory_core_io_writes_1_rsp_valid && s2b_1_rsp_context_channel[0]);
  assign when_DmaSg_l679_1 = (_zz_channels_2_fifo_pop_bytesIncr_value && s2b_1_rsp_context_packet);
  assign when_DmaSg_l681_1 = (_zz_channels_2_fifo_pop_bytesIncr_value && s2b_1_rsp_context_flush);
  assign when_DmaSg_l682_1 = (_zz_channels_2_fifo_pop_bytesIncr_value && s2b_1_rsp_context_packet);
  assign b2s_0_cmd_channelsOh = (((channels_1_channelValid && (! channels_1_pop_memory)) && (channels_1_pop_b2s_portId == 1'b0)) && (! channels_1_fifo_pop_empty));
  assign b2s_0_cmd_veryLastPtr = channels_1_pop_b2s_veryLastPtr;
  assign b2s_0_cmd_address = channels_1_fifo_pop_ptrWithBase;
  assign b2s_0_cmd_context_channel = b2s_0_cmd_channelsOh;
  assign b2s_0_cmd_context_veryLast = ((channels_1_pop_b2s_veryLastValid && (b2s_0_cmd_address[13 : 1] == b2s_0_cmd_veryLastPtr[13 : 1])) && (b2s_0_cmd_address[0 : 0] == 1'b1));
  assign b2s_0_cmd_context_endPacket = channels_1_pop_b2s_veryLastEndPacket;
  assign memory_core_io_reads_0_cmd_valid = (|b2s_0_cmd_channelsOh);
  assign memory_core_io_reads_0_cmd_payload_address = b2s_0_cmd_address[12:0];
  assign memory_core_io_reads_0_cmd_payload_context = {b2s_0_cmd_context_endPacket,{b2s_0_cmd_context_veryLast,b2s_0_cmd_context_channel}};
  assign _zz_b2s_0_rsp_context_channel = memory_core_io_reads_0_rsp_payload_context;
  assign b2s_0_rsp_context_channel = _zz_b2s_0_rsp_context_channel[0 : 0];
  assign b2s_0_rsp_context_veryLast = _zz_b2s_0_rsp_context_channel[1];
  assign b2s_0_rsp_context_endPacket = _zz_b2s_0_rsp_context_channel[2];
  assign io_outputs_0_valid = memory_core_io_reads_0_rsp_valid;
  assign io_outputs_0_payload_data = memory_core_io_reads_0_rsp_payload_data;
  assign io_outputs_0_payload_mask = memory_core_io_reads_0_rsp_payload_mask;
  assign io_outputs_0_payload_sink = channels_1_pop_b2s_sinkId;
  assign io_outputs_0_payload_last = (b2s_0_rsp_context_veryLast && b2s_0_rsp_context_endPacket);
  assign io_outputs_0_fire = (io_outputs_0_valid && io_outputs_0_ready);
  assign when_DmaSg_l725 = (io_outputs_0_fire && b2s_0_rsp_context_veryLast);
  assign when_DmaSg_l726 = b2s_0_rsp_context_channel[0];
  assign b2s_1_cmd_channelsOh = (((channels_3_channelValid && (! channels_3_pop_memory)) && (channels_3_pop_b2s_portId == 1'b0)) && (! channels_3_fifo_pop_empty));
  assign b2s_1_cmd_veryLastPtr = channels_3_pop_b2s_veryLastPtr;
  assign b2s_1_cmd_address = channels_3_fifo_pop_ptrWithBase;
  assign b2s_1_cmd_context_channel = b2s_1_cmd_channelsOh;
  assign b2s_1_cmd_context_veryLast = ((channels_3_pop_b2s_veryLastValid && (b2s_1_cmd_address[13 : 1] == b2s_1_cmd_veryLastPtr[13 : 1])) && (b2s_1_cmd_address[0 : 0] == 1'b1));
  assign b2s_1_cmd_context_endPacket = channels_3_pop_b2s_veryLastEndPacket;
  assign memory_core_io_reads_1_cmd_valid = (|b2s_1_cmd_channelsOh);
  assign memory_core_io_reads_1_cmd_payload_address = b2s_1_cmd_address[12:0];
  assign memory_core_io_reads_1_cmd_payload_context = {b2s_1_cmd_context_endPacket,{b2s_1_cmd_context_veryLast,b2s_1_cmd_context_channel}};
  assign _zz_b2s_1_rsp_context_channel = memory_core_io_reads_1_rsp_payload_context;
  assign b2s_1_rsp_context_channel = _zz_b2s_1_rsp_context_channel[0 : 0];
  assign b2s_1_rsp_context_veryLast = _zz_b2s_1_rsp_context_channel[1];
  assign b2s_1_rsp_context_endPacket = _zz_b2s_1_rsp_context_channel[2];
  assign io_outputs_1_valid = memory_core_io_reads_1_rsp_valid;
  assign io_outputs_1_payload_data = memory_core_io_reads_1_rsp_payload_data;
  assign io_outputs_1_payload_mask = memory_core_io_reads_1_rsp_payload_mask;
  assign io_outputs_1_payload_sink = channels_3_pop_b2s_sinkId;
  assign io_outputs_1_payload_last = (b2s_1_rsp_context_veryLast && b2s_1_rsp_context_endPacket);
  assign io_outputs_1_fire = (io_outputs_1_valid && io_outputs_1_ready);
  assign when_DmaSg_l725_1 = (io_outputs_1_fire && b2s_1_rsp_context_veryLast);
  assign when_DmaSg_l726_1 = b2s_1_rsp_context_channel[0];
  assign _zz_m2b_cmd_s0_priority_masked = channels_1_priority;
  assign _zz_m2b_cmd_s0_priority_masked_1 = channels_3_priority;
  assign _zz_m2b_cmd_s0_priority_masked_2 = (((! channels_3_push_m2b_loadRequest) || (channels_1_push_m2b_loadRequest && (_zz_m2b_cmd_s0_priority_masked_1 < _zz_m2b_cmd_s0_priority_masked))) ? _zz_m2b_cmd_s0_priority_masked : _zz_m2b_cmd_s0_priority_masked_1);
  assign m2b_cmd_s0_priority_masked = {(channels_3_push_m2b_loadRequest && (channels_3_priority == _zz_m2b_cmd_s0_priority_masked_2)),(channels_1_push_m2b_loadRequest && (channels_1_priority == _zz_m2b_cmd_s0_priority_masked_2))};
  assign _zz_m2b_cmd_s0_priority_chosenOh = m2b_cmd_s0_priority_masked;
  assign _zz_m2b_cmd_s0_priority_chosenOh_1 = {_zz_m2b_cmd_s0_priority_chosenOh,_zz_m2b_cmd_s0_priority_chosenOh};
  assign _zz_m2b_cmd_s0_priority_chosenOh_2 = (_zz_m2b_cmd_s0_priority_chosenOh_1 & (~ _zz__zz_m2b_cmd_s0_priority_chosenOh_2));
  assign m2b_cmd_s0_priority_chosenOh = (_zz_m2b_cmd_s0_priority_chosenOh_2[3 : 2] | _zz_m2b_cmd_s0_priority_chosenOh_2[1 : 0]);
  assign _zz_m2b_cmd_s0_priority_chosen = m2b_cmd_s0_priority_chosenOh[1];
  assign m2b_cmd_s0_priority_chosen = _zz_m2b_cmd_s0_priority_chosen;
  assign m2b_cmd_s0_priority_weightLast = _zz_m2b_cmd_s0_priority_weightLast;
  assign m2b_cmd_s0_priority_contextNext = (m2b_cmd_s0_priority_weightLast ? {m2b_cmd_s0_priority_chosenOh[0 : 0],m2b_cmd_s0_priority_chosenOh[1 : 1]} : m2b_cmd_s0_priority_chosenOh);
  assign when_DmaSg_l758 = (! m2b_cmd_s0_valid);
  assign when_DmaSg_l760 = (|{channels_3_push_m2b_loadRequest,channels_1_push_m2b_loadRequest});
  assign when_DmaSg_l763 = (2'b00 == _zz_m2b_cmd_s0_priority_masked_2);
  assign when_DmaSg_l763_1 = (2'b01 == _zz_m2b_cmd_s0_priority_masked_2);
  assign when_DmaSg_l763_2 = (2'b10 == _zz_m2b_cmd_s0_priority_masked_2);
  assign when_DmaSg_l763_3 = (2'b11 == _zz_m2b_cmd_s0_priority_masked_2);
  assign when_DmaSg_l773 = (channels_1_push_m2b_loadRequest && m2b_cmd_s0_priority_chosenOh[0]);
  assign when_DmaSg_l773_1 = (channels_3_push_m2b_loadRequest && m2b_cmd_s0_priority_chosenOh[1]);
  assign m2b_cmd_s0_address = _zz_m2b_cmd_s0_address;
  assign m2b_cmd_s0_bytesLeft = _zz_m2b_cmd_s0_bytesLeft;
  assign m2b_cmd_s0_readAddressBurstRange = m2b_cmd_s0_address[12 : 0];
  assign m2b_cmd_s0_lengthHead = ((~ m2b_cmd_s0_readAddressBurstRange) & _zz_m2b_cmd_s0_lengthHead);
  assign m2b_cmd_s0_length = _zz_m2b_cmd_s0_length[12:0];
  assign m2b_cmd_s0_lastBurst = (m2b_cmd_s0_bytesLeft == _zz_m2b_cmd_s0_lastBurst);
  assign m2b_cmd_s1_context_channel = m2b_cmd_s0_chosen;
  assign m2b_cmd_s1_context_start = m2b_cmd_s1_address[4:0];
  assign m2b_cmd_s1_context_stop = _zz_m2b_cmd_s1_context_stop[4:0];
  assign m2b_cmd_s1_context_last = m2b_cmd_s1_lastBurst;
  assign m2b_cmd_s1_context_length = m2b_cmd_s1_length;
  always @(*) begin
    io_read_cmd_valid = 1'b0;
    if(m2b_cmd_s1_valid) begin
      io_read_cmd_valid = 1'b1;
    end
  end

  assign io_read_cmd_payload_last = 1'b1;
  assign io_read_cmd_payload_fragment_source = m2b_cmd_s0_chosen;
  assign io_read_cmd_payload_fragment_opcode = 1'b0;
  assign io_read_cmd_payload_fragment_address = m2b_cmd_s1_address;
  assign io_read_cmd_payload_fragment_length = m2b_cmd_s1_length;
  assign io_read_cmd_payload_fragment_context = {m2b_cmd_s1_context_last,{m2b_cmd_s1_context_length,{m2b_cmd_s1_context_stop,{m2b_cmd_s1_context_start,m2b_cmd_s1_context_channel}}}};
  assign m2b_cmd_s1_addressNext = (_zz_m2b_cmd_s1_addressNext + 32'h00000001);
  assign m2b_cmd_s1_byteLeftNext = (_zz_m2b_cmd_s1_byteLeftNext - 26'h0000001);
  assign m2b_cmd_s1_fifoPushDecr = (_zz_m2b_cmd_s1_fifoPushDecr >>> 3'd4);
  assign when_DmaSg_l828 = (1'b0 == m2b_cmd_s0_chosen);
  assign when_DmaSg_l828_1 = (1'b1 == m2b_cmd_s0_chosen);
  assign _zz_m2b_rsp_context_channel = io_read_rsp_payload_fragment_context;
  assign m2b_rsp_context_channel = _zz_m2b_rsp_context_channel[0 : 0];
  assign m2b_rsp_context_start = _zz_m2b_rsp_context_channel[5 : 1];
  assign m2b_rsp_context_stop = _zz_m2b_rsp_context_channel[10 : 6];
  assign m2b_rsp_context_length = _zz_m2b_rsp_context_channel[23 : 11];
  assign m2b_rsp_context_last = _zz_m2b_rsp_context_channel[24];
  assign m2b_rsp_veryLast = (m2b_rsp_context_last && io_read_rsp_payload_last);
  assign io_read_rsp_fire = (io_read_rsp_valid && io_read_rsp_ready);
  assign when_DmaSg_l847 = (io_read_rsp_fire && m2b_rsp_veryLast);
  assign when_DmaSg_l848 = (m2b_rsp_context_channel == 1'b0);
  assign when_DmaSg_l848_1 = (m2b_rsp_context_channel == 1'b1);
  always @(*) begin
    memory_core_io_writes_2_cmd_payload_mask[0] = ((! (m2b_rsp_first && (5'h0 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h0))));
    memory_core_io_writes_2_cmd_payload_mask[1] = ((! (m2b_rsp_first && (5'h01 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h01))));
    memory_core_io_writes_2_cmd_payload_mask[2] = ((! (m2b_rsp_first && (5'h02 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h02))));
    memory_core_io_writes_2_cmd_payload_mask[3] = ((! (m2b_rsp_first && (5'h03 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h03))));
    memory_core_io_writes_2_cmd_payload_mask[4] = ((! (m2b_rsp_first && (5'h04 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h04))));
    memory_core_io_writes_2_cmd_payload_mask[5] = ((! (m2b_rsp_first && (5'h05 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h05))));
    memory_core_io_writes_2_cmd_payload_mask[6] = ((! (m2b_rsp_first && (5'h06 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h06))));
    memory_core_io_writes_2_cmd_payload_mask[7] = ((! (m2b_rsp_first && (5'h07 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h07))));
    memory_core_io_writes_2_cmd_payload_mask[8] = ((! (m2b_rsp_first && (5'h08 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h08))));
    memory_core_io_writes_2_cmd_payload_mask[9] = ((! (m2b_rsp_first && (5'h09 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h09))));
    memory_core_io_writes_2_cmd_payload_mask[10] = ((! (m2b_rsp_first && (5'h0a < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h0a))));
    memory_core_io_writes_2_cmd_payload_mask[11] = ((! (m2b_rsp_first && (5'h0b < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h0b))));
    memory_core_io_writes_2_cmd_payload_mask[12] = ((! (m2b_rsp_first && (5'h0c < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h0c))));
    memory_core_io_writes_2_cmd_payload_mask[13] = ((! (m2b_rsp_first && (5'h0d < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h0d))));
    memory_core_io_writes_2_cmd_payload_mask[14] = ((! (m2b_rsp_first && (5'h0e < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h0e))));
    memory_core_io_writes_2_cmd_payload_mask[15] = ((! (m2b_rsp_first && (5'h0f < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h0f))));
    memory_core_io_writes_2_cmd_payload_mask[16] = ((! (m2b_rsp_first && (5'h10 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h10))));
    memory_core_io_writes_2_cmd_payload_mask[17] = ((! (m2b_rsp_first && (5'h11 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h11))));
    memory_core_io_writes_2_cmd_payload_mask[18] = ((! (m2b_rsp_first && (5'h12 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h12))));
    memory_core_io_writes_2_cmd_payload_mask[19] = ((! (m2b_rsp_first && (5'h13 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h13))));
    memory_core_io_writes_2_cmd_payload_mask[20] = ((! (m2b_rsp_first && (5'h14 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h14))));
    memory_core_io_writes_2_cmd_payload_mask[21] = ((! (m2b_rsp_first && (5'h15 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h15))));
    memory_core_io_writes_2_cmd_payload_mask[22] = ((! (m2b_rsp_first && (5'h16 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h16))));
    memory_core_io_writes_2_cmd_payload_mask[23] = ((! (m2b_rsp_first && (5'h17 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h17))));
    memory_core_io_writes_2_cmd_payload_mask[24] = ((! (m2b_rsp_first && (5'h18 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h18))));
    memory_core_io_writes_2_cmd_payload_mask[25] = ((! (m2b_rsp_first && (5'h19 < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h19))));
    memory_core_io_writes_2_cmd_payload_mask[26] = ((! (m2b_rsp_first && (5'h1a < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h1a))));
    memory_core_io_writes_2_cmd_payload_mask[27] = ((! (m2b_rsp_first && (5'h1b < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h1b))));
    memory_core_io_writes_2_cmd_payload_mask[28] = ((! (m2b_rsp_first && (5'h1c < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h1c))));
    memory_core_io_writes_2_cmd_payload_mask[29] = ((! (m2b_rsp_first && (5'h1d < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h1d))));
    memory_core_io_writes_2_cmd_payload_mask[30] = ((! (m2b_rsp_first && (5'h1e < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h1e))));
    memory_core_io_writes_2_cmd_payload_mask[31] = ((! (m2b_rsp_first && (5'h1f < m2b_rsp_context_start))) && (! (io_read_rsp_payload_last && (m2b_rsp_context_stop < 5'h1f))));
  end

  assign m2b_rsp_writeContext_last = m2b_rsp_veryLast;
  assign m2b_rsp_writeContext_lastOfBurst = io_read_rsp_payload_last;
  assign m2b_rsp_writeContext_channel = m2b_rsp_context_channel;
  assign m2b_rsp_writeContext_loadByteInNextBeat = ({1'b0,(io_read_rsp_payload_last ? m2b_rsp_context_stop : 5'h1f)} - {1'b0,(m2b_rsp_first ? m2b_rsp_context_start : 5'h0)});
  assign memory_core_io_writes_2_cmd_payload_address = _zz_io_writes_2_cmd_payload_address[12:0];
  assign io_read_rsp_ready = memory_core_io_writes_2_cmd_ready;
  assign memory_core_io_writes_2_cmd_payload_context = {m2b_rsp_writeContext_loadByteInNextBeat,{m2b_rsp_writeContext_channel,{m2b_rsp_writeContext_lastOfBurst,m2b_rsp_writeContext_last}}};
  assign memory_core_io_writes_2_cmd_fire = (io_read_rsp_valid && memory_core_io_writes_2_cmd_ready);
  assign _zz_m2b_writeRsp_context_last = memory_core_io_writes_2_rsp_payload_context;
  assign m2b_writeRsp_context_last = _zz_m2b_writeRsp_context_last[0];
  assign m2b_writeRsp_context_lastOfBurst = _zz_m2b_writeRsp_context_last[1];
  assign m2b_writeRsp_context_channel = _zz_m2b_writeRsp_context_last[2 : 2];
  assign m2b_writeRsp_context_loadByteInNextBeat = _zz_m2b_writeRsp_context_last[8 : 3];
  assign _zz_channels_1_fifo_pop_bytesIncr_value = (memory_core_io_writes_2_rsp_valid && (m2b_writeRsp_context_channel == 1'b0));
  assign when_DmaSg_l893 = (_zz_channels_1_fifo_pop_bytesIncr_value && m2b_writeRsp_context_lastOfBurst);
  assign _zz_channels_3_fifo_pop_bytesIncr_value = (memory_core_io_writes_2_rsp_valid && (m2b_writeRsp_context_channel == 1'b1));
  assign when_DmaSg_l893_1 = (_zz_channels_3_fifo_pop_bytesIncr_value && m2b_writeRsp_context_lastOfBurst);
  assign _zz_b2m_fsm_arbiter_logic_priority_masked = channels_0_priority;
  assign _zz_b2m_fsm_arbiter_logic_priority_masked_1 = channels_2_priority;
  assign _zz_b2m_fsm_arbiter_logic_priority_masked_2 = (((! channels_2_pop_b2m_request) || (channels_0_pop_b2m_request && (_zz_b2m_fsm_arbiter_logic_priority_masked_1 < _zz_b2m_fsm_arbiter_logic_priority_masked))) ? _zz_b2m_fsm_arbiter_logic_priority_masked : _zz_b2m_fsm_arbiter_logic_priority_masked_1);
  assign b2m_fsm_arbiter_logic_priority_masked = {(channels_2_pop_b2m_request && (channels_2_priority == _zz_b2m_fsm_arbiter_logic_priority_masked_2)),(channels_0_pop_b2m_request && (channels_0_priority == _zz_b2m_fsm_arbiter_logic_priority_masked_2))};
  assign _zz_b2m_fsm_arbiter_logic_priority_chosenOh = b2m_fsm_arbiter_logic_priority_masked;
  assign _zz_b2m_fsm_arbiter_logic_priority_chosenOh_1 = {_zz_b2m_fsm_arbiter_logic_priority_chosenOh,_zz_b2m_fsm_arbiter_logic_priority_chosenOh};
  assign _zz_b2m_fsm_arbiter_logic_priority_chosenOh_2 = (_zz_b2m_fsm_arbiter_logic_priority_chosenOh_1 & (~ _zz__zz_b2m_fsm_arbiter_logic_priority_chosenOh_2));
  assign b2m_fsm_arbiter_logic_priority_chosenOh = (_zz_b2m_fsm_arbiter_logic_priority_chosenOh_2[3 : 2] | _zz_b2m_fsm_arbiter_logic_priority_chosenOh_2[1 : 0]);
  assign _zz_b2m_fsm_arbiter_logic_priority_chosen = b2m_fsm_arbiter_logic_priority_chosenOh[1];
  assign b2m_fsm_arbiter_logic_priority_chosen = _zz_b2m_fsm_arbiter_logic_priority_chosen;
  assign b2m_fsm_arbiter_logic_priority_weightLast = _zz_b2m_fsm_arbiter_logic_priority_weightLast;
  assign b2m_fsm_arbiter_logic_priority_contextNext = (b2m_fsm_arbiter_logic_priority_weightLast ? {b2m_fsm_arbiter_logic_priority_chosenOh[0 : 0],b2m_fsm_arbiter_logic_priority_chosenOh[1 : 1]} : b2m_fsm_arbiter_logic_priority_chosenOh);
  assign when_DmaSg_l758_1 = (! b2m_fsm_arbiter_logic_valid);
  assign when_DmaSg_l760_1 = (|{channels_2_pop_b2m_request,channels_0_pop_b2m_request});
  assign when_DmaSg_l763_4 = (2'b00 == _zz_b2m_fsm_arbiter_logic_priority_masked_2);
  assign when_DmaSg_l763_5 = (2'b01 == _zz_b2m_fsm_arbiter_logic_priority_masked_2);
  assign when_DmaSg_l763_6 = (2'b10 == _zz_b2m_fsm_arbiter_logic_priority_masked_2);
  assign when_DmaSg_l763_7 = (2'b11 == _zz_b2m_fsm_arbiter_logic_priority_masked_2);
  assign when_DmaSg_l773_2 = (channels_0_pop_b2m_request && b2m_fsm_arbiter_logic_priority_chosenOh[0]);
  assign when_DmaSg_l773_3 = (channels_2_pop_b2m_request && b2m_fsm_arbiter_logic_priority_chosenOh[1]);
  assign when_DmaSg_l935 = ((! b2m_fsm_sel_valid) && b2m_fsm_arbiter_logic_valid);
  assign _zz_1 = ({1'd0,1'b1} <<< b2m_fsm_arbiter_logic_chosen);
  assign b2m_fsm_bytesInBurstP1 = ({1'b0,b2m_fsm_sel_bytesInBurst} + _zz_b2m_fsm_bytesInBurstP1);
  assign b2m_fsm_addressNext = (b2m_fsm_sel_address + _zz_b2m_fsm_addressNext);
  assign b2m_fsm_bytesLeftNext = ({1'b0,b2m_fsm_sel_bytesLeft} - _zz_b2m_fsm_bytesLeftNext);
  assign b2m_fsm_isFinalCmd = b2m_fsm_bytesLeftNext[26];
  assign b2m_fsm_s0 = (b2m_fsm_sel_valid && (! b2m_fsm_sel_valid_regNext));
  assign when_DmaSg_l986 = (! b2m_fsm_sel_valid);
  assign _zz_b2m_fsm_sel_bytesInBurst = (b2m_fsm_sel_bytesInFifo - 18'h00001);
  assign _zz_b2m_fsm_sel_bytesInBurst_1 = ((_zz__zz_b2m_fsm_sel_bytesInBurst_1 < b2m_fsm_sel_bytesLeft) ? _zz__zz_b2m_fsm_sel_bytesInBurst_1_1 : b2m_fsm_sel_bytesLeft);
  assign _zz_b2m_fsm_sel_bytesInBurst_2 = (b2m_fsm_sel_bytePerBurst - (_zz__zz_b2m_fsm_sel_bytesInBurst_2 & b2m_fsm_sel_bytePerBurst));
  assign b2m_fsm_fifoCompletion = (_zz_b2m_fsm_fifoCompletion == _zz_b2m_fsm_fifoCompletion_1);
  assign when_DmaSg_l996 = (b2m_fsm_sel_channel == 1'b0);
  assign when_DmaSg_l1001 = (! b2m_fsm_fifoCompletion);
  assign when_DmaSg_l996_1 = (b2m_fsm_sel_channel == 1'b1);
  assign when_DmaSg_l1001_1 = (! b2m_fsm_fifoCompletion);
  assign when_DmaSg_l1013 = (b2m_fsm_sel_valid && b2m_fsm_sel_ready);
  always @(*) begin
    b2m_fsm_sel_ready = 1'b0;
    if(when_DmaSg_l1102) begin
      b2m_fsm_sel_ready = 1'b1;
    end
  end

  assign b2m_fsm_fetch_context_ptr = _zz_b2m_fsm_fetch_context_ptr;
  assign b2m_fsm_fetch_context_toggle = b2m_fsm_toggle;
  assign memory_core_io_reads_2_cmd_payload_address = b2m_fsm_sel_ptr[12:0];
  assign memory_core_io_reads_2_cmd_payload_context = {b2m_fsm_fetch_context_toggle,b2m_fsm_fetch_context_ptr};
  assign when_DmaSg_l1033 = (b2m_fsm_sel_valid && memory_core_io_reads_2_cmd_ready);
  assign _zz_b2m_fsm_aggregate_context_ptr = memory_core_io_reads_2_rsp_payload_context;
  assign b2m_fsm_aggregate_context_ptr = _zz_b2m_fsm_aggregate_context_ptr[13 : 0];
  assign b2m_fsm_aggregate_context_toggle = _zz_b2m_fsm_aggregate_context_ptr[14];
  assign memory_core_io_reads_2_rsp_s2mPipe_valid = (memory_core_io_reads_2_rsp_valid || (! memory_core_io_reads_2_rsp_rValidN));
  assign memory_core_io_reads_2_rsp_s2mPipe_payload_data = (memory_core_io_reads_2_rsp_rValidN ? memory_core_io_reads_2_rsp_payload_data : memory_core_io_reads_2_rsp_rData_data);
  assign memory_core_io_reads_2_rsp_s2mPipe_payload_mask = (memory_core_io_reads_2_rsp_rValidN ? memory_core_io_reads_2_rsp_payload_mask : memory_core_io_reads_2_rsp_rData_mask);
  assign memory_core_io_reads_2_rsp_s2mPipe_payload_context = (memory_core_io_reads_2_rsp_rValidN ? memory_core_io_reads_2_rsp_payload_context : memory_core_io_reads_2_rsp_rData_context);
  assign when_Stream_l445 = (b2m_fsm_aggregate_context_toggle != b2m_fsm_toggle);
  always @(*) begin
    b2m_fsm_aggregate_memoryPort_valid = memory_core_io_reads_2_rsp_s2mPipe_valid;
    if(when_Stream_l445) begin
      b2m_fsm_aggregate_memoryPort_valid = 1'b0;
    end
  end

  always @(*) begin
    memory_core_io_reads_2_rsp_s2mPipe_ready = b2m_fsm_aggregate_memoryPort_ready;
    if(when_Stream_l445) begin
      memory_core_io_reads_2_rsp_s2mPipe_ready = 1'b1;
    end
  end

  assign b2m_fsm_aggregate_memoryPort_payload_data = memory_core_io_reads_2_rsp_s2mPipe_payload_data;
  assign b2m_fsm_aggregate_memoryPort_payload_mask = memory_core_io_reads_2_rsp_s2mPipe_payload_mask;
  assign b2m_fsm_aggregate_memoryPort_payload_context = memory_core_io_reads_2_rsp_s2mPipe_payload_context;
  assign b2m_fsm_aggregate_memoryPort_fire = (b2m_fsm_aggregate_memoryPort_valid && b2m_fsm_aggregate_memoryPort_ready);
  assign when_DmaSg_l1050 = (! (b2m_fsm_sel_valid && (! b2m_fsm_sel_ready)));
  assign b2m_fsm_aggregate_bytesToSkip = _zz_b2m_fsm_aggregate_bytesToSkip;
  assign b2m_fsm_aggregate_bytesToSkipMask = {((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h1f)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= 5'h1e)),{((! b2m_fsm_aggregate_first) || (b2m_fsm_aggregate_bytesToSkip <= _zz_b2m_fsm_aggregate_bytesToSkipMask)),{(_zz_b2m_fsm_aggregate_bytesToSkipMask_1 || _zz_b2m_fsm_aggregate_bytesToSkipMask_2),{_zz_b2m_fsm_aggregate_bytesToSkipMask_3,{_zz_b2m_fsm_aggregate_bytesToSkipMask_4,_zz_b2m_fsm_aggregate_bytesToSkipMask_5}}}}}};
  assign b2m_fsm_aggregate_memoryPort_ready = b2m_fsm_aggregate_engine_io_input_ready;
  assign b2m_fsm_aggregate_engine_io_input_payload_mask = (b2m_fsm_aggregate_memoryPort_payload_mask & b2m_fsm_aggregate_bytesToSkipMask);
  assign b2m_fsm_aggregate_engine_io_offset = b2m_fsm_sel_address[4:0];
  assign b2m_fsm_aggregate_engine_io_flush = (! _zz_io_flush);
  assign b2m_fsm_cmd_maskFirstTrigger = b2m_fsm_sel_address[4:0];
  assign b2m_fsm_cmd_maskLastTriggerComb = (b2m_fsm_cmd_maskFirstTrigger + _zz_b2m_fsm_cmd_maskLastTriggerComb);
  assign b2m_fsm_cmd_maskFirst = {(b2m_fsm_cmd_maskFirstTrigger <= 5'h1f),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h1e),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h1d),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h1c),{(b2m_fsm_cmd_maskFirstTrigger <= 5'h1b),{(b2m_fsm_cmd_maskFirstTrigger <= _zz_b2m_fsm_cmd_maskFirst),{_zz_b2m_fsm_cmd_maskFirst_1,{_zz_b2m_fsm_cmd_maskFirst_2,_zz_b2m_fsm_cmd_maskFirst_3}}}}}}}};
  assign b2m_fsm_cmd_enoughAggregation = (((b2m_fsm_s2 && b2m_fsm_sel_valid) && (! b2m_fsm_aggregate_engine_io_flush)) && (io_write_cmd_payload_last ? ((b2m_fsm_aggregate_engine_io_output_mask & b2m_fsm_cmd_maskLast) == b2m_fsm_cmd_maskLast) : (&b2m_fsm_aggregate_engine_io_output_mask)));
  assign io_write_cmd_fire = (io_write_cmd_valid && io_write_cmd_ready);
  assign io_write_cmd_valid = b2m_fsm_cmd_enoughAggregation;
  assign io_write_cmd_payload_last = (b2m_fsm_beatCounter == 8'h0);
  assign io_write_cmd_payload_fragment_address = b2m_fsm_sel_address;
  assign io_write_cmd_payload_fragment_opcode = 1'b1;
  assign io_write_cmd_payload_fragment_data = b2m_fsm_aggregate_engine_io_output_data;
  assign io_write_cmd_payload_fragment_mask = (~ ((io_write_cmd_payload_first ? (~ b2m_fsm_cmd_maskFirst) : 32'h0) | (io_write_cmd_payload_last ? (~ b2m_fsm_cmd_maskLast) : 32'h0)));
  assign io_write_cmd_payload_fragment_length = b2m_fsm_sel_bytesInBurst;
  assign io_write_cmd_payload_fragment_source = b2m_fsm_sel_channel;
  assign b2m_fsm_cmd_doPtrIncr = (b2m_fsm_sel_valid && (b2m_fsm_aggregate_engine_io_output_consumed || ((io_write_cmd_fire && io_write_cmd_payload_last) && (b2m_fsm_aggregate_engine_io_output_usedUntil == 5'h1f))));
  assign b2m_fsm_cmd_context_channel = b2m_fsm_sel_channel;
  assign b2m_fsm_cmd_context_length = b2m_fsm_sel_bytesInBurst;
  assign b2m_fsm_cmd_context_doPacketSync = (b2m_fsm_sel_packet && b2m_fsm_fifoCompletion);
  assign io_write_cmd_payload_fragment_context = {b2m_fsm_cmd_context_doPacketSync,{b2m_fsm_cmd_context_length,b2m_fsm_cmd_context_channel}};
  assign when_DmaSg_l1102 = (io_write_cmd_fire && io_write_cmd_payload_last);
  assign _zz_2 = ({1'd0,1'b1} <<< b2m_fsm_sel_channel);
  assign _zz_channels_0_pop_b2m_bytesToSkip = (b2m_fsm_aggregate_engine_io_output_usedUntil + 5'h01);
  assign io_write_rsp_ready = 1'b1;
  assign _zz_b2m_rsp_context_channel = io_write_rsp_payload_fragment_context;
  assign b2m_rsp_context_channel = _zz_b2m_rsp_context_channel[0 : 0];
  assign b2m_rsp_context_length = _zz_b2m_rsp_context_channel[13 : 1];
  assign b2m_rsp_context_doPacketSync = _zz_b2m_rsp_context_channel[14];
  assign io_write_rsp_fire = (io_write_rsp_valid && io_write_rsp_ready);
  assign _zz_3 = ({1'd0,1'b1} <<< b2m_rsp_context_channel);
  assign when_DmaSg_l1116 = (b2m_rsp_context_channel == 1'b0);
  assign when_DmaSg_l1116_1 = (b2m_rsp_context_channel == 1'b1);
  always @(*) begin
    io_interrupts = 4'b0000;
    if(channels_0_interrupts_completion_valid) begin
      io_interrupts[0] = 1'b1;
    end
    if(channels_0_interrupts_onChannelCompletion_valid) begin
      io_interrupts[0] = 1'b1;
    end
    if(channels_0_interrupts_s2mPacket_valid) begin
      io_interrupts[0] = 1'b1;
    end
    if(channels_1_interrupts_completion_valid) begin
      io_interrupts[1] = 1'b1;
    end
    if(channels_1_interrupts_onChannelCompletion_valid) begin
      io_interrupts[1] = 1'b1;
    end
    if(channels_2_interrupts_completion_valid) begin
      io_interrupts[2] = 1'b1;
    end
    if(channels_2_interrupts_onChannelCompletion_valid) begin
      io_interrupts[2] = 1'b1;
    end
    if(channels_2_interrupts_s2mPacket_valid) begin
      io_interrupts[2] = 1'b1;
    end
    if(channels_3_interrupts_completion_valid) begin
      io_interrupts[3] = 1'b1;
    end
    if(channels_3_interrupts_onChannelCompletion_valid) begin
      io_interrupts[3] = 1'b1;
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377 = 1'b0;
    case(io_ctrl_PADDR)
      14'h002c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l377_1 = 1'b0;
    case(io_ctrl_PADDR)
      14'h002c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_1 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341 = 1'b0;
    case(io_ctrl_PADDR)
      14'h0054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341_1 = 1'b0;
    case(io_ctrl_PADDR)
      14'h0054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_1 = io_ctrl_PWDATA[2];
  always @(*) begin
    when_BusSlaveFactory_l341_2 = 1'b0;
    case(io_ctrl_PADDR)
      14'h0054 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_2 = io_ctrl_PWDATA[4];
  always @(*) begin
    when_BusSlaveFactory_l377_2 = 1'b0;
    case(io_ctrl_PADDR)
      14'h00ac : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_2 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l377_3 = 1'b0;
    case(io_ctrl_PADDR)
      14'h00ac : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_3 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341_3 = 1'b0;
    case(io_ctrl_PADDR)
      14'h00d4 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_3 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341_4 = 1'b0;
    case(io_ctrl_PADDR)
      14'h00d4 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_4 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_4 = io_ctrl_PWDATA[2];
  always @(*) begin
    when_BusSlaveFactory_l377_4 = 1'b0;
    case(io_ctrl_PADDR)
      14'h012c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_4 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_4 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l377_5 = 1'b0;
    case(io_ctrl_PADDR)
      14'h012c : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_5 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_5 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341_5 = 1'b0;
    case(io_ctrl_PADDR)
      14'h0154 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_5 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_5 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341_6 = 1'b0;
    case(io_ctrl_PADDR)
      14'h0154 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_6 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_6 = io_ctrl_PWDATA[2];
  always @(*) begin
    when_BusSlaveFactory_l341_7 = 1'b0;
    case(io_ctrl_PADDR)
      14'h0154 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_7 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_7 = io_ctrl_PWDATA[4];
  always @(*) begin
    when_BusSlaveFactory_l377_6 = 1'b0;
    case(io_ctrl_PADDR)
      14'h01ac : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_6 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_6 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l377_7 = 1'b0;
    case(io_ctrl_PADDR)
      14'h01ac : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l377_7 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_7 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341_8 = 1'b0;
    case(io_ctrl_PADDR)
      14'h01d4 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_8 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_8 = io_ctrl_PWDATA[0];
  always @(*) begin
    when_BusSlaveFactory_l341_9 = 1'b0;
    case(io_ctrl_PADDR)
      14'h01d4 : begin
        if(ctrl_doWrite) begin
          when_BusSlaveFactory_l341_9 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_9 = io_ctrl_PWDATA[2];
  assign when_Apb3SlaveFactory_l81 = ((io_ctrl_PADDR & (~ 14'h0003)) == 14'h0010);
  assign when_Apb3SlaveFactory_l81_1 = ((io_ctrl_PADDR & (~ 14'h0003)) == 14'h0080);
  assign when_Apb3SlaveFactory_l81_2 = ((io_ctrl_PADDR & (~ 14'h0003)) == 14'h0110);
  assign when_Apb3SlaveFactory_l81_3 = ((io_ctrl_PADDR & (~ 14'h0003)) == 14'h0180);
  assign channels_0_fifo_push_ptrIncr_value = _zz_channels_0_fifo_push_ptrIncr_value;
  assign channels_0_fifo_pop_bytesIncr_value = _zz_channels_0_fifo_pop_bytesIncr_value_1;
  assign channels_0_fifo_pop_bytesDecr_value = channels_0_pop_b2m_decrBytes;
  assign channels_0_fifo_pop_ptrIncr_value = _zz_channels_0_fifo_pop_ptrIncr_value;
  assign channels_1_fifo_push_ptrIncr_value = _zz_channels_1_fifo_push_ptrIncr_value;
  assign channels_1_fifo_pop_bytesIncr_value = _zz_channels_1_fifo_pop_bytesIncr_value_1;
  assign channels_1_fifo_pop_bytesDecr_value = 18'h0;
  assign channels_1_fifo_pop_ptrIncr_value = _zz_channels_1_fifo_pop_ptrIncr_value;
  assign channels_2_fifo_push_ptrIncr_value = _zz_channels_2_fifo_push_ptrIncr_value;
  assign channels_2_fifo_pop_bytesIncr_value = _zz_channels_2_fifo_pop_bytesIncr_value_1;
  assign channels_2_fifo_pop_bytesDecr_value = channels_2_pop_b2m_decrBytes;
  assign channels_2_fifo_pop_ptrIncr_value = _zz_channels_2_fifo_pop_ptrIncr_value;
  assign channels_3_fifo_push_ptrIncr_value = _zz_channels_3_fifo_push_ptrIncr_value;
  assign channels_3_fifo_pop_bytesIncr_value = _zz_channels_3_fifo_pop_bytesIncr_value_1;
  assign channels_3_fifo_pop_bytesDecr_value = 18'h0;
  assign channels_3_fifo_pop_ptrIncr_value = _zz_channels_3_fifo_pop_ptrIncr_value;
  always @(posedge clk) begin
    if(reset) begin
      channels_0_channelValid <= 1'b0;
      channels_0_descriptorValid <= 1'b0;
      channels_0_priority <= 2'b00;
      channels_0_weight <= 2'b00;
      channels_0_ctrl_kick <= 1'b0;
      channels_0_pop_b2m_memPending <= 4'b0000;
      channels_0_interrupts_completion_enable <= 1'b0;
      channels_0_interrupts_completion_valid <= 1'b0;
      channels_0_interrupts_onChannelCompletion_enable <= 1'b0;
      channels_0_interrupts_onChannelCompletion_valid <= 1'b0;
      channels_0_interrupts_s2mPacket_enable <= 1'b0;
      channels_0_interrupts_s2mPacket_valid <= 1'b0;
      channels_1_channelValid <= 1'b0;
      channels_1_descriptorValid <= 1'b0;
      channels_1_priority <= 2'b00;
      channels_1_weight <= 2'b00;
      channels_1_ctrl_kick <= 1'b0;
      channels_1_push_m2b_loadDone <= 1'b1;
      channels_1_push_m2b_memPending <= 4'b0000;
      channels_1_interrupts_completion_enable <= 1'b0;
      channels_1_interrupts_completion_valid <= 1'b0;
      channels_1_interrupts_onChannelCompletion_enable <= 1'b0;
      channels_1_interrupts_onChannelCompletion_valid <= 1'b0;
      channels_2_channelValid <= 1'b0;
      channels_2_descriptorValid <= 1'b0;
      channels_2_priority <= 2'b00;
      channels_2_weight <= 2'b00;
      channels_2_ctrl_kick <= 1'b0;
      channels_2_pop_b2m_memPending <= 4'b0000;
      channels_2_interrupts_completion_enable <= 1'b0;
      channels_2_interrupts_completion_valid <= 1'b0;
      channels_2_interrupts_onChannelCompletion_enable <= 1'b0;
      channels_2_interrupts_onChannelCompletion_valid <= 1'b0;
      channels_2_interrupts_s2mPacket_enable <= 1'b0;
      channels_2_interrupts_s2mPacket_valid <= 1'b0;
      channels_3_channelValid <= 1'b0;
      channels_3_descriptorValid <= 1'b0;
      channels_3_priority <= 2'b00;
      channels_3_weight <= 2'b00;
      channels_3_ctrl_kick <= 1'b0;
      channels_3_push_m2b_loadDone <= 1'b1;
      channels_3_push_m2b_memPending <= 4'b0000;
      channels_3_interrupts_completion_enable <= 1'b0;
      channels_3_interrupts_completion_valid <= 1'b0;
      channels_3_interrupts_onChannelCompletion_enable <= 1'b0;
      channels_3_interrupts_onChannelCompletion_valid <= 1'b0;
      io_inputs_0_payload_last_regNextWhen <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_1 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_2 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_3 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_4 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_5 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_6 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_7 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_8 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_9 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_10 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_11 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_12 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_13 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_14 <= 1'b1;
      io_inputs_0_payload_last_regNextWhen_15 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_1 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_2 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_3 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_4 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_5 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_6 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_7 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_8 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_9 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_10 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_11 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_12 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_13 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_14 <= 1'b1;
      io_inputs_1_payload_last_regNextWhen_15 <= 1'b1;
      m2b_cmd_s0_valid <= 1'b0;
      m2b_cmd_s0_priority_roundRobins_0 <= 2'b01;
      m2b_cmd_s0_priority_roundRobins_1 <= 2'b01;
      m2b_cmd_s0_priority_roundRobins_2 <= 2'b01;
      m2b_cmd_s0_priority_roundRobins_3 <= 2'b01;
      m2b_cmd_s0_priority_counter <= 2'b00;
      m2b_cmd_s1_valid <= 1'b0;
      m2b_rsp_first <= 1'b1;
      b2m_fsm_sel_valid <= 1'b0;
      b2m_fsm_arbiter_logic_valid <= 1'b0;
      b2m_fsm_arbiter_logic_priority_roundRobins_0 <= 2'b01;
      b2m_fsm_arbiter_logic_priority_roundRobins_1 <= 2'b01;
      b2m_fsm_arbiter_logic_priority_roundRobins_2 <= 2'b01;
      b2m_fsm_arbiter_logic_priority_roundRobins_3 <= 2'b01;
      b2m_fsm_arbiter_logic_priority_counter <= 2'b00;
      b2m_fsm_sel_valid_regNext <= 1'b0;
      b2m_fsm_s1 <= 1'b0;
      b2m_fsm_s2 <= 1'b0;
      b2m_fsm_toggle <= 1'b0;
      memory_core_io_reads_2_rsp_rValidN <= 1'b1;
      _zz_io_flush <= 1'b0;
      io_write_cmd_payload_first <= 1'b1;
    end else begin
      if(channels_0_channelStart) begin
        channels_0_channelValid <= 1'b1;
      end
      if(channels_0_channelCompletion) begin
        channels_0_channelValid <= 1'b0;
      end
      if(channels_0_descriptorStart) begin
        channels_0_descriptorValid <= 1'b1;
      end
      if(channels_0_descriptorCompletion) begin
        channels_0_descriptorValid <= 1'b0;
      end
      channels_0_ctrl_kick <= 1'b0;
      if(channels_0_channelCompletion) begin
        channels_0_ctrl_kick <= 1'b0;
      end
      channels_0_pop_b2m_memPending <= (_zz_channels_0_pop_b2m_memPending - _zz_channels_0_pop_b2m_memPending_3);
      if(when_DmaSg_l255) begin
        channels_0_interrupts_completion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_1) begin
        channels_0_interrupts_completion_valid <= 1'b0;
      end
      if(when_DmaSg_l255_2) begin
        channels_0_interrupts_onChannelCompletion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_3) begin
        channels_0_interrupts_onChannelCompletion_valid <= 1'b0;
      end
      if(channels_0_pop_b2m_packetSync) begin
        channels_0_interrupts_s2mPacket_valid <= 1'b1;
      end
      if(when_DmaSg_l255_4) begin
        channels_0_interrupts_s2mPacket_valid <= 1'b0;
      end
      if(channels_1_channelStart) begin
        channels_1_channelValid <= 1'b1;
      end
      if(channels_1_channelCompletion) begin
        channels_1_channelValid <= 1'b0;
      end
      if(channels_1_descriptorStart) begin
        channels_1_descriptorValid <= 1'b1;
      end
      if(channels_1_descriptorCompletion) begin
        channels_1_descriptorValid <= 1'b0;
      end
      channels_1_ctrl_kick <= 1'b0;
      if(channels_1_channelCompletion) begin
        channels_1_ctrl_kick <= 1'b0;
      end
      channels_1_push_m2b_memPending <= (_zz_channels_1_push_m2b_memPending - _zz_channels_1_push_m2b_memPending_3);
      if(channels_1_descriptorStart) begin
        channels_1_push_m2b_loadDone <= 1'b0;
      end
      if(when_DmaSg_l255_5) begin
        channels_1_interrupts_completion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_6) begin
        channels_1_interrupts_completion_valid <= 1'b0;
      end
      if(when_DmaSg_l255_7) begin
        channels_1_interrupts_onChannelCompletion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_8) begin
        channels_1_interrupts_onChannelCompletion_valid <= 1'b0;
      end
      if(channels_2_channelStart) begin
        channels_2_channelValid <= 1'b1;
      end
      if(channels_2_channelCompletion) begin
        channels_2_channelValid <= 1'b0;
      end
      if(channels_2_descriptorStart) begin
        channels_2_descriptorValid <= 1'b1;
      end
      if(channels_2_descriptorCompletion) begin
        channels_2_descriptorValid <= 1'b0;
      end
      channels_2_ctrl_kick <= 1'b0;
      if(channels_2_channelCompletion) begin
        channels_2_ctrl_kick <= 1'b0;
      end
      channels_2_pop_b2m_memPending <= (_zz_channels_2_pop_b2m_memPending - _zz_channels_2_pop_b2m_memPending_3);
      if(when_DmaSg_l255_9) begin
        channels_2_interrupts_completion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_10) begin
        channels_2_interrupts_completion_valid <= 1'b0;
      end
      if(when_DmaSg_l255_11) begin
        channels_2_interrupts_onChannelCompletion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_12) begin
        channels_2_interrupts_onChannelCompletion_valid <= 1'b0;
      end
      if(channels_2_pop_b2m_packetSync) begin
        channels_2_interrupts_s2mPacket_valid <= 1'b1;
      end
      if(when_DmaSg_l255_13) begin
        channels_2_interrupts_s2mPacket_valid <= 1'b0;
      end
      if(channels_3_channelStart) begin
        channels_3_channelValid <= 1'b1;
      end
      if(channels_3_channelCompletion) begin
        channels_3_channelValid <= 1'b0;
      end
      if(channels_3_descriptorStart) begin
        channels_3_descriptorValid <= 1'b1;
      end
      if(channels_3_descriptorCompletion) begin
        channels_3_descriptorValid <= 1'b0;
      end
      channels_3_ctrl_kick <= 1'b0;
      if(channels_3_channelCompletion) begin
        channels_3_ctrl_kick <= 1'b0;
      end
      channels_3_push_m2b_memPending <= (_zz_channels_3_push_m2b_memPending - _zz_channels_3_push_m2b_memPending_3);
      if(channels_3_descriptorStart) begin
        channels_3_push_m2b_loadDone <= 1'b0;
      end
      if(when_DmaSg_l255_14) begin
        channels_3_interrupts_completion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_15) begin
        channels_3_interrupts_completion_valid <= 1'b0;
      end
      if(when_DmaSg_l255_16) begin
        channels_3_interrupts_onChannelCompletion_valid <= 1'b1;
      end
      if(when_DmaSg_l255_17) begin
        channels_3_interrupts_onChannelCompletion_valid <= 1'b0;
      end
      if(when_package_l12) begin
        io_inputs_0_payload_last_regNextWhen <= io_inputs_0_payload_last;
      end
      if(when_package_l12_1) begin
        io_inputs_0_payload_last_regNextWhen_1 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_2) begin
        io_inputs_0_payload_last_regNextWhen_2 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_3) begin
        io_inputs_0_payload_last_regNextWhen_3 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_4) begin
        io_inputs_0_payload_last_regNextWhen_4 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_5) begin
        io_inputs_0_payload_last_regNextWhen_5 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_6) begin
        io_inputs_0_payload_last_regNextWhen_6 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_7) begin
        io_inputs_0_payload_last_regNextWhen_7 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_8) begin
        io_inputs_0_payload_last_regNextWhen_8 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_9) begin
        io_inputs_0_payload_last_regNextWhen_9 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_10) begin
        io_inputs_0_payload_last_regNextWhen_10 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_11) begin
        io_inputs_0_payload_last_regNextWhen_11 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_12) begin
        io_inputs_0_payload_last_regNextWhen_12 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_13) begin
        io_inputs_0_payload_last_regNextWhen_13 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_14) begin
        io_inputs_0_payload_last_regNextWhen_14 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_15) begin
        io_inputs_0_payload_last_regNextWhen_15 <= io_inputs_0_payload_last;
      end
      if(when_package_l12_16) begin
        io_inputs_1_payload_last_regNextWhen <= io_inputs_1_payload_last;
      end
      if(when_package_l12_17) begin
        io_inputs_1_payload_last_regNextWhen_1 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_18) begin
        io_inputs_1_payload_last_regNextWhen_2 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_19) begin
        io_inputs_1_payload_last_regNextWhen_3 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_20) begin
        io_inputs_1_payload_last_regNextWhen_4 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_21) begin
        io_inputs_1_payload_last_regNextWhen_5 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_22) begin
        io_inputs_1_payload_last_regNextWhen_6 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_23) begin
        io_inputs_1_payload_last_regNextWhen_7 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_24) begin
        io_inputs_1_payload_last_regNextWhen_8 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_25) begin
        io_inputs_1_payload_last_regNextWhen_9 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_26) begin
        io_inputs_1_payload_last_regNextWhen_10 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_27) begin
        io_inputs_1_payload_last_regNextWhen_11 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_28) begin
        io_inputs_1_payload_last_regNextWhen_12 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_29) begin
        io_inputs_1_payload_last_regNextWhen_13 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_30) begin
        io_inputs_1_payload_last_regNextWhen_14 <= io_inputs_1_payload_last;
      end
      if(when_package_l12_31) begin
        io_inputs_1_payload_last_regNextWhen_15 <= io_inputs_1_payload_last;
      end
      if(when_DmaSg_l758) begin
        if(when_DmaSg_l760) begin
          m2b_cmd_s0_valid <= 1'b1;
          if(when_DmaSg_l763) begin
            m2b_cmd_s0_priority_roundRobins_0 <= m2b_cmd_s0_priority_contextNext;
          end
          if(when_DmaSg_l763_1) begin
            m2b_cmd_s0_priority_roundRobins_1 <= m2b_cmd_s0_priority_contextNext;
          end
          if(when_DmaSg_l763_2) begin
            m2b_cmd_s0_priority_roundRobins_2 <= m2b_cmd_s0_priority_contextNext;
          end
          if(when_DmaSg_l763_3) begin
            m2b_cmd_s0_priority_roundRobins_3 <= m2b_cmd_s0_priority_contextNext;
          end
          m2b_cmd_s0_priority_counter <= (m2b_cmd_s0_priority_counter + 2'b01);
          if(m2b_cmd_s0_priority_weightLast) begin
            m2b_cmd_s0_priority_counter <= 2'b00;
          end
        end
      end
      if(m2b_cmd_s0_valid) begin
        m2b_cmd_s1_valid <= 1'b1;
      end
      if(m2b_cmd_s1_valid) begin
        if(io_read_cmd_ready) begin
          m2b_cmd_s0_valid <= 1'b0;
          m2b_cmd_s1_valid <= 1'b0;
          if(when_DmaSg_l828) begin
            if(m2b_cmd_s1_lastBurst) begin
              channels_1_push_m2b_loadDone <= 1'b1;
            end
          end
          if(when_DmaSg_l828_1) begin
            if(m2b_cmd_s1_lastBurst) begin
              channels_3_push_m2b_loadDone <= 1'b1;
            end
          end
        end
      end
      if(io_read_rsp_fire) begin
        m2b_rsp_first <= io_read_rsp_payload_last;
      end
      if(when_DmaSg_l758_1) begin
        if(when_DmaSg_l760_1) begin
          b2m_fsm_arbiter_logic_valid <= 1'b1;
          if(when_DmaSg_l763_4) begin
            b2m_fsm_arbiter_logic_priority_roundRobins_0 <= b2m_fsm_arbiter_logic_priority_contextNext;
          end
          if(when_DmaSg_l763_5) begin
            b2m_fsm_arbiter_logic_priority_roundRobins_1 <= b2m_fsm_arbiter_logic_priority_contextNext;
          end
          if(when_DmaSg_l763_6) begin
            b2m_fsm_arbiter_logic_priority_roundRobins_2 <= b2m_fsm_arbiter_logic_priority_contextNext;
          end
          if(when_DmaSg_l763_7) begin
            b2m_fsm_arbiter_logic_priority_roundRobins_3 <= b2m_fsm_arbiter_logic_priority_contextNext;
          end
          b2m_fsm_arbiter_logic_priority_counter <= (b2m_fsm_arbiter_logic_priority_counter + 2'b01);
          if(b2m_fsm_arbiter_logic_priority_weightLast) begin
            b2m_fsm_arbiter_logic_priority_counter <= 2'b00;
          end
        end
      end
      if(b2m_fsm_sel_ready) begin
        b2m_fsm_sel_valid <= 1'b0;
        if(b2m_fsm_sel_valid) begin
          b2m_fsm_arbiter_logic_valid <= 1'b0;
        end
      end
      if(when_DmaSg_l935) begin
        b2m_fsm_sel_valid <= 1'b1;
      end
      b2m_fsm_sel_valid_regNext <= b2m_fsm_sel_valid;
      b2m_fsm_s1 <= b2m_fsm_s0;
      if(b2m_fsm_s1) begin
        b2m_fsm_s2 <= 1'b1;
      end
      if(when_DmaSg_l986) begin
        b2m_fsm_s2 <= 1'b0;
      end
      if(when_DmaSg_l1013) begin
        b2m_fsm_toggle <= (! b2m_fsm_toggle);
      end
      if(memory_core_io_reads_2_rsp_valid) begin
        memory_core_io_reads_2_rsp_rValidN <= 1'b0;
      end
      if(memory_core_io_reads_2_rsp_s2mPipe_ready) begin
        memory_core_io_reads_2_rsp_rValidN <= 1'b1;
      end
      _zz_io_flush <= (b2m_fsm_sel_valid && (! b2m_fsm_sel_ready));
      if(io_write_cmd_fire) begin
        io_write_cmd_payload_first <= io_write_cmd_payload_last;
      end
      if(when_BusSlaveFactory_l377_1) begin
        if(when_BusSlaveFactory_l379_1) begin
          channels_0_ctrl_kick <= _zz_channels_0_ctrl_kick[0];
        end
      end
      if(when_BusSlaveFactory_l341) begin
        if(when_BusSlaveFactory_l347) begin
          channels_0_interrupts_completion_valid <= _zz_channels_0_interrupts_completion_valid[0];
        end
      end
      if(when_BusSlaveFactory_l341_1) begin
        if(when_BusSlaveFactory_l347_1) begin
          channels_0_interrupts_onChannelCompletion_valid <= _zz_channels_0_interrupts_onChannelCompletion_valid[0];
        end
      end
      if(when_BusSlaveFactory_l341_2) begin
        if(when_BusSlaveFactory_l347_2) begin
          channels_0_interrupts_s2mPacket_valid <= _zz_channels_0_interrupts_s2mPacket_valid[0];
        end
      end
      if(when_BusSlaveFactory_l377_3) begin
        if(when_BusSlaveFactory_l379_3) begin
          channels_1_ctrl_kick <= _zz_channels_1_ctrl_kick[0];
        end
      end
      if(when_BusSlaveFactory_l341_3) begin
        if(when_BusSlaveFactory_l347_3) begin
          channels_1_interrupts_completion_valid <= _zz_channels_1_interrupts_completion_valid[0];
        end
      end
      if(when_BusSlaveFactory_l341_4) begin
        if(when_BusSlaveFactory_l347_4) begin
          channels_1_interrupts_onChannelCompletion_valid <= _zz_channels_1_interrupts_onChannelCompletion_valid[0];
        end
      end
      if(when_BusSlaveFactory_l377_5) begin
        if(when_BusSlaveFactory_l379_5) begin
          channels_2_ctrl_kick <= _zz_channels_2_ctrl_kick[0];
        end
      end
      if(when_BusSlaveFactory_l341_5) begin
        if(when_BusSlaveFactory_l347_5) begin
          channels_2_interrupts_completion_valid <= _zz_channels_2_interrupts_completion_valid[0];
        end
      end
      if(when_BusSlaveFactory_l341_6) begin
        if(when_BusSlaveFactory_l347_6) begin
          channels_2_interrupts_onChannelCompletion_valid <= _zz_channels_2_interrupts_onChannelCompletion_valid[0];
        end
      end
      if(when_BusSlaveFactory_l341_7) begin
        if(when_BusSlaveFactory_l347_7) begin
          channels_2_interrupts_s2mPacket_valid <= _zz_channels_2_interrupts_s2mPacket_valid[0];
        end
      end
      if(when_BusSlaveFactory_l377_7) begin
        if(when_BusSlaveFactory_l379_7) begin
          channels_3_ctrl_kick <= _zz_channels_3_ctrl_kick[0];
        end
      end
      if(when_BusSlaveFactory_l341_8) begin
        if(when_BusSlaveFactory_l347_8) begin
          channels_3_interrupts_completion_valid <= _zz_channels_3_interrupts_completion_valid[0];
        end
      end
      if(when_BusSlaveFactory_l341_9) begin
        if(when_BusSlaveFactory_l347_9) begin
          channels_3_interrupts_onChannelCompletion_valid <= _zz_channels_3_interrupts_onChannelCompletion_valid[0];
        end
      end
      case(io_ctrl_PADDR)
        14'h0044 : begin
          if(ctrl_doWrite) begin
            channels_0_priority <= io_ctrl_PWDATA[1 : 0];
            channels_0_weight <= io_ctrl_PWDATA[9 : 8];
          end
        end
        14'h0050 : begin
          if(ctrl_doWrite) begin
            channels_0_interrupts_completion_enable <= io_ctrl_PWDATA[0];
            channels_0_interrupts_onChannelCompletion_enable <= io_ctrl_PWDATA[2];
            channels_0_interrupts_s2mPacket_enable <= io_ctrl_PWDATA[4];
          end
        end
        14'h00c4 : begin
          if(ctrl_doWrite) begin
            channels_1_priority <= io_ctrl_PWDATA[1 : 0];
            channels_1_weight <= io_ctrl_PWDATA[9 : 8];
          end
        end
        14'h00d0 : begin
          if(ctrl_doWrite) begin
            channels_1_interrupts_completion_enable <= io_ctrl_PWDATA[0];
            channels_1_interrupts_onChannelCompletion_enable <= io_ctrl_PWDATA[2];
          end
        end
        14'h0144 : begin
          if(ctrl_doWrite) begin
            channels_2_priority <= io_ctrl_PWDATA[1 : 0];
            channels_2_weight <= io_ctrl_PWDATA[9 : 8];
          end
        end
        14'h0150 : begin
          if(ctrl_doWrite) begin
            channels_2_interrupts_completion_enable <= io_ctrl_PWDATA[0];
            channels_2_interrupts_onChannelCompletion_enable <= io_ctrl_PWDATA[2];
            channels_2_interrupts_s2mPacket_enable <= io_ctrl_PWDATA[4];
          end
        end
        14'h01c4 : begin
          if(ctrl_doWrite) begin
            channels_3_priority <= io_ctrl_PWDATA[1 : 0];
            channels_3_weight <= io_ctrl_PWDATA[9 : 8];
          end
        end
        14'h01d0 : begin
          if(ctrl_doWrite) begin
            channels_3_interrupts_completion_enable <= io_ctrl_PWDATA[0];
            channels_3_interrupts_onChannelCompletion_enable <= io_ctrl_PWDATA[2];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    channels_0_fifo_push_ptr <= (channels_0_fifo_push_ptr + channels_0_fifo_push_ptrIncr_value);
    if(channels_0_channelStart) begin
      channels_0_fifo_push_ptr <= 14'h0;
    end
    channels_0_fifo_pop_ptr <= (channels_0_fifo_pop_ptr + channels_0_fifo_pop_ptrIncr_value);
    channels_0_fifo_pop_withOverride_backup <= channels_0_fifo_pop_withOverride_backupNext;
    if(when_DmaSg_l409) begin
      channels_0_fifo_pop_withOverride_valid <= 1'b0;
    end
    if(channels_0_fifo_pop_withOverride_load) begin
      channels_0_fifo_pop_withOverride_valid <= 1'b1;
    end
    channels_0_fifo_pop_withOverride_exposed <= ((! channels_0_fifo_pop_withOverride_valid) ? channels_0_fifo_pop_withOverride_backupNext : _zz_channels_0_fifo_pop_withOverride_exposed);
    if(channels_0_channelStart) begin
      channels_0_fifo_pop_withOverride_backup <= 18'h0;
      channels_0_fifo_pop_withOverride_valid <= 1'b0;
    end
    if(channels_0_channelStart) begin
      channels_0_push_s2b_packetLock <= 1'b0;
    end
    if(channels_0_pop_b2m_fire) begin
      channels_0_pop_b2m_flush <= 1'b0;
    end
    if(when_DmaSg_l505) begin
      channels_0_pop_b2m_packet <= 1'b0;
    end
    if(when_DmaSg_l523) begin
      channels_0_pop_b2m_flush <= 1'b0;
      channels_0_pop_b2m_packet <= 1'b0;
    end
    if(channels_0_pop_b2m_packetSync) begin
      channels_0_push_s2b_packetLock <= 1'b0;
    end
    if(channels_0_channelStart) begin
      channels_0_pop_b2m_bytesToSkip <= 5'h0;
      channels_0_pop_b2m_flush <= 1'b0;
    end
    if(channels_0_descriptorStart) begin
      channels_0_pop_b2m_bytesLeft <= {1'd0, channels_0_bytes};
      channels_0_pop_b2m_waitFinalRsp <= 1'b0;
    end
    if(channels_0_channelValid) begin
      if(!channels_0_channelStop) begin
        if(when_DmaSg_l575) begin
          if(when_DmaSg_l578) begin
            channels_0_pop_b2m_address <= (_zz_channels_0_pop_b2m_address - 32'h00000001);
          end
          if(when_DmaSg_l593) begin
            channels_0_channelStop <= 1'b1;
          end
        end
      end
    end
    channels_0_fifo_pop_ptrIncr_value_regNext <= channels_0_fifo_pop_ptrIncr_value;
    channels_0_fifo_push_available <= (_zz_channels_0_fifo_push_available - (channels_0_push_memory ? channels_0_fifo_push_availableDecr : channels_0_fifo_push_ptrIncr_value));
    if(channels_0_channelStart) begin
      channels_0_fifo_push_ptr <= 14'h0;
      channels_0_fifo_push_available <= (channels_0_fifo_words + 14'h0001);
      channels_0_fifo_pop_ptr <= 14'h0;
    end
    channels_1_fifo_push_ptr <= (channels_1_fifo_push_ptr + channels_1_fifo_push_ptrIncr_value);
    if(channels_1_channelStart) begin
      channels_1_fifo_push_ptr <= 14'h0;
    end
    channels_1_fifo_pop_ptr <= (channels_1_fifo_pop_ptr + channels_1_fifo_pop_ptrIncr_value);
    channels_1_fifo_pop_withoutOverride_exposed <= (_zz_channels_1_fifo_pop_withoutOverride_exposed - channels_1_fifo_pop_bytesDecr_value);
    if(channels_1_channelStart) begin
      channels_1_fifo_pop_withoutOverride_exposed <= 18'h0;
    end
    if(channels_1_descriptorStart) begin
      channels_1_push_m2b_bytesLeft <= channels_1_bytes;
    end
    if(when_DmaSg_l474) begin
      channels_1_pop_b2s_veryLastValid <= 1'b1;
    end
    if(channels_1_pop_b2s_veryLastTrigger) begin
      channels_1_pop_b2s_veryLastPtr <= channels_1_fifo_push_ptrWithBase;
      channels_1_pop_b2s_veryLastEndPacket <= channels_1_pop_b2s_last;
    end
    if(channels_1_channelStart) begin
      channels_1_pop_b2s_veryLastValid <= 1'b0;
    end
    if(channels_1_channelValid) begin
      if(!channels_1_channelStop) begin
        if(when_DmaSg_l575_1) begin
          if(when_DmaSg_l578_1) begin
            channels_1_push_m2b_address <= (_zz_channels_1_push_m2b_address - 32'h00000001);
          end
          if(when_DmaSg_l593_1) begin
            channels_1_channelStop <= 1'b1;
          end
        end
      end
    end
    channels_1_fifo_pop_ptrIncr_value_regNext <= channels_1_fifo_pop_ptrIncr_value;
    channels_1_fifo_push_available <= (_zz_channels_1_fifo_push_available - (channels_1_push_memory ? channels_1_fifo_push_availableDecr : channels_1_fifo_push_ptrIncr_value));
    if(channels_1_channelStart) begin
      channels_1_fifo_push_ptr <= 14'h0;
      channels_1_fifo_push_available <= (channels_1_fifo_words + 14'h0001);
      channels_1_fifo_pop_ptr <= 14'h0;
    end
    channels_2_fifo_push_ptr <= (channels_2_fifo_push_ptr + channels_2_fifo_push_ptrIncr_value);
    if(channels_2_channelStart) begin
      channels_2_fifo_push_ptr <= 14'h0;
    end
    channels_2_fifo_pop_ptr <= (channels_2_fifo_pop_ptr + channels_2_fifo_pop_ptrIncr_value);
    channels_2_fifo_pop_withOverride_backup <= channels_2_fifo_pop_withOverride_backupNext;
    if(when_DmaSg_l409_1) begin
      channels_2_fifo_pop_withOverride_valid <= 1'b0;
    end
    if(channels_2_fifo_pop_withOverride_load) begin
      channels_2_fifo_pop_withOverride_valid <= 1'b1;
    end
    channels_2_fifo_pop_withOverride_exposed <= ((! channels_2_fifo_pop_withOverride_valid) ? channels_2_fifo_pop_withOverride_backupNext : _zz_channels_2_fifo_pop_withOverride_exposed);
    if(channels_2_channelStart) begin
      channels_2_fifo_pop_withOverride_backup <= 18'h0;
      channels_2_fifo_pop_withOverride_valid <= 1'b0;
    end
    if(channels_2_channelStart) begin
      channels_2_push_s2b_packetLock <= 1'b0;
    end
    if(channels_2_pop_b2m_fire) begin
      channels_2_pop_b2m_flush <= 1'b0;
    end
    if(when_DmaSg_l505_1) begin
      channels_2_pop_b2m_packet <= 1'b0;
    end
    if(when_DmaSg_l523_1) begin
      channels_2_pop_b2m_flush <= 1'b0;
      channels_2_pop_b2m_packet <= 1'b0;
    end
    if(channels_2_pop_b2m_packetSync) begin
      channels_2_push_s2b_packetLock <= 1'b0;
    end
    if(channels_2_channelStart) begin
      channels_2_pop_b2m_bytesToSkip <= 5'h0;
      channels_2_pop_b2m_flush <= 1'b0;
    end
    if(channels_2_descriptorStart) begin
      channels_2_pop_b2m_bytesLeft <= {1'd0, channels_2_bytes};
      channels_2_pop_b2m_waitFinalRsp <= 1'b0;
    end
    if(channels_2_channelValid) begin
      if(!channels_2_channelStop) begin
        if(when_DmaSg_l575_2) begin
          if(when_DmaSg_l578_2) begin
            channels_2_pop_b2m_address <= (_zz_channels_2_pop_b2m_address - 32'h00000001);
          end
          if(when_DmaSg_l593_2) begin
            channels_2_channelStop <= 1'b1;
          end
        end
      end
    end
    channels_2_fifo_pop_ptrIncr_value_regNext <= channels_2_fifo_pop_ptrIncr_value;
    channels_2_fifo_push_available <= (_zz_channels_2_fifo_push_available - (channels_2_push_memory ? channels_2_fifo_push_availableDecr : channels_2_fifo_push_ptrIncr_value));
    if(channels_2_channelStart) begin
      channels_2_fifo_push_ptr <= 14'h0;
      channels_2_fifo_push_available <= (channels_2_fifo_words + 14'h0001);
      channels_2_fifo_pop_ptr <= 14'h0;
    end
    channels_3_fifo_push_ptr <= (channels_3_fifo_push_ptr + channels_3_fifo_push_ptrIncr_value);
    if(channels_3_channelStart) begin
      channels_3_fifo_push_ptr <= 14'h0;
    end
    channels_3_fifo_pop_ptr <= (channels_3_fifo_pop_ptr + channels_3_fifo_pop_ptrIncr_value);
    channels_3_fifo_pop_withoutOverride_exposed <= (_zz_channels_3_fifo_pop_withoutOverride_exposed - channels_3_fifo_pop_bytesDecr_value);
    if(channels_3_channelStart) begin
      channels_3_fifo_pop_withoutOverride_exposed <= 18'h0;
    end
    if(channels_3_descriptorStart) begin
      channels_3_push_m2b_bytesLeft <= channels_3_bytes;
    end
    if(when_DmaSg_l474_1) begin
      channels_3_pop_b2s_veryLastValid <= 1'b1;
    end
    if(channels_3_pop_b2s_veryLastTrigger) begin
      channels_3_pop_b2s_veryLastPtr <= channels_3_fifo_push_ptrWithBase;
      channels_3_pop_b2s_veryLastEndPacket <= channels_3_pop_b2s_last;
    end
    if(channels_3_channelStart) begin
      channels_3_pop_b2s_veryLastValid <= 1'b0;
    end
    if(channels_3_channelValid) begin
      if(!channels_3_channelStop) begin
        if(when_DmaSg_l575_3) begin
          if(when_DmaSg_l578_3) begin
            channels_3_push_m2b_address <= (_zz_channels_3_push_m2b_address - 32'h00000001);
          end
          if(when_DmaSg_l593_3) begin
            channels_3_channelStop <= 1'b1;
          end
        end
      end
    end
    channels_3_fifo_pop_ptrIncr_value_regNext <= channels_3_fifo_pop_ptrIncr_value;
    channels_3_fifo_push_available <= (_zz_channels_3_fifo_push_available - (channels_3_push_memory ? channels_3_fifo_push_availableDecr : channels_3_fifo_push_ptrIncr_value));
    if(channels_3_channelStart) begin
      channels_3_fifo_push_ptr <= 14'h0;
      channels_3_fifo_push_available <= (channels_3_fifo_words + 14'h0001);
      channels_3_fifo_pop_ptr <= 14'h0;
    end
    if(when_DmaSg_l665) begin
      channels_0_push_s2b_waitFirst <= 1'b0;
      if(io_inputs_0_payload_last) begin
        channels_0_push_s2b_packetLock <= 1'b1;
      end
    end
    if(when_DmaSg_l681) begin
      channels_0_pop_b2m_flush <= 1'b1;
    end
    if(when_DmaSg_l682) begin
      channels_0_pop_b2m_packet <= 1'b1;
    end
    if(when_DmaSg_l665_1) begin
      channels_2_push_s2b_waitFirst <= 1'b0;
      if(io_inputs_1_payload_last) begin
        channels_2_push_s2b_packetLock <= 1'b1;
      end
    end
    if(when_DmaSg_l681_1) begin
      channels_2_pop_b2m_flush <= 1'b1;
    end
    if(when_DmaSg_l682_1) begin
      channels_2_pop_b2m_packet <= 1'b1;
    end
    if(when_DmaSg_l725) begin
      if(when_DmaSg_l726) begin
        channels_1_pop_b2s_veryLastValid <= 1'b0;
      end
    end
    if(when_DmaSg_l725_1) begin
      if(when_DmaSg_l726_1) begin
        channels_3_pop_b2s_veryLastValid <= 1'b0;
      end
    end
    if(when_DmaSg_l758) begin
      m2b_cmd_s0_chosen <= m2b_cmd_s0_priority_chosen;
    end
    m2b_cmd_s1_address <= m2b_cmd_s0_address;
    m2b_cmd_s1_length <= m2b_cmd_s0_length;
    m2b_cmd_s1_lastBurst <= m2b_cmd_s0_lastBurst;
    m2b_cmd_s1_bytesLeft <= m2b_cmd_s0_bytesLeft;
    if(m2b_cmd_s1_valid) begin
      if(io_read_cmd_ready) begin
        if(when_DmaSg_l828) begin
          channels_1_push_m2b_address <= m2b_cmd_s1_addressNext;
          channels_1_push_m2b_bytesLeft <= m2b_cmd_s1_byteLeftNext;
        end
        if(when_DmaSg_l828_1) begin
          channels_3_push_m2b_address <= m2b_cmd_s1_addressNext;
          channels_3_push_m2b_bytesLeft <= m2b_cmd_s1_byteLeftNext;
        end
      end
    end
    if(when_DmaSg_l758_1) begin
      b2m_fsm_arbiter_logic_chosen <= b2m_fsm_arbiter_logic_priority_chosen;
    end
    if(when_DmaSg_l935) begin
      b2m_fsm_sel_channel <= b2m_fsm_arbiter_logic_chosen;
      b2m_fsm_sel_address <= _zz_b2m_fsm_sel_address;
      b2m_fsm_sel_ptr <= _zz_b2m_fsm_sel_ptr;
      b2m_fsm_sel_ptrMask <= _zz_b2m_fsm_sel_ptrMask;
      b2m_fsm_sel_bytePerBurst <= _zz_b2m_fsm_sel_bytePerBurst;
      b2m_fsm_sel_bytesInFifo <= _zz_b2m_fsm_sel_bytesInFifo;
      b2m_fsm_sel_flush <= _zz_b2m_fsm_sel_flush;
      b2m_fsm_sel_packet <= _zz_b2m_fsm_sel_packet;
      b2m_fsm_sel_bytesLeft <= _zz_b2m_fsm_sel_bytesLeft[25:0];
    end
    if(b2m_fsm_s0) begin
      b2m_fsm_sel_bytesInBurst <= _zz_b2m_fsm_sel_bytesInBurst_3[12:0];
    end
    if(b2m_fsm_s1) begin
      b2m_fsm_beatCounter <= (_zz_b2m_fsm_beatCounter >>> 3'd5);
      if(when_DmaSg_l996) begin
        channels_0_pop_b2m_address <= b2m_fsm_addressNext;
        channels_0_pop_b2m_bytesLeft <= b2m_fsm_bytesLeftNext;
        if(b2m_fsm_isFinalCmd) begin
          channels_0_pop_b2m_waitFinalRsp <= 1'b1;
        end
        if(when_DmaSg_l1001) begin
          if(b2m_fsm_sel_flush) begin
            channels_0_pop_b2m_flush <= 1'b1;
          end
          if(b2m_fsm_sel_packet) begin
            channels_0_pop_b2m_packet <= 1'b1;
          end
        end
      end
      if(when_DmaSg_l996_1) begin
        channels_2_pop_b2m_address <= b2m_fsm_addressNext;
        channels_2_pop_b2m_bytesLeft <= b2m_fsm_bytesLeftNext;
        if(b2m_fsm_isFinalCmd) begin
          channels_2_pop_b2m_waitFinalRsp <= 1'b1;
        end
        if(when_DmaSg_l1001_1) begin
          if(b2m_fsm_sel_flush) begin
            channels_2_pop_b2m_flush <= 1'b1;
          end
          if(b2m_fsm_sel_packet) begin
            channels_2_pop_b2m_packet <= 1'b1;
          end
        end
      end
    end
    if(when_DmaSg_l1033) begin
      b2m_fsm_sel_ptr <= ((b2m_fsm_sel_ptr & (~ b2m_fsm_sel_ptrMask)) | (_zz_b2m_fsm_sel_ptr_1 & b2m_fsm_sel_ptrMask));
    end
    if(memory_core_io_reads_2_rsp_rValidN) begin
      memory_core_io_reads_2_rsp_rData_data <= memory_core_io_reads_2_rsp_payload_data;
      memory_core_io_reads_2_rsp_rData_mask <= memory_core_io_reads_2_rsp_payload_mask;
      memory_core_io_reads_2_rsp_rData_context <= memory_core_io_reads_2_rsp_payload_context;
    end
    if(b2m_fsm_aggregate_memoryPort_fire) begin
      b2m_fsm_aggregate_first <= 1'b0;
    end
    if(when_DmaSg_l1050) begin
      b2m_fsm_aggregate_first <= 1'b1;
    end
    b2m_fsm_cmd_maskLastTriggerReg <= b2m_fsm_cmd_maskLastTriggerComb;
    b2m_fsm_cmd_maskLast <= {(5'h1f <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h1e <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h1d <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h1c <= b2m_fsm_cmd_maskLastTriggerComb),{(5'h1b <= b2m_fsm_cmd_maskLastTriggerComb),{(_zz_b2m_fsm_cmd_maskLast <= b2m_fsm_cmd_maskLastTriggerComb),{_zz_b2m_fsm_cmd_maskLast_1,{_zz_b2m_fsm_cmd_maskLast_2,_zz_b2m_fsm_cmd_maskLast_3}}}}}}}};
    if(io_write_cmd_fire) begin
      b2m_fsm_beatCounter <= (b2m_fsm_beatCounter - 8'h01);
    end
    if(when_DmaSg_l1102) begin
      if(_zz_2[0]) begin
        channels_0_pop_b2m_bytesToSkip <= _zz_channels_0_pop_b2m_bytesToSkip;
      end
      if(_zz_2[1]) begin
        channels_2_pop_b2m_bytesToSkip <= _zz_channels_0_pop_b2m_bytesToSkip;
      end
    end
    case(io_ctrl_PADDR)
      14'h000c : begin
        if(ctrl_doWrite) begin
          channels_0_push_memory <= io_ctrl_PWDATA[12];
          channels_0_push_s2b_completionOnLast <= io_ctrl_PWDATA[13];
          channels_0_push_s2b_waitFirst <= io_ctrl_PWDATA[14];
        end
      end
      14'h001c : begin
        if(ctrl_doWrite) begin
          channels_0_pop_memory <= io_ctrl_PWDATA[12];
        end
      end
      14'h002c : begin
        if(ctrl_doWrite) begin
          channels_0_channelStop <= io_ctrl_PWDATA[2];
          channels_0_selfRestart <= io_ctrl_PWDATA[1];
        end
      end
      14'h0020 : begin
        if(ctrl_doWrite) begin
          channels_0_bytes <= io_ctrl_PWDATA[25 : 0];
        end
      end
      14'h008c : begin
        if(ctrl_doWrite) begin
          channels_1_push_memory <= io_ctrl_PWDATA[12];
        end
      end
      14'h0098 : begin
        if(ctrl_doWrite) begin
          channels_1_pop_b2s_portId <= io_ctrl_PWDATA[0 : 0];
          channels_1_pop_b2s_sinkId <= io_ctrl_PWDATA[19 : 16];
        end
      end
      14'h009c : begin
        if(ctrl_doWrite) begin
          channels_1_pop_memory <= io_ctrl_PWDATA[12];
          channels_1_pop_b2s_last <= io_ctrl_PWDATA[13];
        end
      end
      14'h00ac : begin
        if(ctrl_doWrite) begin
          channels_1_channelStop <= io_ctrl_PWDATA[2];
          channels_1_selfRestart <= io_ctrl_PWDATA[1];
        end
      end
      14'h00a0 : begin
        if(ctrl_doWrite) begin
          channels_1_bytes <= io_ctrl_PWDATA[25 : 0];
        end
      end
      14'h010c : begin
        if(ctrl_doWrite) begin
          channels_2_push_memory <= io_ctrl_PWDATA[12];
          channels_2_push_s2b_completionOnLast <= io_ctrl_PWDATA[13];
          channels_2_push_s2b_waitFirst <= io_ctrl_PWDATA[14];
        end
      end
      14'h011c : begin
        if(ctrl_doWrite) begin
          channels_2_pop_memory <= io_ctrl_PWDATA[12];
        end
      end
      14'h012c : begin
        if(ctrl_doWrite) begin
          channels_2_channelStop <= io_ctrl_PWDATA[2];
          channels_2_selfRestart <= io_ctrl_PWDATA[1];
        end
      end
      14'h0120 : begin
        if(ctrl_doWrite) begin
          channels_2_bytes <= io_ctrl_PWDATA[25 : 0];
        end
      end
      14'h018c : begin
        if(ctrl_doWrite) begin
          channels_3_push_memory <= io_ctrl_PWDATA[12];
        end
      end
      14'h0198 : begin
        if(ctrl_doWrite) begin
          channels_3_pop_b2s_portId <= io_ctrl_PWDATA[0 : 0];
          channels_3_pop_b2s_sinkId <= io_ctrl_PWDATA[19 : 16];
        end
      end
      14'h019c : begin
        if(ctrl_doWrite) begin
          channels_3_pop_memory <= io_ctrl_PWDATA[12];
          channels_3_pop_b2s_last <= io_ctrl_PWDATA[13];
        end
      end
      14'h01ac : begin
        if(ctrl_doWrite) begin
          channels_3_channelStop <= io_ctrl_PWDATA[2];
          channels_3_selfRestart <= io_ctrl_PWDATA[1];
        end
      end
      14'h01a0 : begin
        if(ctrl_doWrite) begin
          channels_3_bytes <= io_ctrl_PWDATA[25 : 0];
        end
      end
      default : begin
      end
    endcase
    if(when_Apb3SlaveFactory_l81) begin
      if(ctrl_doWrite) begin
        channels_0_pop_b2m_address[31 : 0] <= io_ctrl_PWDATA[31 : 0];
      end
    end
    if(when_Apb3SlaveFactory_l81_1) begin
      if(ctrl_doWrite) begin
        channels_1_push_m2b_address[31 : 0] <= io_ctrl_PWDATA[31 : 0];
      end
    end
    if(when_Apb3SlaveFactory_l81_2) begin
      if(ctrl_doWrite) begin
        channels_2_pop_b2m_address[31 : 0] <= io_ctrl_PWDATA[31 : 0];
      end
    end
    if(when_Apb3SlaveFactory_l81_3) begin
      if(ctrl_doWrite) begin
        channels_3_push_m2b_address[31 : 0] <= io_ctrl_PWDATA[31 : 0];
      end
    end
  end


endmodule

module EfxDMA_BufferCC_9 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          dat3_o_clk,
  input  wire          dat3_o_reset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge dat3_o_clk) begin
    if(dat3_o_reset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//EfxDMA_BufferCC_8 replaced by EfxDMA_BufferCC_3

module EfxDMA_BufferCC_7 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          dat1_o_clk,
  input  wire          dat1_o_reset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge dat1_o_clk) begin
    if(dat1_o_reset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//EfxDMA_BufferCC_6 replaced by EfxDMA_BufferCC_3

//EfxDMA_BufferCC_5 replaced by EfxDMA_BufferCC_3

module EfxDMA_BufferCC_4 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          dat2_i_clk,
  input  wire          dat2_i_reset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge dat2_i_clk) begin
    if(dat2_i_reset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module EfxDMA_BufferCC_3 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          clk,
  input  wire          reset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk) begin
    if(reset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module EfxDMA_BufferCC_2 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          dat0_i_clk,
  input  wire          dat0_i_reset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge dat0_i_clk) begin
    if(dat0_i_reset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module EfxDMA_BmbContextRemover_1 (
  input  wire          io_input_cmd_valid,
  output reg           io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [12:0]   io_input_cmd_payload_fragment_length,
  input  wire [255:0]  io_input_cmd_payload_fragment_data,
  input  wire [31:0]   io_input_cmd_payload_fragment_mask,
  input  wire [15:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [15:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [12:0]   io_output_cmd_payload_fragment_length,
  output wire [255:0]  io_output_cmd_payload_fragment_data,
  output wire [31:0]   io_output_cmd_payload_fragment_mask,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire          clk,
  input  wire          reset
);

  reg                 fifoFork_thrown_translated_fifo_io_pop_ready;
  wire                fifoFork_thrown_translated_fifo_io_push_ready;
  wire                fifoFork_thrown_translated_fifo_io_pop_valid;
  wire       [15:0]   fifoFork_thrown_translated_fifo_io_pop_payload_context;
  wire       [2:0]    fifoFork_thrown_translated_fifo_io_occupancy;
  wire       [2:0]    fifoFork_thrown_translated_fifo_io_availability;
  wire                fifoFork_valid;
  reg                 fifoFork_ready;
  wire                fifoFork_payload_last;
  wire       [0:0]    fifoFork_payload_fragment_opcode;
  wire       [31:0]   fifoFork_payload_fragment_address;
  wire       [12:0]   fifoFork_payload_fragment_length;
  wire       [255:0]  fifoFork_payload_fragment_data;
  wire       [31:0]   fifoFork_payload_fragment_mask;
  wire       [15:0]   fifoFork_payload_fragment_context;
  wire                cmdFork_valid;
  wire                cmdFork_ready;
  wire                cmdFork_payload_last;
  wire       [0:0]    cmdFork_payload_fragment_opcode;
  wire       [31:0]   cmdFork_payload_fragment_address;
  wire       [12:0]   cmdFork_payload_fragment_length;
  wire       [255:0]  cmdFork_payload_fragment_data;
  wire       [31:0]   cmdFork_payload_fragment_mask;
  wire       [15:0]   cmdFork_payload_fragment_context;
  reg                 io_input_cmd_fork2_logic_linkEnable_0;
  reg                 io_input_cmd_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                fifoFork_fire;
  wire                cmdFork_fire;
  wire       [15:0]   pushCtx_context;
  reg                 fifoFork_payload_first;
  wire                when_Stream_l445;
  reg                 fifoFork_thrown_valid;
  wire                fifoFork_thrown_ready;
  wire                fifoFork_thrown_payload_last;
  wire       [0:0]    fifoFork_thrown_payload_fragment_opcode;
  wire       [31:0]   fifoFork_thrown_payload_fragment_address;
  wire       [12:0]   fifoFork_thrown_payload_fragment_length;
  wire       [255:0]  fifoFork_thrown_payload_fragment_data;
  wire       [31:0]   fifoFork_thrown_payload_fragment_mask;
  wire       [15:0]   fifoFork_thrown_payload_fragment_context;
  wire                fifoFork_thrown_translated_valid;
  wire                fifoFork_thrown_translated_ready;
  wire       [15:0]   fifoFork_thrown_translated_payload_context;
  wire                popCtx_valid;
  wire                popCtx_ready;
  wire       [15:0]   popCtx_payload_context;
  reg                 fifoFork_thrown_translated_fifo_io_pop_rValid;
  reg        [15:0]   fifoFork_thrown_translated_fifo_io_pop_rData_context;
  wire                when_Stream_l375;
  wire                _zz_io_input_rsp_valid;

  EfxDMA_StreamFifo_1 fifoFork_thrown_translated_fifo (
    .io_push_valid           (fifoFork_thrown_translated_valid                            ), //i
    .io_push_ready           (fifoFork_thrown_translated_fifo_io_push_ready               ), //o
    .io_push_payload_context (fifoFork_thrown_translated_payload_context[15:0]            ), //i
    .io_pop_valid            (fifoFork_thrown_translated_fifo_io_pop_valid                ), //o
    .io_pop_ready            (fifoFork_thrown_translated_fifo_io_pop_ready                ), //i
    .io_pop_payload_context  (fifoFork_thrown_translated_fifo_io_pop_payload_context[15:0]), //o
    .io_flush                (1'b0                                                        ), //i
    .io_occupancy            (fifoFork_thrown_translated_fifo_io_occupancy[2:0]           ), //o
    .io_availability         (fifoFork_thrown_translated_fifo_io_availability[2:0]        ), //o
    .clk                     (clk                                                         ), //i
    .reset                   (reset                                                       )  //i
  );
  always @(*) begin
    io_input_cmd_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_input_cmd_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_input_cmd_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! fifoFork_ready) && io_input_cmd_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdFork_ready) && io_input_cmd_fork2_logic_linkEnable_1);
  assign fifoFork_valid = (io_input_cmd_valid && io_input_cmd_fork2_logic_linkEnable_0);
  assign fifoFork_payload_last = io_input_cmd_payload_last;
  assign fifoFork_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign fifoFork_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign fifoFork_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign fifoFork_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign fifoFork_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign fifoFork_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign fifoFork_fire = (fifoFork_valid && fifoFork_ready);
  assign cmdFork_valid = (io_input_cmd_valid && io_input_cmd_fork2_logic_linkEnable_1);
  assign cmdFork_payload_last = io_input_cmd_payload_last;
  assign cmdFork_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign cmdFork_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign cmdFork_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign cmdFork_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign cmdFork_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign cmdFork_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign cmdFork_fire = (cmdFork_valid && cmdFork_ready);
  assign io_output_cmd_valid = cmdFork_valid;
  assign cmdFork_ready = io_output_cmd_ready;
  assign io_output_cmd_payload_last = cmdFork_payload_last;
  assign io_output_cmd_payload_fragment_opcode = cmdFork_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = cmdFork_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = cmdFork_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = cmdFork_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = cmdFork_payload_fragment_mask;
  assign pushCtx_context = fifoFork_payload_fragment_context;
  assign when_Stream_l445 = (! fifoFork_payload_first);
  always @(*) begin
    fifoFork_thrown_valid = fifoFork_valid;
    if(when_Stream_l445) begin
      fifoFork_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    fifoFork_ready = fifoFork_thrown_ready;
    if(when_Stream_l445) begin
      fifoFork_ready = 1'b1;
    end
  end

  assign fifoFork_thrown_payload_last = fifoFork_payload_last;
  assign fifoFork_thrown_payload_fragment_opcode = fifoFork_payload_fragment_opcode;
  assign fifoFork_thrown_payload_fragment_address = fifoFork_payload_fragment_address;
  assign fifoFork_thrown_payload_fragment_length = fifoFork_payload_fragment_length;
  assign fifoFork_thrown_payload_fragment_data = fifoFork_payload_fragment_data;
  assign fifoFork_thrown_payload_fragment_mask = fifoFork_payload_fragment_mask;
  assign fifoFork_thrown_payload_fragment_context = fifoFork_payload_fragment_context;
  assign fifoFork_thrown_translated_valid = fifoFork_thrown_valid;
  assign fifoFork_thrown_ready = fifoFork_thrown_translated_ready;
  assign fifoFork_thrown_translated_payload_context = pushCtx_context;
  assign fifoFork_thrown_translated_ready = fifoFork_thrown_translated_fifo_io_push_ready;
  always @(*) begin
    fifoFork_thrown_translated_fifo_io_pop_ready = popCtx_ready;
    if(when_Stream_l375) begin
      fifoFork_thrown_translated_fifo_io_pop_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCtx_valid);
  assign popCtx_valid = fifoFork_thrown_translated_fifo_io_pop_rValid;
  assign popCtx_payload_context = fifoFork_thrown_translated_fifo_io_pop_rData_context;
  assign popCtx_ready = ((io_output_rsp_valid && io_output_rsp_payload_last) && io_input_rsp_ready);
  assign _zz_io_input_rsp_valid = (! (! popCtx_valid));
  assign io_output_rsp_ready = (io_input_rsp_ready && _zz_io_input_rsp_valid);
  assign io_input_rsp_valid = (io_output_rsp_valid && _zz_io_input_rsp_valid);
  assign io_input_rsp_payload_last = io_output_rsp_payload_last;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_context = popCtx_payload_context;
  always @(posedge clk) begin
    if(reset) begin
      io_input_cmd_fork2_logic_linkEnable_0 <= 1'b1;
      io_input_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      fifoFork_payload_first <= 1'b1;
      fifoFork_thrown_translated_fifo_io_pop_rValid <= 1'b0;
    end else begin
      if(fifoFork_fire) begin
        io_input_cmd_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdFork_fire) begin
        io_input_cmd_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_cmd_ready) begin
        io_input_cmd_fork2_logic_linkEnable_0 <= 1'b1;
        io_input_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(fifoFork_fire) begin
        fifoFork_payload_first <= fifoFork_payload_last;
      end
      if(fifoFork_thrown_translated_fifo_io_pop_ready) begin
        fifoFork_thrown_translated_fifo_io_pop_rValid <= fifoFork_thrown_translated_fifo_io_pop_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(fifoFork_thrown_translated_fifo_io_pop_ready) begin
      fifoFork_thrown_translated_fifo_io_pop_rData_context <= fifoFork_thrown_translated_fifo_io_pop_payload_context;
    end
  end


endmodule

module EfxDMA_BmbContextRemover (
  input  wire          io_input_cmd_valid,
  output reg           io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [12:0]   io_input_cmd_payload_fragment_length,
  input  wire [25:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [255:0]  io_input_rsp_payload_fragment_data,
  output wire [25:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [12:0]   io_output_cmd_payload_fragment_length,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [255:0]  io_output_rsp_payload_fragment_data,
  input  wire          clk,
  input  wire          reset
);

  reg                 fifoFork_thrown_translated_fifo_io_pop_ready;
  wire                fifoFork_thrown_translated_fifo_io_push_ready;
  wire                fifoFork_thrown_translated_fifo_io_pop_valid;
  wire       [25:0]   fifoFork_thrown_translated_fifo_io_pop_payload_context;
  wire       [2:0]    fifoFork_thrown_translated_fifo_io_occupancy;
  wire       [2:0]    fifoFork_thrown_translated_fifo_io_availability;
  wire                fifoFork_valid;
  reg                 fifoFork_ready;
  wire                fifoFork_payload_last;
  wire       [0:0]    fifoFork_payload_fragment_opcode;
  wire       [31:0]   fifoFork_payload_fragment_address;
  wire       [12:0]   fifoFork_payload_fragment_length;
  wire       [25:0]   fifoFork_payload_fragment_context;
  wire                cmdFork_valid;
  wire                cmdFork_ready;
  wire                cmdFork_payload_last;
  wire       [0:0]    cmdFork_payload_fragment_opcode;
  wire       [31:0]   cmdFork_payload_fragment_address;
  wire       [12:0]   cmdFork_payload_fragment_length;
  wire       [25:0]   cmdFork_payload_fragment_context;
  reg                 io_input_cmd_fork2_logic_linkEnable_0;
  reg                 io_input_cmd_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                fifoFork_fire;
  wire                cmdFork_fire;
  wire       [25:0]   pushCtx_context;
  reg                 fifoFork_payload_first;
  wire                when_Stream_l445;
  reg                 fifoFork_thrown_valid;
  wire                fifoFork_thrown_ready;
  wire                fifoFork_thrown_payload_last;
  wire       [0:0]    fifoFork_thrown_payload_fragment_opcode;
  wire       [31:0]   fifoFork_thrown_payload_fragment_address;
  wire       [12:0]   fifoFork_thrown_payload_fragment_length;
  wire       [25:0]   fifoFork_thrown_payload_fragment_context;
  wire                fifoFork_thrown_translated_valid;
  wire                fifoFork_thrown_translated_ready;
  wire       [25:0]   fifoFork_thrown_translated_payload_context;
  wire                popCtx_valid;
  wire                popCtx_ready;
  wire       [25:0]   popCtx_payload_context;
  reg                 fifoFork_thrown_translated_fifo_io_pop_rValid;
  reg        [25:0]   fifoFork_thrown_translated_fifo_io_pop_rData_context;
  wire                when_Stream_l375;
  wire                _zz_io_input_rsp_valid;

  EfxDMA_StreamFifo fifoFork_thrown_translated_fifo (
    .io_push_valid           (fifoFork_thrown_translated_valid                            ), //i
    .io_push_ready           (fifoFork_thrown_translated_fifo_io_push_ready               ), //o
    .io_push_payload_context (fifoFork_thrown_translated_payload_context[25:0]            ), //i
    .io_pop_valid            (fifoFork_thrown_translated_fifo_io_pop_valid                ), //o
    .io_pop_ready            (fifoFork_thrown_translated_fifo_io_pop_ready                ), //i
    .io_pop_payload_context  (fifoFork_thrown_translated_fifo_io_pop_payload_context[25:0]), //o
    .io_flush                (1'b0                                                        ), //i
    .io_occupancy            (fifoFork_thrown_translated_fifo_io_occupancy[2:0]           ), //o
    .io_availability         (fifoFork_thrown_translated_fifo_io_availability[2:0]        ), //o
    .clk                     (clk                                                         ), //i
    .reset                   (reset                                                       )  //i
  );
  always @(*) begin
    io_input_cmd_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_input_cmd_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_input_cmd_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! fifoFork_ready) && io_input_cmd_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdFork_ready) && io_input_cmd_fork2_logic_linkEnable_1);
  assign fifoFork_valid = (io_input_cmd_valid && io_input_cmd_fork2_logic_linkEnable_0);
  assign fifoFork_payload_last = io_input_cmd_payload_last;
  assign fifoFork_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign fifoFork_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign fifoFork_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign fifoFork_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign fifoFork_fire = (fifoFork_valid && fifoFork_ready);
  assign cmdFork_valid = (io_input_cmd_valid && io_input_cmd_fork2_logic_linkEnable_1);
  assign cmdFork_payload_last = io_input_cmd_payload_last;
  assign cmdFork_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign cmdFork_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign cmdFork_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign cmdFork_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign cmdFork_fire = (cmdFork_valid && cmdFork_ready);
  assign io_output_cmd_valid = cmdFork_valid;
  assign cmdFork_ready = io_output_cmd_ready;
  assign io_output_cmd_payload_last = cmdFork_payload_last;
  assign io_output_cmd_payload_fragment_opcode = cmdFork_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = cmdFork_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = cmdFork_payload_fragment_length;
  assign pushCtx_context = fifoFork_payload_fragment_context;
  assign when_Stream_l445 = (! fifoFork_payload_first);
  always @(*) begin
    fifoFork_thrown_valid = fifoFork_valid;
    if(when_Stream_l445) begin
      fifoFork_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    fifoFork_ready = fifoFork_thrown_ready;
    if(when_Stream_l445) begin
      fifoFork_ready = 1'b1;
    end
  end

  assign fifoFork_thrown_payload_last = fifoFork_payload_last;
  assign fifoFork_thrown_payload_fragment_opcode = fifoFork_payload_fragment_opcode;
  assign fifoFork_thrown_payload_fragment_address = fifoFork_payload_fragment_address;
  assign fifoFork_thrown_payload_fragment_length = fifoFork_payload_fragment_length;
  assign fifoFork_thrown_payload_fragment_context = fifoFork_payload_fragment_context;
  assign fifoFork_thrown_translated_valid = fifoFork_thrown_valid;
  assign fifoFork_thrown_ready = fifoFork_thrown_translated_ready;
  assign fifoFork_thrown_translated_payload_context = pushCtx_context;
  assign fifoFork_thrown_translated_ready = fifoFork_thrown_translated_fifo_io_push_ready;
  always @(*) begin
    fifoFork_thrown_translated_fifo_io_pop_ready = popCtx_ready;
    if(when_Stream_l375) begin
      fifoFork_thrown_translated_fifo_io_pop_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCtx_valid);
  assign popCtx_valid = fifoFork_thrown_translated_fifo_io_pop_rValid;
  assign popCtx_payload_context = fifoFork_thrown_translated_fifo_io_pop_rData_context;
  assign popCtx_ready = ((io_output_rsp_valid && io_output_rsp_payload_last) && io_input_rsp_ready);
  assign _zz_io_input_rsp_valid = (! (! popCtx_valid));
  assign io_output_rsp_ready = (io_input_rsp_ready && _zz_io_input_rsp_valid);
  assign io_input_rsp_valid = (io_output_rsp_valid && _zz_io_input_rsp_valid);
  assign io_input_rsp_payload_last = io_output_rsp_payload_last;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = popCtx_payload_context;
  always @(posedge clk) begin
    if(reset) begin
      io_input_cmd_fork2_logic_linkEnable_0 <= 1'b1;
      io_input_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      fifoFork_payload_first <= 1'b1;
      fifoFork_thrown_translated_fifo_io_pop_rValid <= 1'b0;
    end else begin
      if(fifoFork_fire) begin
        io_input_cmd_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdFork_fire) begin
        io_input_cmd_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_cmd_ready) begin
        io_input_cmd_fork2_logic_linkEnable_0 <= 1'b1;
        io_input_cmd_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(fifoFork_fire) begin
        fifoFork_payload_first <= fifoFork_payload_last;
      end
      if(fifoFork_thrown_translated_fifo_io_pop_ready) begin
        fifoFork_thrown_translated_fifo_io_pop_rValid <= fifoFork_thrown_translated_fifo_io_pop_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(fifoFork_thrown_translated_fifo_io_pop_ready) begin
      fifoFork_thrown_translated_fifo_io_pop_rData_context <= fifoFork_thrown_translated_fifo_io_pop_payload_context;
    end
  end


endmodule

module EfxDMA_FlowCCUnsafeByToggle_1 (
  input  wire          io_input_valid,
  input  wire [31:0]   io_input_payload_PRDATA,
  input  wire          io_input_payload_PSLVERROR,
  output wire          io_output_valid,
  output wire [31:0]   io_output_payload_PRDATA,
  output wire          io_output_payload_PSLVERROR,
  input  wire          clk,
  input  wire          reset,
  input  wire          ctrl_clk,
  input  wire          ctrl_reset
);

  wire                inputArea_target_buffercc_io_dataOut;
  reg                 inputArea_target;
  reg        [31:0]   inputArea_data_PRDATA;
  reg                 inputArea_data_PSLVERROR;
  wire                outputArea_target;
  reg                 outputArea_hit;
  wire                outputArea_flow_valid;
  wire       [31:0]   outputArea_flow_payload_PRDATA;
  wire                outputArea_flow_payload_PSLVERROR;
  reg                 outputArea_flow_m2sPipe_valid;
  (* async_reg = "true" *) reg        [31:0]   outputArea_flow_m2sPipe_payload_PRDATA;
  (* async_reg = "true" *) reg                 outputArea_flow_m2sPipe_payload_PSLVERROR;

  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC_1 inputArea_target_buffercc (
    .io_dataIn  (inputArea_target                    ), //i
    .io_dataOut (inputArea_target_buffercc_io_dataOut), //o
    .ctrl_clk   (ctrl_clk                            ), //i
    .ctrl_reset (ctrl_reset                          )  //i
  );
  assign outputArea_target = inputArea_target_buffercc_io_dataOut;
  assign outputArea_flow_valid = (outputArea_target != outputArea_hit);
  assign outputArea_flow_payload_PRDATA = inputArea_data_PRDATA;
  assign outputArea_flow_payload_PSLVERROR = inputArea_data_PSLVERROR;
  assign io_output_valid = outputArea_flow_m2sPipe_valid;
  assign io_output_payload_PRDATA = outputArea_flow_m2sPipe_payload_PRDATA;
  assign io_output_payload_PSLVERROR = outputArea_flow_m2sPipe_payload_PSLVERROR;
  always @(posedge clk) begin
    if(reset) begin
      inputArea_target <= 1'b0;
    end else begin
      if(io_input_valid) begin
        inputArea_target <= (! inputArea_target);
      end
    end
  end

  always @(posedge clk) begin
    if(io_input_valid) begin
      inputArea_data_PRDATA <= io_input_payload_PRDATA;
      inputArea_data_PSLVERROR <= io_input_payload_PSLVERROR;
    end
  end

  always @(posedge ctrl_clk) begin
    if(ctrl_reset) begin
      outputArea_flow_m2sPipe_valid <= 1'b0;
      outputArea_hit <= 1'b0;
    end else begin
      outputArea_hit <= outputArea_target;
      outputArea_flow_m2sPipe_valid <= outputArea_flow_valid;
    end
  end

  always @(posedge ctrl_clk) begin
    if(outputArea_flow_valid) begin
      outputArea_flow_m2sPipe_payload_PRDATA <= outputArea_flow_payload_PRDATA;
      outputArea_flow_m2sPipe_payload_PSLVERROR <= outputArea_flow_payload_PSLVERROR;
    end
  end


endmodule

module EfxDMA_FlowCCUnsafeByToggle (
  input  wire          io_input_valid,
  input  wire [13:0]   io_input_payload_PADDR,
  input  wire          io_input_payload_PWRITE,
  input  wire [31:0]   io_input_payload_PWDATA,
  output wire          io_output_valid,
  output wire [13:0]   io_output_payload_PADDR,
  output wire          io_output_payload_PWRITE,
  output wire [31:0]   io_output_payload_PWDATA,
  input  wire          ctrl_clk,
  input  wire          ctrl_reset,
  input  wire          clk,
  input  wire          reset
);

  wire                inputArea_target_buffercc_io_dataOut;
  reg                 inputArea_target;
  reg        [13:0]   inputArea_data_PADDR;
  reg                 inputArea_data_PWRITE;
  reg        [31:0]   inputArea_data_PWDATA;
  wire                outputArea_target;
  reg                 outputArea_hit;
  wire                outputArea_flow_valid;
  wire       [13:0]   outputArea_flow_payload_PADDR;
  wire                outputArea_flow_payload_PWRITE;
  wire       [31:0]   outputArea_flow_payload_PWDATA;

  (* keep_hierarchy = "TRUE" *) EfxDMA_BufferCC inputArea_target_buffercc (
    .io_dataIn  (inputArea_target                    ), //i
    .io_dataOut (inputArea_target_buffercc_io_dataOut), //o
    .clk        (clk                                 ), //i
    .reset      (reset                               )  //i
  );
  assign outputArea_target = inputArea_target_buffercc_io_dataOut;
  assign outputArea_flow_valid = (outputArea_target != outputArea_hit);
  assign outputArea_flow_payload_PADDR = inputArea_data_PADDR;
  assign outputArea_flow_payload_PWRITE = inputArea_data_PWRITE;
  assign outputArea_flow_payload_PWDATA = inputArea_data_PWDATA;
  assign io_output_valid = outputArea_flow_valid;
  assign io_output_payload_PADDR = outputArea_flow_payload_PADDR;
  assign io_output_payload_PWRITE = outputArea_flow_payload_PWRITE;
  assign io_output_payload_PWDATA = outputArea_flow_payload_PWDATA;
  always @(posedge ctrl_clk) begin
    if(ctrl_reset) begin
      inputArea_target <= 1'b0;
    end else begin
      if(io_input_valid) begin
        inputArea_target <= (! inputArea_target);
      end
    end
  end

  always @(posedge ctrl_clk) begin
    if(io_input_valid) begin
      inputArea_data_PADDR <= io_input_payload_PADDR;
      inputArea_data_PWRITE <= io_input_payload_PWRITE;
      inputArea_data_PWDATA <= io_input_payload_PWDATA;
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      outputArea_hit <= 1'b0;
    end else begin
      outputArea_hit <= outputArea_target;
    end
  end


endmodule

module EfxDMA_Aggregator (
  input  wire          io_input_valid,
  output reg           io_input_ready,
  input  wire [255:0]  io_input_payload_data,
  input  wire [31:0]   io_input_payload_mask,
  output reg  [255:0]  io_output_data,
  output reg  [31:0]   io_output_mask,
  input  wire          io_output_enough,
  input  wire          io_output_consume,
  output wire          io_output_consumed,
  input  wire [4:0]    io_output_lastByteUsed,
  output wire [4:0]    io_output_usedUntil,
  input  wire          io_flush,
  input  wire [4:0]    io_offset,
  input  wire [12:0]   io_burstLength,
  input  wire          clk,
  input  wire          reset
);

  reg        [0:0]    _zz_s0_countOnesLogic_0_1;
  wire       [0:0]    _zz_s0_countOnesLogic_0_2;
  reg        [1:0]    _zz_s0_countOnesLogic_1_1;
  wire       [1:0]    _zz_s0_countOnesLogic_1_2;
  reg        [1:0]    _zz_s0_countOnesLogic_2_1;
  wire       [2:0]    _zz_s0_countOnesLogic_2_2;
  reg        [2:0]    _zz_s0_countOnesLogic_3_9;
  wire       [2:0]    _zz_s0_countOnesLogic_3_10;
  reg        [2:0]    _zz_s0_countOnesLogic_3_11;
  wire       [2:0]    _zz_s0_countOnesLogic_3_12;
  wire       [0:0]    _zz_s0_countOnesLogic_3_13;
  reg        [2:0]    _zz_s0_countOnesLogic_4_9;
  wire       [2:0]    _zz_s0_countOnesLogic_4_10;
  reg        [2:0]    _zz_s0_countOnesLogic_4_11;
  wire       [2:0]    _zz_s0_countOnesLogic_4_12;
  wire       [1:0]    _zz_s0_countOnesLogic_4_13;
  reg        [2:0]    _zz_s0_countOnesLogic_5_9;
  wire       [2:0]    _zz_s0_countOnesLogic_5_10;
  reg        [2:0]    _zz_s0_countOnesLogic_5_11;
  wire       [2:0]    _zz_s0_countOnesLogic_5_12;
  wire       [2:0]    _zz_s0_countOnesLogic_6_9;
  reg        [2:0]    _zz_s0_countOnesLogic_6_10;
  wire       [2:0]    _zz_s0_countOnesLogic_6_11;
  reg        [2:0]    _zz_s0_countOnesLogic_6_12;
  wire       [2:0]    _zz_s0_countOnesLogic_6_13;
  reg        [2:0]    _zz_s0_countOnesLogic_6_14;
  wire       [2:0]    _zz_s0_countOnesLogic_6_15;
  wire       [0:0]    _zz_s0_countOnesLogic_6_16;
  wire       [3:0]    _zz_s0_countOnesLogic_7_9;
  reg        [3:0]    _zz_s0_countOnesLogic_7_10;
  wire       [2:0]    _zz_s0_countOnesLogic_7_11;
  reg        [3:0]    _zz_s0_countOnesLogic_7_12;
  wire       [2:0]    _zz_s0_countOnesLogic_7_13;
  reg        [3:0]    _zz_s0_countOnesLogic_7_14;
  wire       [2:0]    _zz_s0_countOnesLogic_7_15;
  wire       [1:0]    _zz_s0_countOnesLogic_7_16;
  wire       [3:0]    _zz_s0_countOnesLogic_8_9;
  reg        [3:0]    _zz_s0_countOnesLogic_8_10;
  wire       [2:0]    _zz_s0_countOnesLogic_8_11;
  reg        [3:0]    _zz_s0_countOnesLogic_8_12;
  wire       [2:0]    _zz_s0_countOnesLogic_8_13;
  reg        [3:0]    _zz_s0_countOnesLogic_8_14;
  wire       [2:0]    _zz_s0_countOnesLogic_8_15;
  wire       [3:0]    _zz_s0_countOnesLogic_9_9;
  reg        [3:0]    _zz_s0_countOnesLogic_9_10;
  wire       [2:0]    _zz_s0_countOnesLogic_9_11;
  reg        [3:0]    _zz_s0_countOnesLogic_9_12;
  wire       [2:0]    _zz_s0_countOnesLogic_9_13;
  wire       [3:0]    _zz_s0_countOnesLogic_9_14;
  reg        [3:0]    _zz_s0_countOnesLogic_9_15;
  wire       [2:0]    _zz_s0_countOnesLogic_9_16;
  reg        [3:0]    _zz_s0_countOnesLogic_9_17;
  wire       [2:0]    _zz_s0_countOnesLogic_9_18;
  wire       [0:0]    _zz_s0_countOnesLogic_9_19;
  wire       [3:0]    _zz_s0_countOnesLogic_10_9;
  reg        [3:0]    _zz_s0_countOnesLogic_10_10;
  wire       [2:0]    _zz_s0_countOnesLogic_10_11;
  reg        [3:0]    _zz_s0_countOnesLogic_10_12;
  wire       [2:0]    _zz_s0_countOnesLogic_10_13;
  wire       [3:0]    _zz_s0_countOnesLogic_10_14;
  reg        [3:0]    _zz_s0_countOnesLogic_10_15;
  wire       [2:0]    _zz_s0_countOnesLogic_10_16;
  reg        [3:0]    _zz_s0_countOnesLogic_10_17;
  wire       [2:0]    _zz_s0_countOnesLogic_10_18;
  wire       [1:0]    _zz_s0_countOnesLogic_10_19;
  wire       [3:0]    _zz_s0_countOnesLogic_11_9;
  reg        [3:0]    _zz_s0_countOnesLogic_11_10;
  wire       [2:0]    _zz_s0_countOnesLogic_11_11;
  reg        [3:0]    _zz_s0_countOnesLogic_11_12;
  wire       [2:0]    _zz_s0_countOnesLogic_11_13;
  wire       [3:0]    _zz_s0_countOnesLogic_11_14;
  reg        [3:0]    _zz_s0_countOnesLogic_11_15;
  wire       [2:0]    _zz_s0_countOnesLogic_11_16;
  reg        [3:0]    _zz_s0_countOnesLogic_11_17;
  wire       [2:0]    _zz_s0_countOnesLogic_11_18;
  wire       [3:0]    _zz_s0_countOnesLogic_12_9;
  wire       [3:0]    _zz_s0_countOnesLogic_12_10;
  reg        [3:0]    _zz_s0_countOnesLogic_12_11;
  wire       [2:0]    _zz_s0_countOnesLogic_12_12;
  reg        [3:0]    _zz_s0_countOnesLogic_12_13;
  wire       [2:0]    _zz_s0_countOnesLogic_12_14;
  wire       [3:0]    _zz_s0_countOnesLogic_12_15;
  reg        [3:0]    _zz_s0_countOnesLogic_12_16;
  wire       [2:0]    _zz_s0_countOnesLogic_12_17;
  reg        [3:0]    _zz_s0_countOnesLogic_12_18;
  wire       [2:0]    _zz_s0_countOnesLogic_12_19;
  reg        [3:0]    _zz_s0_countOnesLogic_12_20;
  wire       [2:0]    _zz_s0_countOnesLogic_12_21;
  wire       [0:0]    _zz_s0_countOnesLogic_12_22;
  wire       [3:0]    _zz_s0_countOnesLogic_13_9;
  wire       [3:0]    _zz_s0_countOnesLogic_13_10;
  reg        [3:0]    _zz_s0_countOnesLogic_13_11;
  wire       [2:0]    _zz_s0_countOnesLogic_13_12;
  reg        [3:0]    _zz_s0_countOnesLogic_13_13;
  wire       [2:0]    _zz_s0_countOnesLogic_13_14;
  wire       [3:0]    _zz_s0_countOnesLogic_13_15;
  reg        [3:0]    _zz_s0_countOnesLogic_13_16;
  wire       [2:0]    _zz_s0_countOnesLogic_13_17;
  reg        [3:0]    _zz_s0_countOnesLogic_13_18;
  wire       [2:0]    _zz_s0_countOnesLogic_13_19;
  reg        [3:0]    _zz_s0_countOnesLogic_13_20;
  wire       [2:0]    _zz_s0_countOnesLogic_13_21;
  wire       [1:0]    _zz_s0_countOnesLogic_13_22;
  wire       [3:0]    _zz_s0_countOnesLogic_14_9;
  wire       [3:0]    _zz_s0_countOnesLogic_14_10;
  reg        [3:0]    _zz_s0_countOnesLogic_14_11;
  wire       [2:0]    _zz_s0_countOnesLogic_14_12;
  reg        [3:0]    _zz_s0_countOnesLogic_14_13;
  wire       [2:0]    _zz_s0_countOnesLogic_14_14;
  wire       [3:0]    _zz_s0_countOnesLogic_14_15;
  reg        [3:0]    _zz_s0_countOnesLogic_14_16;
  wire       [2:0]    _zz_s0_countOnesLogic_14_17;
  reg        [3:0]    _zz_s0_countOnesLogic_14_18;
  wire       [2:0]    _zz_s0_countOnesLogic_14_19;
  reg        [3:0]    _zz_s0_countOnesLogic_14_20;
  wire       [2:0]    _zz_s0_countOnesLogic_14_21;
  wire       [4:0]    _zz_s0_countOnesLogic_15_9;
  wire       [4:0]    _zz_s0_countOnesLogic_15_10;
  reg        [4:0]    _zz_s0_countOnesLogic_15_11;
  wire       [2:0]    _zz_s0_countOnesLogic_15_12;
  reg        [4:0]    _zz_s0_countOnesLogic_15_13;
  wire       [2:0]    _zz_s0_countOnesLogic_15_14;
  wire       [4:0]    _zz_s0_countOnesLogic_15_15;
  reg        [4:0]    _zz_s0_countOnesLogic_15_16;
  wire       [2:0]    _zz_s0_countOnesLogic_15_17;
  reg        [4:0]    _zz_s0_countOnesLogic_15_18;
  wire       [2:0]    _zz_s0_countOnesLogic_15_19;
  wire       [4:0]    _zz_s0_countOnesLogic_15_20;
  reg        [4:0]    _zz_s0_countOnesLogic_15_21;
  wire       [2:0]    _zz_s0_countOnesLogic_15_22;
  reg        [4:0]    _zz_s0_countOnesLogic_15_23;
  wire       [2:0]    _zz_s0_countOnesLogic_15_24;
  wire       [0:0]    _zz_s0_countOnesLogic_15_25;
  wire       [4:0]    _zz_s0_countOnesLogic_16_9;
  wire       [4:0]    _zz_s0_countOnesLogic_16_10;
  reg        [4:0]    _zz_s0_countOnesLogic_16_11;
  wire       [2:0]    _zz_s0_countOnesLogic_16_12;
  reg        [4:0]    _zz_s0_countOnesLogic_16_13;
  wire       [2:0]    _zz_s0_countOnesLogic_16_14;
  wire       [4:0]    _zz_s0_countOnesLogic_16_15;
  reg        [4:0]    _zz_s0_countOnesLogic_16_16;
  wire       [2:0]    _zz_s0_countOnesLogic_16_17;
  reg        [4:0]    _zz_s0_countOnesLogic_16_18;
  wire       [2:0]    _zz_s0_countOnesLogic_16_19;
  wire       [4:0]    _zz_s0_countOnesLogic_16_20;
  reg        [4:0]    _zz_s0_countOnesLogic_16_21;
  wire       [2:0]    _zz_s0_countOnesLogic_16_22;
  reg        [4:0]    _zz_s0_countOnesLogic_16_23;
  wire       [2:0]    _zz_s0_countOnesLogic_16_24;
  wire       [1:0]    _zz_s0_countOnesLogic_16_25;
  wire       [4:0]    _zz_s0_countOnesLogic_17_9;
  wire       [4:0]    _zz_s0_countOnesLogic_17_10;
  reg        [4:0]    _zz_s0_countOnesLogic_17_11;
  wire       [2:0]    _zz_s0_countOnesLogic_17_12;
  reg        [4:0]    _zz_s0_countOnesLogic_17_13;
  wire       [2:0]    _zz_s0_countOnesLogic_17_14;
  wire       [4:0]    _zz_s0_countOnesLogic_17_15;
  reg        [4:0]    _zz_s0_countOnesLogic_17_16;
  wire       [2:0]    _zz_s0_countOnesLogic_17_17;
  reg        [4:0]    _zz_s0_countOnesLogic_17_18;
  wire       [2:0]    _zz_s0_countOnesLogic_17_19;
  wire       [4:0]    _zz_s0_countOnesLogic_17_20;
  reg        [4:0]    _zz_s0_countOnesLogic_17_21;
  wire       [2:0]    _zz_s0_countOnesLogic_17_22;
  reg        [4:0]    _zz_s0_countOnesLogic_17_23;
  wire       [2:0]    _zz_s0_countOnesLogic_17_24;
  wire       [4:0]    _zz_s0_countOnesLogic_18_9;
  wire       [4:0]    _zz_s0_countOnesLogic_18_10;
  reg        [4:0]    _zz_s0_countOnesLogic_18_11;
  wire       [2:0]    _zz_s0_countOnesLogic_18_12;
  reg        [4:0]    _zz_s0_countOnesLogic_18_13;
  wire       [2:0]    _zz_s0_countOnesLogic_18_14;
  wire       [4:0]    _zz_s0_countOnesLogic_18_15;
  reg        [4:0]    _zz_s0_countOnesLogic_18_16;
  wire       [2:0]    _zz_s0_countOnesLogic_18_17;
  reg        [4:0]    _zz_s0_countOnesLogic_18_18;
  wire       [2:0]    _zz_s0_countOnesLogic_18_19;
  wire       [4:0]    _zz_s0_countOnesLogic_18_20;
  wire       [4:0]    _zz_s0_countOnesLogic_18_21;
  reg        [4:0]    _zz_s0_countOnesLogic_18_22;
  wire       [2:0]    _zz_s0_countOnesLogic_18_23;
  reg        [4:0]    _zz_s0_countOnesLogic_18_24;
  wire       [2:0]    _zz_s0_countOnesLogic_18_25;
  reg        [4:0]    _zz_s0_countOnesLogic_18_26;
  wire       [2:0]    _zz_s0_countOnesLogic_18_27;
  wire       [0:0]    _zz_s0_countOnesLogic_18_28;
  wire       [4:0]    _zz_s0_countOnesLogic_19_9;
  wire       [4:0]    _zz_s0_countOnesLogic_19_10;
  reg        [4:0]    _zz_s0_countOnesLogic_19_11;
  wire       [2:0]    _zz_s0_countOnesLogic_19_12;
  reg        [4:0]    _zz_s0_countOnesLogic_19_13;
  wire       [2:0]    _zz_s0_countOnesLogic_19_14;
  wire       [4:0]    _zz_s0_countOnesLogic_19_15;
  reg        [4:0]    _zz_s0_countOnesLogic_19_16;
  wire       [2:0]    _zz_s0_countOnesLogic_19_17;
  reg        [4:0]    _zz_s0_countOnesLogic_19_18;
  wire       [2:0]    _zz_s0_countOnesLogic_19_19;
  wire       [4:0]    _zz_s0_countOnesLogic_19_20;
  wire       [4:0]    _zz_s0_countOnesLogic_19_21;
  reg        [4:0]    _zz_s0_countOnesLogic_19_22;
  wire       [2:0]    _zz_s0_countOnesLogic_19_23;
  reg        [4:0]    _zz_s0_countOnesLogic_19_24;
  wire       [2:0]    _zz_s0_countOnesLogic_19_25;
  reg        [4:0]    _zz_s0_countOnesLogic_19_26;
  wire       [2:0]    _zz_s0_countOnesLogic_19_27;
  wire       [1:0]    _zz_s0_countOnesLogic_19_28;
  wire       [4:0]    _zz_s0_countOnesLogic_20_9;
  wire       [4:0]    _zz_s0_countOnesLogic_20_10;
  reg        [4:0]    _zz_s0_countOnesLogic_20_11;
  wire       [2:0]    _zz_s0_countOnesLogic_20_12;
  reg        [4:0]    _zz_s0_countOnesLogic_20_13;
  wire       [2:0]    _zz_s0_countOnesLogic_20_14;
  wire       [4:0]    _zz_s0_countOnesLogic_20_15;
  reg        [4:0]    _zz_s0_countOnesLogic_20_16;
  wire       [2:0]    _zz_s0_countOnesLogic_20_17;
  reg        [4:0]    _zz_s0_countOnesLogic_20_18;
  wire       [2:0]    _zz_s0_countOnesLogic_20_19;
  wire       [4:0]    _zz_s0_countOnesLogic_20_20;
  wire       [4:0]    _zz_s0_countOnesLogic_20_21;
  reg        [4:0]    _zz_s0_countOnesLogic_20_22;
  wire       [2:0]    _zz_s0_countOnesLogic_20_23;
  reg        [4:0]    _zz_s0_countOnesLogic_20_24;
  wire       [2:0]    _zz_s0_countOnesLogic_20_25;
  reg        [4:0]    _zz_s0_countOnesLogic_20_26;
  wire       [2:0]    _zz_s0_countOnesLogic_20_27;
  wire       [4:0]    _zz_s0_countOnesLogic_21_9;
  wire       [4:0]    _zz_s0_countOnesLogic_21_10;
  reg        [4:0]    _zz_s0_countOnesLogic_21_11;
  wire       [2:0]    _zz_s0_countOnesLogic_21_12;
  reg        [4:0]    _zz_s0_countOnesLogic_21_13;
  wire       [2:0]    _zz_s0_countOnesLogic_21_14;
  wire       [4:0]    _zz_s0_countOnesLogic_21_15;
  reg        [4:0]    _zz_s0_countOnesLogic_21_16;
  wire       [2:0]    _zz_s0_countOnesLogic_21_17;
  reg        [4:0]    _zz_s0_countOnesLogic_21_18;
  wire       [2:0]    _zz_s0_countOnesLogic_21_19;
  wire       [4:0]    _zz_s0_countOnesLogic_21_20;
  wire       [4:0]    _zz_s0_countOnesLogic_21_21;
  reg        [4:0]    _zz_s0_countOnesLogic_21_22;
  wire       [2:0]    _zz_s0_countOnesLogic_21_23;
  reg        [4:0]    _zz_s0_countOnesLogic_21_24;
  wire       [2:0]    _zz_s0_countOnesLogic_21_25;
  wire       [4:0]    _zz_s0_countOnesLogic_21_26;
  reg        [4:0]    _zz_s0_countOnesLogic_21_27;
  wire       [2:0]    _zz_s0_countOnesLogic_21_28;
  reg        [4:0]    _zz_s0_countOnesLogic_21_29;
  wire       [2:0]    _zz_s0_countOnesLogic_21_30;
  wire       [0:0]    _zz_s0_countOnesLogic_21_31;
  wire       [4:0]    _zz_s0_countOnesLogic_22_9;
  wire       [4:0]    _zz_s0_countOnesLogic_22_10;
  reg        [4:0]    _zz_s0_countOnesLogic_22_11;
  wire       [2:0]    _zz_s0_countOnesLogic_22_12;
  reg        [4:0]    _zz_s0_countOnesLogic_22_13;
  wire       [2:0]    _zz_s0_countOnesLogic_22_14;
  wire       [4:0]    _zz_s0_countOnesLogic_22_15;
  reg        [4:0]    _zz_s0_countOnesLogic_22_16;
  wire       [2:0]    _zz_s0_countOnesLogic_22_17;
  reg        [4:0]    _zz_s0_countOnesLogic_22_18;
  wire       [2:0]    _zz_s0_countOnesLogic_22_19;
  wire       [4:0]    _zz_s0_countOnesLogic_22_20;
  wire       [4:0]    _zz_s0_countOnesLogic_22_21;
  reg        [4:0]    _zz_s0_countOnesLogic_22_22;
  wire       [2:0]    _zz_s0_countOnesLogic_22_23;
  reg        [4:0]    _zz_s0_countOnesLogic_22_24;
  wire       [2:0]    _zz_s0_countOnesLogic_22_25;
  wire       [4:0]    _zz_s0_countOnesLogic_22_26;
  reg        [4:0]    _zz_s0_countOnesLogic_22_27;
  wire       [2:0]    _zz_s0_countOnesLogic_22_28;
  reg        [4:0]    _zz_s0_countOnesLogic_22_29;
  wire       [2:0]    _zz_s0_countOnesLogic_22_30;
  wire       [1:0]    _zz_s0_countOnesLogic_22_31;
  wire       [4:0]    _zz_s0_countOnesLogic_23_9;
  wire       [4:0]    _zz_s0_countOnesLogic_23_10;
  reg        [4:0]    _zz_s0_countOnesLogic_23_11;
  wire       [2:0]    _zz_s0_countOnesLogic_23_12;
  reg        [4:0]    _zz_s0_countOnesLogic_23_13;
  wire       [2:0]    _zz_s0_countOnesLogic_23_14;
  wire       [4:0]    _zz_s0_countOnesLogic_23_15;
  reg        [4:0]    _zz_s0_countOnesLogic_23_16;
  wire       [2:0]    _zz_s0_countOnesLogic_23_17;
  reg        [4:0]    _zz_s0_countOnesLogic_23_18;
  wire       [2:0]    _zz_s0_countOnesLogic_23_19;
  wire       [4:0]    _zz_s0_countOnesLogic_23_20;
  wire       [4:0]    _zz_s0_countOnesLogic_23_21;
  reg        [4:0]    _zz_s0_countOnesLogic_23_22;
  wire       [2:0]    _zz_s0_countOnesLogic_23_23;
  reg        [4:0]    _zz_s0_countOnesLogic_23_24;
  wire       [2:0]    _zz_s0_countOnesLogic_23_25;
  wire       [4:0]    _zz_s0_countOnesLogic_23_26;
  reg        [4:0]    _zz_s0_countOnesLogic_23_27;
  wire       [2:0]    _zz_s0_countOnesLogic_23_28;
  reg        [4:0]    _zz_s0_countOnesLogic_23_29;
  wire       [2:0]    _zz_s0_countOnesLogic_23_30;
  wire       [4:0]    _zz_s0_countOnesLogic_24_9;
  wire       [4:0]    _zz_s0_countOnesLogic_24_10;
  wire       [4:0]    _zz_s0_countOnesLogic_24_11;
  reg        [4:0]    _zz_s0_countOnesLogic_24_12;
  wire       [2:0]    _zz_s0_countOnesLogic_24_13;
  reg        [4:0]    _zz_s0_countOnesLogic_24_14;
  wire       [2:0]    _zz_s0_countOnesLogic_24_15;
  wire       [4:0]    _zz_s0_countOnesLogic_24_16;
  reg        [4:0]    _zz_s0_countOnesLogic_24_17;
  wire       [2:0]    _zz_s0_countOnesLogic_24_18;
  reg        [4:0]    _zz_s0_countOnesLogic_24_19;
  wire       [2:0]    _zz_s0_countOnesLogic_24_20;
  wire       [4:0]    _zz_s0_countOnesLogic_24_21;
  wire       [4:0]    _zz_s0_countOnesLogic_24_22;
  reg        [4:0]    _zz_s0_countOnesLogic_24_23;
  wire       [2:0]    _zz_s0_countOnesLogic_24_24;
  reg        [4:0]    _zz_s0_countOnesLogic_24_25;
  wire       [2:0]    _zz_s0_countOnesLogic_24_26;
  wire       [4:0]    _zz_s0_countOnesLogic_24_27;
  reg        [4:0]    _zz_s0_countOnesLogic_24_28;
  wire       [2:0]    _zz_s0_countOnesLogic_24_29;
  reg        [4:0]    _zz_s0_countOnesLogic_24_30;
  wire       [2:0]    _zz_s0_countOnesLogic_24_31;
  reg        [4:0]    _zz_s0_countOnesLogic_24_32;
  wire       [2:0]    _zz_s0_countOnesLogic_24_33;
  wire       [0:0]    _zz_s0_countOnesLogic_24_34;
  wire       [4:0]    _zz_s0_countOnesLogic_25_9;
  wire       [4:0]    _zz_s0_countOnesLogic_25_10;
  wire       [4:0]    _zz_s0_countOnesLogic_25_11;
  reg        [4:0]    _zz_s0_countOnesLogic_25_12;
  wire       [2:0]    _zz_s0_countOnesLogic_25_13;
  reg        [4:0]    _zz_s0_countOnesLogic_25_14;
  wire       [2:0]    _zz_s0_countOnesLogic_25_15;
  wire       [4:0]    _zz_s0_countOnesLogic_25_16;
  reg        [4:0]    _zz_s0_countOnesLogic_25_17;
  wire       [2:0]    _zz_s0_countOnesLogic_25_18;
  reg        [4:0]    _zz_s0_countOnesLogic_25_19;
  wire       [2:0]    _zz_s0_countOnesLogic_25_20;
  wire       [4:0]    _zz_s0_countOnesLogic_25_21;
  wire       [4:0]    _zz_s0_countOnesLogic_25_22;
  reg        [4:0]    _zz_s0_countOnesLogic_25_23;
  wire       [2:0]    _zz_s0_countOnesLogic_25_24;
  reg        [4:0]    _zz_s0_countOnesLogic_25_25;
  wire       [2:0]    _zz_s0_countOnesLogic_25_26;
  wire       [4:0]    _zz_s0_countOnesLogic_25_27;
  reg        [4:0]    _zz_s0_countOnesLogic_25_28;
  wire       [2:0]    _zz_s0_countOnesLogic_25_29;
  reg        [4:0]    _zz_s0_countOnesLogic_25_30;
  wire       [2:0]    _zz_s0_countOnesLogic_25_31;
  reg        [4:0]    _zz_s0_countOnesLogic_25_32;
  wire       [2:0]    _zz_s0_countOnesLogic_25_33;
  wire       [1:0]    _zz_s0_countOnesLogic_25_34;
  wire       [4:0]    _zz_s0_countOnesLogic_26_9;
  wire       [4:0]    _zz_s0_countOnesLogic_26_10;
  wire       [4:0]    _zz_s0_countOnesLogic_26_11;
  reg        [4:0]    _zz_s0_countOnesLogic_26_12;
  wire       [2:0]    _zz_s0_countOnesLogic_26_13;
  reg        [4:0]    _zz_s0_countOnesLogic_26_14;
  wire       [2:0]    _zz_s0_countOnesLogic_26_15;
  wire       [4:0]    _zz_s0_countOnesLogic_26_16;
  reg        [4:0]    _zz_s0_countOnesLogic_26_17;
  wire       [2:0]    _zz_s0_countOnesLogic_26_18;
  reg        [4:0]    _zz_s0_countOnesLogic_26_19;
  wire       [2:0]    _zz_s0_countOnesLogic_26_20;
  wire       [4:0]    _zz_s0_countOnesLogic_26_21;
  wire       [4:0]    _zz_s0_countOnesLogic_26_22;
  reg        [4:0]    _zz_s0_countOnesLogic_26_23;
  wire       [2:0]    _zz_s0_countOnesLogic_26_24;
  reg        [4:0]    _zz_s0_countOnesLogic_26_25;
  wire       [2:0]    _zz_s0_countOnesLogic_26_26;
  wire       [4:0]    _zz_s0_countOnesLogic_26_27;
  reg        [4:0]    _zz_s0_countOnesLogic_26_28;
  wire       [2:0]    _zz_s0_countOnesLogic_26_29;
  reg        [4:0]    _zz_s0_countOnesLogic_26_30;
  wire       [2:0]    _zz_s0_countOnesLogic_26_31;
  reg        [4:0]    _zz_s0_countOnesLogic_26_32;
  wire       [2:0]    _zz_s0_countOnesLogic_26_33;
  wire       [4:0]    _zz_s0_countOnesLogic_27_9;
  wire       [4:0]    _zz_s0_countOnesLogic_27_10;
  wire       [4:0]    _zz_s0_countOnesLogic_27_11;
  reg        [4:0]    _zz_s0_countOnesLogic_27_12;
  wire       [2:0]    _zz_s0_countOnesLogic_27_13;
  reg        [4:0]    _zz_s0_countOnesLogic_27_14;
  wire       [2:0]    _zz_s0_countOnesLogic_27_15;
  wire       [4:0]    _zz_s0_countOnesLogic_27_16;
  reg        [4:0]    _zz_s0_countOnesLogic_27_17;
  wire       [2:0]    _zz_s0_countOnesLogic_27_18;
  reg        [4:0]    _zz_s0_countOnesLogic_27_19;
  wire       [2:0]    _zz_s0_countOnesLogic_27_20;
  wire       [4:0]    _zz_s0_countOnesLogic_27_21;
  wire       [4:0]    _zz_s0_countOnesLogic_27_22;
  reg        [4:0]    _zz_s0_countOnesLogic_27_23;
  wire       [2:0]    _zz_s0_countOnesLogic_27_24;
  reg        [4:0]    _zz_s0_countOnesLogic_27_25;
  wire       [2:0]    _zz_s0_countOnesLogic_27_26;
  wire       [4:0]    _zz_s0_countOnesLogic_27_27;
  reg        [4:0]    _zz_s0_countOnesLogic_27_28;
  wire       [2:0]    _zz_s0_countOnesLogic_27_29;
  reg        [4:0]    _zz_s0_countOnesLogic_27_30;
  wire       [2:0]    _zz_s0_countOnesLogic_27_31;
  wire       [4:0]    _zz_s0_countOnesLogic_27_32;
  reg        [4:0]    _zz_s0_countOnesLogic_27_33;
  wire       [2:0]    _zz_s0_countOnesLogic_27_34;
  reg        [4:0]    _zz_s0_countOnesLogic_27_35;
  wire       [2:0]    _zz_s0_countOnesLogic_27_36;
  wire       [0:0]    _zz_s0_countOnesLogic_27_37;
  wire       [4:0]    _zz_s0_countOnesLogic_28_9;
  wire       [4:0]    _zz_s0_countOnesLogic_28_10;
  wire       [4:0]    _zz_s0_countOnesLogic_28_11;
  reg        [4:0]    _zz_s0_countOnesLogic_28_12;
  wire       [2:0]    _zz_s0_countOnesLogic_28_13;
  reg        [4:0]    _zz_s0_countOnesLogic_28_14;
  wire       [2:0]    _zz_s0_countOnesLogic_28_15;
  wire       [4:0]    _zz_s0_countOnesLogic_28_16;
  reg        [4:0]    _zz_s0_countOnesLogic_28_17;
  wire       [2:0]    _zz_s0_countOnesLogic_28_18;
  reg        [4:0]    _zz_s0_countOnesLogic_28_19;
  wire       [2:0]    _zz_s0_countOnesLogic_28_20;
  wire       [4:0]    _zz_s0_countOnesLogic_28_21;
  wire       [4:0]    _zz_s0_countOnesLogic_28_22;
  reg        [4:0]    _zz_s0_countOnesLogic_28_23;
  wire       [2:0]    _zz_s0_countOnesLogic_28_24;
  reg        [4:0]    _zz_s0_countOnesLogic_28_25;
  wire       [2:0]    _zz_s0_countOnesLogic_28_26;
  wire       [4:0]    _zz_s0_countOnesLogic_28_27;
  reg        [4:0]    _zz_s0_countOnesLogic_28_28;
  wire       [2:0]    _zz_s0_countOnesLogic_28_29;
  reg        [4:0]    _zz_s0_countOnesLogic_28_30;
  wire       [2:0]    _zz_s0_countOnesLogic_28_31;
  wire       [4:0]    _zz_s0_countOnesLogic_28_32;
  reg        [4:0]    _zz_s0_countOnesLogic_28_33;
  wire       [2:0]    _zz_s0_countOnesLogic_28_34;
  reg        [4:0]    _zz_s0_countOnesLogic_28_35;
  wire       [2:0]    _zz_s0_countOnesLogic_28_36;
  wire       [1:0]    _zz_s0_countOnesLogic_28_37;
  wire       [4:0]    _zz_s0_countOnesLogic_29_9;
  wire       [4:0]    _zz_s0_countOnesLogic_29_10;
  wire       [4:0]    _zz_s0_countOnesLogic_29_11;
  reg        [4:0]    _zz_s0_countOnesLogic_29_12;
  wire       [2:0]    _zz_s0_countOnesLogic_29_13;
  reg        [4:0]    _zz_s0_countOnesLogic_29_14;
  wire       [2:0]    _zz_s0_countOnesLogic_29_15;
  wire       [4:0]    _zz_s0_countOnesLogic_29_16;
  reg        [4:0]    _zz_s0_countOnesLogic_29_17;
  wire       [2:0]    _zz_s0_countOnesLogic_29_18;
  reg        [4:0]    _zz_s0_countOnesLogic_29_19;
  wire       [2:0]    _zz_s0_countOnesLogic_29_20;
  wire       [4:0]    _zz_s0_countOnesLogic_29_21;
  wire       [4:0]    _zz_s0_countOnesLogic_29_22;
  reg        [4:0]    _zz_s0_countOnesLogic_29_23;
  wire       [2:0]    _zz_s0_countOnesLogic_29_24;
  reg        [4:0]    _zz_s0_countOnesLogic_29_25;
  wire       [2:0]    _zz_s0_countOnesLogic_29_26;
  wire       [4:0]    _zz_s0_countOnesLogic_29_27;
  reg        [4:0]    _zz_s0_countOnesLogic_29_28;
  wire       [2:0]    _zz_s0_countOnesLogic_29_29;
  reg        [4:0]    _zz_s0_countOnesLogic_29_30;
  wire       [2:0]    _zz_s0_countOnesLogic_29_31;
  wire       [4:0]    _zz_s0_countOnesLogic_29_32;
  reg        [4:0]    _zz_s0_countOnesLogic_29_33;
  wire       [2:0]    _zz_s0_countOnesLogic_29_34;
  reg        [4:0]    _zz_s0_countOnesLogic_29_35;
  wire       [2:0]    _zz_s0_countOnesLogic_29_36;
  wire       [4:0]    _zz_s0_countOnesLogic_30_9;
  wire       [4:0]    _zz_s0_countOnesLogic_30_10;
  wire       [4:0]    _zz_s0_countOnesLogic_30_11;
  reg        [4:0]    _zz_s0_countOnesLogic_30_12;
  wire       [2:0]    _zz_s0_countOnesLogic_30_13;
  reg        [4:0]    _zz_s0_countOnesLogic_30_14;
  wire       [2:0]    _zz_s0_countOnesLogic_30_15;
  wire       [4:0]    _zz_s0_countOnesLogic_30_16;
  reg        [4:0]    _zz_s0_countOnesLogic_30_17;
  wire       [2:0]    _zz_s0_countOnesLogic_30_18;
  reg        [4:0]    _zz_s0_countOnesLogic_30_19;
  wire       [2:0]    _zz_s0_countOnesLogic_30_20;
  wire       [4:0]    _zz_s0_countOnesLogic_30_21;
  wire       [4:0]    _zz_s0_countOnesLogic_30_22;
  reg        [4:0]    _zz_s0_countOnesLogic_30_23;
  wire       [2:0]    _zz_s0_countOnesLogic_30_24;
  reg        [4:0]    _zz_s0_countOnesLogic_30_25;
  wire       [2:0]    _zz_s0_countOnesLogic_30_26;
  wire       [4:0]    _zz_s0_countOnesLogic_30_27;
  reg        [4:0]    _zz_s0_countOnesLogic_30_28;
  wire       [2:0]    _zz_s0_countOnesLogic_30_29;
  reg        [4:0]    _zz_s0_countOnesLogic_30_30;
  wire       [2:0]    _zz_s0_countOnesLogic_30_31;
  wire       [4:0]    _zz_s0_countOnesLogic_30_32;
  wire       [4:0]    _zz_s0_countOnesLogic_30_33;
  reg        [4:0]    _zz_s0_countOnesLogic_30_34;
  wire       [2:0]    _zz_s0_countOnesLogic_30_35;
  reg        [4:0]    _zz_s0_countOnesLogic_30_36;
  wire       [2:0]    _zz_s0_countOnesLogic_30_37;
  reg        [4:0]    _zz_s0_countOnesLogic_30_38;
  wire       [2:0]    _zz_s0_countOnesLogic_30_39;
  wire       [0:0]    _zz_s0_countOnesLogic_30_40;
  wire       [5:0]    _zz_s0_countOnesLogic_31_8;
  wire       [5:0]    _zz_s0_countOnesLogic_31_9;
  wire       [5:0]    _zz_s0_countOnesLogic_31_10;
  reg        [5:0]    _zz_s0_countOnesLogic_31_11;
  wire       [2:0]    _zz_s0_countOnesLogic_31_12;
  reg        [5:0]    _zz_s0_countOnesLogic_31_13;
  wire       [2:0]    _zz_s0_countOnesLogic_31_14;
  wire       [5:0]    _zz_s0_countOnesLogic_31_15;
  reg        [5:0]    _zz_s0_countOnesLogic_31_16;
  wire       [2:0]    _zz_s0_countOnesLogic_31_17;
  reg        [5:0]    _zz_s0_countOnesLogic_31_18;
  wire       [2:0]    _zz_s0_countOnesLogic_31_19;
  wire       [5:0]    _zz_s0_countOnesLogic_31_20;
  wire       [5:0]    _zz_s0_countOnesLogic_31_21;
  reg        [5:0]    _zz_s0_countOnesLogic_31_22;
  wire       [2:0]    _zz_s0_countOnesLogic_31_23;
  reg        [5:0]    _zz_s0_countOnesLogic_31_24;
  wire       [2:0]    _zz_s0_countOnesLogic_31_25;
  wire       [5:0]    _zz_s0_countOnesLogic_31_26;
  reg        [5:0]    _zz_s0_countOnesLogic_31_27;
  wire       [2:0]    _zz_s0_countOnesLogic_31_28;
  reg        [5:0]    _zz_s0_countOnesLogic_31_29;
  wire       [2:0]    _zz_s0_countOnesLogic_31_30;
  wire       [5:0]    _zz_s0_countOnesLogic_31_31;
  wire       [5:0]    _zz_s0_countOnesLogic_31_32;
  reg        [5:0]    _zz_s0_countOnesLogic_31_33;
  wire       [2:0]    _zz_s0_countOnesLogic_31_34;
  reg        [5:0]    _zz_s0_countOnesLogic_31_35;
  wire       [2:0]    _zz_s0_countOnesLogic_31_36;
  reg        [5:0]    _zz_s0_countOnesLogic_31_37;
  wire       [2:0]    _zz_s0_countOnesLogic_31_38;
  wire       [1:0]    _zz_s0_countOnesLogic_31_39;
  wire       [5:0]    _zz_s1_offsetNext;
  wire       [13:0]   _zz_s1_byteCounter;
  wire       [4:0]    _zz_s1_inputIndexes_1;
  wire       [4:0]    _zz_s1_inputIndexes_2;
  wire       [4:0]    _zz_s1_inputIndexes_3;
  wire       [4:0]    _zz_s1_inputIndexes_4;
  wire       [4:0]    _zz_s1_inputIndexes_5;
  wire       [4:0]    _zz_s1_inputIndexes_6;
  wire       [4:0]    _zz_s1_inputIndexes_7;
  wire       [4:0]    _zz_s1_inputIndexes_8;
  wire       [4:0]    _zz_s1_inputIndexes_9;
  wire       [4:0]    _zz_s1_inputIndexes_10;
  wire       [4:0]    _zz_s1_inputIndexes_11;
  wire       [4:0]    _zz_s1_inputIndexes_12;
  wire       [4:0]    _zz_s1_inputIndexes_13;
  wire       [4:0]    _zz_s1_inputIndexes_14;
  wire       [4:0]    _zz_s1_inputIndexes_15;
  wire       [0:0]    _zz_s1_outputPayload_selValid_992;
  wire       [22:0]   _zz_s1_outputPayload_selValid_993;
  wire       [0:0]    _zz_s1_outputPayload_selValid_994;
  wire       [11:0]   _zz_s1_outputPayload_selValid_995;
  wire       [0:0]    _zz_s1_outputPayload_selValid_996;
  wire       [0:0]    _zz_s1_outputPayload_selValid_997;
  wire       [0:0]    _zz_s1_outputPayload_selValid_998;
  wire       [22:0]   _zz_s1_outputPayload_selValid_999;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1000;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1001;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1002;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1003;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1004;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1005;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1006;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1007;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1008;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1009;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1010;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1011;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1012;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1013;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1014;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1015;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1016;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1017;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1018;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1019;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1020;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1021;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1022;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1023;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1024;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1025;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1026;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1027;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1028;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1029;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1030;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1031;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1032;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1033;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1034;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1035;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1036;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1037;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1038;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1039;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1040;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1041;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1042;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1043;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1044;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1045;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1046;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1047;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1048;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1049;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1050;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1051;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1052;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1053;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1054;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1055;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1056;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1057;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1058;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1059;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1060;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1061;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1062;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1063;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1064;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1065;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1066;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1067;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1068;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1069;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1070;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1071;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1072;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1073;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1074;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1075;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1076;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1077;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1078;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1079;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1080;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1081;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1082;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1083;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1084;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1085;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1086;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1087;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1088;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1089;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1090;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1091;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1092;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1093;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1094;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1095;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1096;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1097;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1098;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1099;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1100;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1101;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1102;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1103;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1104;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1105;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1106;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1107;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1108;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1109;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1110;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1111;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1112;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1113;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1114;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1115;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1116;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1117;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1118;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1119;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1120;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1121;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1122;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1123;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1124;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1125;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1126;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1127;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1128;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1129;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1130;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1131;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1132;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1133;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1134;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1135;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1136;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1137;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1138;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1139;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1140;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1141;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1142;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1143;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1144;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1145;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1146;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1147;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1148;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1149;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1150;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1151;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1152;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1153;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1154;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1155;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1156;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1157;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1158;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1159;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1160;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1161;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1162;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1163;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1164;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1165;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1166;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1167;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1168;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1169;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1170;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1171;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1172;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1173;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1174;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1175;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1176;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1177;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1178;
  wire       [22:0]   _zz_s1_outputPayload_selValid_1179;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1180;
  wire       [11:0]   _zz_s1_outputPayload_selValid_1181;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1182;
  wire       [0:0]    _zz_s1_outputPayload_selValid_1183;
  wire       [13:0]   _zz_when_DmaSg_l1464;
  reg        [7:0]    _zz_s2_byteLogic_0_inputData;
  reg        [7:0]    _zz_s2_byteLogic_1_inputData;
  reg        [7:0]    _zz_s2_byteLogic_2_inputData;
  reg        [7:0]    _zz_s2_byteLogic_3_inputData;
  reg        [7:0]    _zz_s2_byteLogic_4_inputData;
  reg        [7:0]    _zz_s2_byteLogic_5_inputData;
  reg        [7:0]    _zz_s2_byteLogic_6_inputData;
  reg        [7:0]    _zz_s2_byteLogic_7_inputData;
  reg        [7:0]    _zz_s2_byteLogic_8_inputData;
  reg        [7:0]    _zz_s2_byteLogic_9_inputData;
  reg        [7:0]    _zz_s2_byteLogic_10_inputData;
  reg        [7:0]    _zz_s2_byteLogic_11_inputData;
  reg        [7:0]    _zz_s2_byteLogic_12_inputData;
  reg        [7:0]    _zz_s2_byteLogic_13_inputData;
  reg        [7:0]    _zz_s2_byteLogic_14_inputData;
  reg        [7:0]    _zz_s2_byteLogic_15_inputData;
  reg        [7:0]    _zz_s2_byteLogic_16_inputData;
  reg        [7:0]    _zz_s2_byteLogic_17_inputData;
  reg        [7:0]    _zz_s2_byteLogic_18_inputData;
  reg        [7:0]    _zz_s2_byteLogic_19_inputData;
  reg        [7:0]    _zz_s2_byteLogic_20_inputData;
  reg        [7:0]    _zz_s2_byteLogic_21_inputData;
  reg        [7:0]    _zz_s2_byteLogic_22_inputData;
  reg        [7:0]    _zz_s2_byteLogic_23_inputData;
  reg        [7:0]    _zz_s2_byteLogic_24_inputData;
  reg        [7:0]    _zz_s2_byteLogic_25_inputData;
  reg        [7:0]    _zz_s2_byteLogic_26_inputData;
  reg        [7:0]    _zz_s2_byteLogic_27_inputData;
  reg        [7:0]    _zz_s2_byteLogic_28_inputData;
  reg        [7:0]    _zz_s2_byteLogic_29_inputData;
  reg        [7:0]    _zz_s2_byteLogic_30_inputData;
  reg        [7:0]    _zz_s2_byteLogic_31_inputData;
  reg        [4:0]    _zz_io_output_usedUntil_5;
  wire       [4:0]    _zz_io_output_usedUntil_6;
  wire                s0_input_valid;
  wire                s0_input_ready;
  wire       [255:0]  s0_input_payload_data;
  wire       [31:0]   s0_input_payload_mask;
  reg                 io_input_rValid;
  reg        [255:0]  io_input_rData_data;
  reg        [31:0]   io_input_rData_mask;
  wire                when_Stream_l375;
  wire                _zz_s0_countOnesLogic_0;
  wire                _zz_s0_countOnesLogic_1;
  wire                _zz_s0_countOnesLogic_2;
  wire                _zz_s0_countOnesLogic_3;
  wire                _zz_s0_countOnesLogic_4;
  wire                _zz_s0_countOnesLogic_5;
  wire                _zz_s0_countOnesLogic_6;
  wire                _zz_s0_countOnesLogic_7;
  wire                _zz_s0_countOnesLogic_8;
  wire                _zz_s0_countOnesLogic_9;
  wire                _zz_s0_countOnesLogic_10;
  wire                _zz_s0_countOnesLogic_11;
  wire                _zz_s0_countOnesLogic_12;
  wire                _zz_s0_countOnesLogic_13;
  wire                _zz_s0_countOnesLogic_14;
  wire                _zz_s0_countOnesLogic_15;
  wire                _zz_s0_countOnesLogic_16;
  wire                _zz_s0_countOnesLogic_17;
  wire                _zz_s0_countOnesLogic_18;
  wire                _zz_s0_countOnesLogic_19;
  wire                _zz_s0_countOnesLogic_20;
  wire                _zz_s0_countOnesLogic_21;
  wire                _zz_s0_countOnesLogic_22;
  wire                _zz_s0_countOnesLogic_23;
  wire                _zz_s0_countOnesLogic_24;
  wire                _zz_s0_countOnesLogic_25;
  wire                _zz_s0_countOnesLogic_26;
  wire                _zz_s0_countOnesLogic_27;
  wire                _zz_s0_countOnesLogic_28;
  wire                _zz_s0_countOnesLogic_29;
  wire                _zz_s0_countOnesLogic_30;
  wire       [0:0]    s0_countOnesLogic_0;
  wire       [1:0]    s0_countOnesLogic_1;
  wire       [1:0]    s0_countOnesLogic_2;
  wire       [2:0]    _zz_s0_countOnesLogic_3_1;
  wire       [2:0]    _zz_s0_countOnesLogic_3_2;
  wire       [2:0]    _zz_s0_countOnesLogic_3_3;
  wire       [2:0]    _zz_s0_countOnesLogic_3_4;
  wire       [2:0]    _zz_s0_countOnesLogic_3_5;
  wire       [2:0]    _zz_s0_countOnesLogic_3_6;
  wire       [2:0]    _zz_s0_countOnesLogic_3_7;
  wire       [2:0]    _zz_s0_countOnesLogic_3_8;
  wire       [2:0]    s0_countOnesLogic_3;
  wire       [2:0]    _zz_s0_countOnesLogic_4_1;
  wire       [2:0]    _zz_s0_countOnesLogic_4_2;
  wire       [2:0]    _zz_s0_countOnesLogic_4_3;
  wire       [2:0]    _zz_s0_countOnesLogic_4_4;
  wire       [2:0]    _zz_s0_countOnesLogic_4_5;
  wire       [2:0]    _zz_s0_countOnesLogic_4_6;
  wire       [2:0]    _zz_s0_countOnesLogic_4_7;
  wire       [2:0]    _zz_s0_countOnesLogic_4_8;
  wire       [2:0]    s0_countOnesLogic_4;
  wire       [2:0]    _zz_s0_countOnesLogic_5_1;
  wire       [2:0]    _zz_s0_countOnesLogic_5_2;
  wire       [2:0]    _zz_s0_countOnesLogic_5_3;
  wire       [2:0]    _zz_s0_countOnesLogic_5_4;
  wire       [2:0]    _zz_s0_countOnesLogic_5_5;
  wire       [2:0]    _zz_s0_countOnesLogic_5_6;
  wire       [2:0]    _zz_s0_countOnesLogic_5_7;
  wire       [2:0]    _zz_s0_countOnesLogic_5_8;
  wire       [2:0]    s0_countOnesLogic_5;
  wire       [2:0]    _zz_s0_countOnesLogic_6_1;
  wire       [2:0]    _zz_s0_countOnesLogic_6_2;
  wire       [2:0]    _zz_s0_countOnesLogic_6_3;
  wire       [2:0]    _zz_s0_countOnesLogic_6_4;
  wire       [2:0]    _zz_s0_countOnesLogic_6_5;
  wire       [2:0]    _zz_s0_countOnesLogic_6_6;
  wire       [2:0]    _zz_s0_countOnesLogic_6_7;
  wire       [2:0]    _zz_s0_countOnesLogic_6_8;
  wire       [2:0]    s0_countOnesLogic_6;
  wire       [3:0]    _zz_s0_countOnesLogic_7_1;
  wire       [3:0]    _zz_s0_countOnesLogic_7_2;
  wire       [3:0]    _zz_s0_countOnesLogic_7_3;
  wire       [3:0]    _zz_s0_countOnesLogic_7_4;
  wire       [3:0]    _zz_s0_countOnesLogic_7_5;
  wire       [3:0]    _zz_s0_countOnesLogic_7_6;
  wire       [3:0]    _zz_s0_countOnesLogic_7_7;
  wire       [3:0]    _zz_s0_countOnesLogic_7_8;
  wire       [3:0]    s0_countOnesLogic_7;
  wire       [3:0]    _zz_s0_countOnesLogic_8_1;
  wire       [3:0]    _zz_s0_countOnesLogic_8_2;
  wire       [3:0]    _zz_s0_countOnesLogic_8_3;
  wire       [3:0]    _zz_s0_countOnesLogic_8_4;
  wire       [3:0]    _zz_s0_countOnesLogic_8_5;
  wire       [3:0]    _zz_s0_countOnesLogic_8_6;
  wire       [3:0]    _zz_s0_countOnesLogic_8_7;
  wire       [3:0]    _zz_s0_countOnesLogic_8_8;
  wire       [3:0]    s0_countOnesLogic_8;
  wire       [3:0]    _zz_s0_countOnesLogic_9_1;
  wire       [3:0]    _zz_s0_countOnesLogic_9_2;
  wire       [3:0]    _zz_s0_countOnesLogic_9_3;
  wire       [3:0]    _zz_s0_countOnesLogic_9_4;
  wire       [3:0]    _zz_s0_countOnesLogic_9_5;
  wire       [3:0]    _zz_s0_countOnesLogic_9_6;
  wire       [3:0]    _zz_s0_countOnesLogic_9_7;
  wire       [3:0]    _zz_s0_countOnesLogic_9_8;
  wire       [3:0]    s0_countOnesLogic_9;
  wire       [3:0]    _zz_s0_countOnesLogic_10_1;
  wire       [3:0]    _zz_s0_countOnesLogic_10_2;
  wire       [3:0]    _zz_s0_countOnesLogic_10_3;
  wire       [3:0]    _zz_s0_countOnesLogic_10_4;
  wire       [3:0]    _zz_s0_countOnesLogic_10_5;
  wire       [3:0]    _zz_s0_countOnesLogic_10_6;
  wire       [3:0]    _zz_s0_countOnesLogic_10_7;
  wire       [3:0]    _zz_s0_countOnesLogic_10_8;
  wire       [3:0]    s0_countOnesLogic_10;
  wire       [3:0]    _zz_s0_countOnesLogic_11_1;
  wire       [3:0]    _zz_s0_countOnesLogic_11_2;
  wire       [3:0]    _zz_s0_countOnesLogic_11_3;
  wire       [3:0]    _zz_s0_countOnesLogic_11_4;
  wire       [3:0]    _zz_s0_countOnesLogic_11_5;
  wire       [3:0]    _zz_s0_countOnesLogic_11_6;
  wire       [3:0]    _zz_s0_countOnesLogic_11_7;
  wire       [3:0]    _zz_s0_countOnesLogic_11_8;
  wire       [3:0]    s0_countOnesLogic_11;
  wire       [3:0]    _zz_s0_countOnesLogic_12_1;
  wire       [3:0]    _zz_s0_countOnesLogic_12_2;
  wire       [3:0]    _zz_s0_countOnesLogic_12_3;
  wire       [3:0]    _zz_s0_countOnesLogic_12_4;
  wire       [3:0]    _zz_s0_countOnesLogic_12_5;
  wire       [3:0]    _zz_s0_countOnesLogic_12_6;
  wire       [3:0]    _zz_s0_countOnesLogic_12_7;
  wire       [3:0]    _zz_s0_countOnesLogic_12_8;
  wire       [3:0]    s0_countOnesLogic_12;
  wire       [3:0]    _zz_s0_countOnesLogic_13_1;
  wire       [3:0]    _zz_s0_countOnesLogic_13_2;
  wire       [3:0]    _zz_s0_countOnesLogic_13_3;
  wire       [3:0]    _zz_s0_countOnesLogic_13_4;
  wire       [3:0]    _zz_s0_countOnesLogic_13_5;
  wire       [3:0]    _zz_s0_countOnesLogic_13_6;
  wire       [3:0]    _zz_s0_countOnesLogic_13_7;
  wire       [3:0]    _zz_s0_countOnesLogic_13_8;
  wire       [3:0]    s0_countOnesLogic_13;
  wire       [3:0]    _zz_s0_countOnesLogic_14_1;
  wire       [3:0]    _zz_s0_countOnesLogic_14_2;
  wire       [3:0]    _zz_s0_countOnesLogic_14_3;
  wire       [3:0]    _zz_s0_countOnesLogic_14_4;
  wire       [3:0]    _zz_s0_countOnesLogic_14_5;
  wire       [3:0]    _zz_s0_countOnesLogic_14_6;
  wire       [3:0]    _zz_s0_countOnesLogic_14_7;
  wire       [3:0]    _zz_s0_countOnesLogic_14_8;
  wire       [3:0]    s0_countOnesLogic_14;
  wire       [4:0]    _zz_s0_countOnesLogic_15_1;
  wire       [4:0]    _zz_s0_countOnesLogic_15_2;
  wire       [4:0]    _zz_s0_countOnesLogic_15_3;
  wire       [4:0]    _zz_s0_countOnesLogic_15_4;
  wire       [4:0]    _zz_s0_countOnesLogic_15_5;
  wire       [4:0]    _zz_s0_countOnesLogic_15_6;
  wire       [4:0]    _zz_s0_countOnesLogic_15_7;
  wire       [4:0]    _zz_s0_countOnesLogic_15_8;
  wire       [4:0]    s0_countOnesLogic_15;
  wire       [4:0]    _zz_s0_countOnesLogic_16_1;
  wire       [4:0]    _zz_s0_countOnesLogic_16_2;
  wire       [4:0]    _zz_s0_countOnesLogic_16_3;
  wire       [4:0]    _zz_s0_countOnesLogic_16_4;
  wire       [4:0]    _zz_s0_countOnesLogic_16_5;
  wire       [4:0]    _zz_s0_countOnesLogic_16_6;
  wire       [4:0]    _zz_s0_countOnesLogic_16_7;
  wire       [4:0]    _zz_s0_countOnesLogic_16_8;
  wire       [4:0]    s0_countOnesLogic_16;
  wire       [4:0]    _zz_s0_countOnesLogic_17_1;
  wire       [4:0]    _zz_s0_countOnesLogic_17_2;
  wire       [4:0]    _zz_s0_countOnesLogic_17_3;
  wire       [4:0]    _zz_s0_countOnesLogic_17_4;
  wire       [4:0]    _zz_s0_countOnesLogic_17_5;
  wire       [4:0]    _zz_s0_countOnesLogic_17_6;
  wire       [4:0]    _zz_s0_countOnesLogic_17_7;
  wire       [4:0]    _zz_s0_countOnesLogic_17_8;
  wire       [4:0]    s0_countOnesLogic_17;
  wire       [4:0]    _zz_s0_countOnesLogic_18_1;
  wire       [4:0]    _zz_s0_countOnesLogic_18_2;
  wire       [4:0]    _zz_s0_countOnesLogic_18_3;
  wire       [4:0]    _zz_s0_countOnesLogic_18_4;
  wire       [4:0]    _zz_s0_countOnesLogic_18_5;
  wire       [4:0]    _zz_s0_countOnesLogic_18_6;
  wire       [4:0]    _zz_s0_countOnesLogic_18_7;
  wire       [4:0]    _zz_s0_countOnesLogic_18_8;
  wire       [4:0]    s0_countOnesLogic_18;
  wire       [4:0]    _zz_s0_countOnesLogic_19_1;
  wire       [4:0]    _zz_s0_countOnesLogic_19_2;
  wire       [4:0]    _zz_s0_countOnesLogic_19_3;
  wire       [4:0]    _zz_s0_countOnesLogic_19_4;
  wire       [4:0]    _zz_s0_countOnesLogic_19_5;
  wire       [4:0]    _zz_s0_countOnesLogic_19_6;
  wire       [4:0]    _zz_s0_countOnesLogic_19_7;
  wire       [4:0]    _zz_s0_countOnesLogic_19_8;
  wire       [4:0]    s0_countOnesLogic_19;
  wire       [4:0]    _zz_s0_countOnesLogic_20_1;
  wire       [4:0]    _zz_s0_countOnesLogic_20_2;
  wire       [4:0]    _zz_s0_countOnesLogic_20_3;
  wire       [4:0]    _zz_s0_countOnesLogic_20_4;
  wire       [4:0]    _zz_s0_countOnesLogic_20_5;
  wire       [4:0]    _zz_s0_countOnesLogic_20_6;
  wire       [4:0]    _zz_s0_countOnesLogic_20_7;
  wire       [4:0]    _zz_s0_countOnesLogic_20_8;
  wire       [4:0]    s0_countOnesLogic_20;
  wire       [4:0]    _zz_s0_countOnesLogic_21_1;
  wire       [4:0]    _zz_s0_countOnesLogic_21_2;
  wire       [4:0]    _zz_s0_countOnesLogic_21_3;
  wire       [4:0]    _zz_s0_countOnesLogic_21_4;
  wire       [4:0]    _zz_s0_countOnesLogic_21_5;
  wire       [4:0]    _zz_s0_countOnesLogic_21_6;
  wire       [4:0]    _zz_s0_countOnesLogic_21_7;
  wire       [4:0]    _zz_s0_countOnesLogic_21_8;
  wire       [4:0]    s0_countOnesLogic_21;
  wire       [4:0]    _zz_s0_countOnesLogic_22_1;
  wire       [4:0]    _zz_s0_countOnesLogic_22_2;
  wire       [4:0]    _zz_s0_countOnesLogic_22_3;
  wire       [4:0]    _zz_s0_countOnesLogic_22_4;
  wire       [4:0]    _zz_s0_countOnesLogic_22_5;
  wire       [4:0]    _zz_s0_countOnesLogic_22_6;
  wire       [4:0]    _zz_s0_countOnesLogic_22_7;
  wire       [4:0]    _zz_s0_countOnesLogic_22_8;
  wire       [4:0]    s0_countOnesLogic_22;
  wire       [4:0]    _zz_s0_countOnesLogic_23_1;
  wire       [4:0]    _zz_s0_countOnesLogic_23_2;
  wire       [4:0]    _zz_s0_countOnesLogic_23_3;
  wire       [4:0]    _zz_s0_countOnesLogic_23_4;
  wire       [4:0]    _zz_s0_countOnesLogic_23_5;
  wire       [4:0]    _zz_s0_countOnesLogic_23_6;
  wire       [4:0]    _zz_s0_countOnesLogic_23_7;
  wire       [4:0]    _zz_s0_countOnesLogic_23_8;
  wire       [4:0]    s0_countOnesLogic_23;
  wire       [4:0]    _zz_s0_countOnesLogic_24_1;
  wire       [4:0]    _zz_s0_countOnesLogic_24_2;
  wire       [4:0]    _zz_s0_countOnesLogic_24_3;
  wire       [4:0]    _zz_s0_countOnesLogic_24_4;
  wire       [4:0]    _zz_s0_countOnesLogic_24_5;
  wire       [4:0]    _zz_s0_countOnesLogic_24_6;
  wire       [4:0]    _zz_s0_countOnesLogic_24_7;
  wire       [4:0]    _zz_s0_countOnesLogic_24_8;
  wire       [4:0]    s0_countOnesLogic_24;
  wire       [4:0]    _zz_s0_countOnesLogic_25_1;
  wire       [4:0]    _zz_s0_countOnesLogic_25_2;
  wire       [4:0]    _zz_s0_countOnesLogic_25_3;
  wire       [4:0]    _zz_s0_countOnesLogic_25_4;
  wire       [4:0]    _zz_s0_countOnesLogic_25_5;
  wire       [4:0]    _zz_s0_countOnesLogic_25_6;
  wire       [4:0]    _zz_s0_countOnesLogic_25_7;
  wire       [4:0]    _zz_s0_countOnesLogic_25_8;
  wire       [4:0]    s0_countOnesLogic_25;
  wire       [4:0]    _zz_s0_countOnesLogic_26_1;
  wire       [4:0]    _zz_s0_countOnesLogic_26_2;
  wire       [4:0]    _zz_s0_countOnesLogic_26_3;
  wire       [4:0]    _zz_s0_countOnesLogic_26_4;
  wire       [4:0]    _zz_s0_countOnesLogic_26_5;
  wire       [4:0]    _zz_s0_countOnesLogic_26_6;
  wire       [4:0]    _zz_s0_countOnesLogic_26_7;
  wire       [4:0]    _zz_s0_countOnesLogic_26_8;
  wire       [4:0]    s0_countOnesLogic_26;
  wire       [4:0]    _zz_s0_countOnesLogic_27_1;
  wire       [4:0]    _zz_s0_countOnesLogic_27_2;
  wire       [4:0]    _zz_s0_countOnesLogic_27_3;
  wire       [4:0]    _zz_s0_countOnesLogic_27_4;
  wire       [4:0]    _zz_s0_countOnesLogic_27_5;
  wire       [4:0]    _zz_s0_countOnesLogic_27_6;
  wire       [4:0]    _zz_s0_countOnesLogic_27_7;
  wire       [4:0]    _zz_s0_countOnesLogic_27_8;
  wire       [4:0]    s0_countOnesLogic_27;
  wire       [4:0]    _zz_s0_countOnesLogic_28_1;
  wire       [4:0]    _zz_s0_countOnesLogic_28_2;
  wire       [4:0]    _zz_s0_countOnesLogic_28_3;
  wire       [4:0]    _zz_s0_countOnesLogic_28_4;
  wire       [4:0]    _zz_s0_countOnesLogic_28_5;
  wire       [4:0]    _zz_s0_countOnesLogic_28_6;
  wire       [4:0]    _zz_s0_countOnesLogic_28_7;
  wire       [4:0]    _zz_s0_countOnesLogic_28_8;
  wire       [4:0]    s0_countOnesLogic_28;
  wire       [4:0]    _zz_s0_countOnesLogic_29_1;
  wire       [4:0]    _zz_s0_countOnesLogic_29_2;
  wire       [4:0]    _zz_s0_countOnesLogic_29_3;
  wire       [4:0]    _zz_s0_countOnesLogic_29_4;
  wire       [4:0]    _zz_s0_countOnesLogic_29_5;
  wire       [4:0]    _zz_s0_countOnesLogic_29_6;
  wire       [4:0]    _zz_s0_countOnesLogic_29_7;
  wire       [4:0]    _zz_s0_countOnesLogic_29_8;
  wire       [4:0]    s0_countOnesLogic_29;
  wire       [4:0]    _zz_s0_countOnesLogic_30_1;
  wire       [4:0]    _zz_s0_countOnesLogic_30_2;
  wire       [4:0]    _zz_s0_countOnesLogic_30_3;
  wire       [4:0]    _zz_s0_countOnesLogic_30_4;
  wire       [4:0]    _zz_s0_countOnesLogic_30_5;
  wire       [4:0]    _zz_s0_countOnesLogic_30_6;
  wire       [4:0]    _zz_s0_countOnesLogic_30_7;
  wire       [4:0]    _zz_s0_countOnesLogic_30_8;
  wire       [4:0]    s0_countOnesLogic_30;
  wire       [5:0]    _zz_s0_countOnesLogic_31;
  wire       [5:0]    _zz_s0_countOnesLogic_31_1;
  wire       [5:0]    _zz_s0_countOnesLogic_31_2;
  wire       [5:0]    _zz_s0_countOnesLogic_31_3;
  wire       [5:0]    _zz_s0_countOnesLogic_31_4;
  wire       [5:0]    _zz_s0_countOnesLogic_31_5;
  wire       [5:0]    _zz_s0_countOnesLogic_31_6;
  wire       [5:0]    _zz_s0_countOnesLogic_31_7;
  wire       [5:0]    s0_countOnesLogic_31;
  wire       [255:0]  s0_outputPayload_cmd_data;
  wire       [31:0]   s0_outputPayload_cmd_mask;
  wire       [0:0]    s0_outputPayload_countOnes_0;
  wire       [1:0]    s0_outputPayload_countOnes_1;
  wire       [1:0]    s0_outputPayload_countOnes_2;
  wire       [2:0]    s0_outputPayload_countOnes_3;
  wire       [2:0]    s0_outputPayload_countOnes_4;
  wire       [2:0]    s0_outputPayload_countOnes_5;
  wire       [2:0]    s0_outputPayload_countOnes_6;
  wire       [3:0]    s0_outputPayload_countOnes_7;
  wire       [3:0]    s0_outputPayload_countOnes_8;
  wire       [3:0]    s0_outputPayload_countOnes_9;
  wire       [3:0]    s0_outputPayload_countOnes_10;
  wire       [3:0]    s0_outputPayload_countOnes_11;
  wire       [3:0]    s0_outputPayload_countOnes_12;
  wire       [3:0]    s0_outputPayload_countOnes_13;
  wire       [3:0]    s0_outputPayload_countOnes_14;
  wire       [4:0]    s0_outputPayload_countOnes_15;
  wire       [4:0]    s0_outputPayload_countOnes_16;
  wire       [4:0]    s0_outputPayload_countOnes_17;
  wire       [4:0]    s0_outputPayload_countOnes_18;
  wire       [4:0]    s0_outputPayload_countOnes_19;
  wire       [4:0]    s0_outputPayload_countOnes_20;
  wire       [4:0]    s0_outputPayload_countOnes_21;
  wire       [4:0]    s0_outputPayload_countOnes_22;
  wire       [4:0]    s0_outputPayload_countOnes_23;
  wire       [4:0]    s0_outputPayload_countOnes_24;
  wire       [4:0]    s0_outputPayload_countOnes_25;
  wire       [4:0]    s0_outputPayload_countOnes_26;
  wire       [4:0]    s0_outputPayload_countOnes_27;
  wire       [4:0]    s0_outputPayload_countOnes_28;
  wire       [4:0]    s0_outputPayload_countOnes_29;
  wire       [4:0]    s0_outputPayload_countOnes_30;
  wire       [5:0]    s0_outputPayload_countOnes_31;
  wire                s0_output_valid;
  reg                 s0_output_ready;
  wire       [255:0]  s0_output_payload_cmd_data;
  wire       [31:0]   s0_output_payload_cmd_mask;
  wire       [0:0]    s0_output_payload_countOnes_0;
  wire       [1:0]    s0_output_payload_countOnes_1;
  wire       [1:0]    s0_output_payload_countOnes_2;
  wire       [2:0]    s0_output_payload_countOnes_3;
  wire       [2:0]    s0_output_payload_countOnes_4;
  wire       [2:0]    s0_output_payload_countOnes_5;
  wire       [2:0]    s0_output_payload_countOnes_6;
  wire       [3:0]    s0_output_payload_countOnes_7;
  wire       [3:0]    s0_output_payload_countOnes_8;
  wire       [3:0]    s0_output_payload_countOnes_9;
  wire       [3:0]    s0_output_payload_countOnes_10;
  wire       [3:0]    s0_output_payload_countOnes_11;
  wire       [3:0]    s0_output_payload_countOnes_12;
  wire       [3:0]    s0_output_payload_countOnes_13;
  wire       [3:0]    s0_output_payload_countOnes_14;
  wire       [4:0]    s0_output_payload_countOnes_15;
  wire       [4:0]    s0_output_payload_countOnes_16;
  wire       [4:0]    s0_output_payload_countOnes_17;
  wire       [4:0]    s0_output_payload_countOnes_18;
  wire       [4:0]    s0_output_payload_countOnes_19;
  wire       [4:0]    s0_output_payload_countOnes_20;
  wire       [4:0]    s0_output_payload_countOnes_21;
  wire       [4:0]    s0_output_payload_countOnes_22;
  wire       [4:0]    s0_output_payload_countOnes_23;
  wire       [4:0]    s0_output_payload_countOnes_24;
  wire       [4:0]    s0_output_payload_countOnes_25;
  wire       [4:0]    s0_output_payload_countOnes_26;
  wire       [4:0]    s0_output_payload_countOnes_27;
  wire       [4:0]    s0_output_payload_countOnes_28;
  wire       [4:0]    s0_output_payload_countOnes_29;
  wire       [4:0]    s0_output_payload_countOnes_30;
  wire       [5:0]    s0_output_payload_countOnes_31;
  wire                s1_input_valid;
  wire                s1_input_ready;
  wire       [255:0]  s1_input_payload_cmd_data;
  wire       [31:0]   s1_input_payload_cmd_mask;
  wire       [0:0]    s1_input_payload_countOnes_0;
  wire       [1:0]    s1_input_payload_countOnes_1;
  wire       [1:0]    s1_input_payload_countOnes_2;
  wire       [2:0]    s1_input_payload_countOnes_3;
  wire       [2:0]    s1_input_payload_countOnes_4;
  wire       [2:0]    s1_input_payload_countOnes_5;
  wire       [2:0]    s1_input_payload_countOnes_6;
  wire       [3:0]    s1_input_payload_countOnes_7;
  wire       [3:0]    s1_input_payload_countOnes_8;
  wire       [3:0]    s1_input_payload_countOnes_9;
  wire       [3:0]    s1_input_payload_countOnes_10;
  wire       [3:0]    s1_input_payload_countOnes_11;
  wire       [3:0]    s1_input_payload_countOnes_12;
  wire       [3:0]    s1_input_payload_countOnes_13;
  wire       [3:0]    s1_input_payload_countOnes_14;
  wire       [4:0]    s1_input_payload_countOnes_15;
  wire       [4:0]    s1_input_payload_countOnes_16;
  wire       [4:0]    s1_input_payload_countOnes_17;
  wire       [4:0]    s1_input_payload_countOnes_18;
  wire       [4:0]    s1_input_payload_countOnes_19;
  wire       [4:0]    s1_input_payload_countOnes_20;
  wire       [4:0]    s1_input_payload_countOnes_21;
  wire       [4:0]    s1_input_payload_countOnes_22;
  wire       [4:0]    s1_input_payload_countOnes_23;
  wire       [4:0]    s1_input_payload_countOnes_24;
  wire       [4:0]    s1_input_payload_countOnes_25;
  wire       [4:0]    s1_input_payload_countOnes_26;
  wire       [4:0]    s1_input_payload_countOnes_27;
  wire       [4:0]    s1_input_payload_countOnes_28;
  wire       [4:0]    s1_input_payload_countOnes_29;
  wire       [4:0]    s1_input_payload_countOnes_30;
  wire       [5:0]    s1_input_payload_countOnes_31;
  reg                 s0_output_rValid;
  reg        [255:0]  s0_output_rData_cmd_data;
  reg        [31:0]   s0_output_rData_cmd_mask;
  reg        [0:0]    s0_output_rData_countOnes_0;
  reg        [1:0]    s0_output_rData_countOnes_1;
  reg        [1:0]    s0_output_rData_countOnes_2;
  reg        [2:0]    s0_output_rData_countOnes_3;
  reg        [2:0]    s0_output_rData_countOnes_4;
  reg        [2:0]    s0_output_rData_countOnes_5;
  reg        [2:0]    s0_output_rData_countOnes_6;
  reg        [3:0]    s0_output_rData_countOnes_7;
  reg        [3:0]    s0_output_rData_countOnes_8;
  reg        [3:0]    s0_output_rData_countOnes_9;
  reg        [3:0]    s0_output_rData_countOnes_10;
  reg        [3:0]    s0_output_rData_countOnes_11;
  reg        [3:0]    s0_output_rData_countOnes_12;
  reg        [3:0]    s0_output_rData_countOnes_13;
  reg        [3:0]    s0_output_rData_countOnes_14;
  reg        [4:0]    s0_output_rData_countOnes_15;
  reg        [4:0]    s0_output_rData_countOnes_16;
  reg        [4:0]    s0_output_rData_countOnes_17;
  reg        [4:0]    s0_output_rData_countOnes_18;
  reg        [4:0]    s0_output_rData_countOnes_19;
  reg        [4:0]    s0_output_rData_countOnes_20;
  reg        [4:0]    s0_output_rData_countOnes_21;
  reg        [4:0]    s0_output_rData_countOnes_22;
  reg        [4:0]    s0_output_rData_countOnes_23;
  reg        [4:0]    s0_output_rData_countOnes_24;
  reg        [4:0]    s0_output_rData_countOnes_25;
  reg        [4:0]    s0_output_rData_countOnes_26;
  reg        [4:0]    s0_output_rData_countOnes_27;
  reg        [4:0]    s0_output_rData_countOnes_28;
  reg        [4:0]    s0_output_rData_countOnes_29;
  reg        [4:0]    s0_output_rData_countOnes_30;
  reg        [5:0]    s0_output_rData_countOnes_31;
  wire                when_Stream_l375_1;
  reg        [4:0]    s1_offset;
  wire       [5:0]    s1_offsetNext;
  wire                s1_input_fire;
  reg        [13:0]   s1_byteCounter;
  wire       [4:0]    s1_inputIndexes_0;
  wire       [4:0]    s1_inputIndexes_1;
  wire       [4:0]    s1_inputIndexes_2;
  wire       [4:0]    s1_inputIndexes_3;
  wire       [4:0]    s1_inputIndexes_4;
  wire       [4:0]    s1_inputIndexes_5;
  wire       [4:0]    s1_inputIndexes_6;
  wire       [4:0]    s1_inputIndexes_7;
  wire       [4:0]    s1_inputIndexes_8;
  wire       [4:0]    s1_inputIndexes_9;
  wire       [4:0]    s1_inputIndexes_10;
  wire       [4:0]    s1_inputIndexes_11;
  wire       [4:0]    s1_inputIndexes_12;
  wire       [4:0]    s1_inputIndexes_13;
  wire       [4:0]    s1_inputIndexes_14;
  wire       [4:0]    s1_inputIndexes_15;
  wire       [4:0]    s1_inputIndexes_16;
  wire       [4:0]    s1_inputIndexes_17;
  wire       [4:0]    s1_inputIndexes_18;
  wire       [4:0]    s1_inputIndexes_19;
  wire       [4:0]    s1_inputIndexes_20;
  wire       [4:0]    s1_inputIndexes_21;
  wire       [4:0]    s1_inputIndexes_22;
  wire       [4:0]    s1_inputIndexes_23;
  wire       [4:0]    s1_inputIndexes_24;
  wire       [4:0]    s1_inputIndexes_25;
  wire       [4:0]    s1_inputIndexes_26;
  wire       [4:0]    s1_inputIndexes_27;
  wire       [4:0]    s1_inputIndexes_28;
  wire       [4:0]    s1_inputIndexes_29;
  wire       [4:0]    s1_inputIndexes_30;
  wire       [4:0]    s1_inputIndexes_31;
  wire       [255:0]  s1_outputPayload_cmd_data;
  wire       [31:0]   s1_outputPayload_cmd_mask;
  wire       [4:0]    s1_outputPayload_index_0;
  wire       [4:0]    s1_outputPayload_index_1;
  wire       [4:0]    s1_outputPayload_index_2;
  wire       [4:0]    s1_outputPayload_index_3;
  wire       [4:0]    s1_outputPayload_index_4;
  wire       [4:0]    s1_outputPayload_index_5;
  wire       [4:0]    s1_outputPayload_index_6;
  wire       [4:0]    s1_outputPayload_index_7;
  wire       [4:0]    s1_outputPayload_index_8;
  wire       [4:0]    s1_outputPayload_index_9;
  wire       [4:0]    s1_outputPayload_index_10;
  wire       [4:0]    s1_outputPayload_index_11;
  wire       [4:0]    s1_outputPayload_index_12;
  wire       [4:0]    s1_outputPayload_index_13;
  wire       [4:0]    s1_outputPayload_index_14;
  wire       [4:0]    s1_outputPayload_index_15;
  wire       [4:0]    s1_outputPayload_index_16;
  wire       [4:0]    s1_outputPayload_index_17;
  wire       [4:0]    s1_outputPayload_index_18;
  wire       [4:0]    s1_outputPayload_index_19;
  wire       [4:0]    s1_outputPayload_index_20;
  wire       [4:0]    s1_outputPayload_index_21;
  wire       [4:0]    s1_outputPayload_index_22;
  wire       [4:0]    s1_outputPayload_index_23;
  wire       [4:0]    s1_outputPayload_index_24;
  wire       [4:0]    s1_outputPayload_index_25;
  wire       [4:0]    s1_outputPayload_index_26;
  wire       [4:0]    s1_outputPayload_index_27;
  wire       [4:0]    s1_outputPayload_index_28;
  wire       [4:0]    s1_outputPayload_index_29;
  wire       [4:0]    s1_outputPayload_index_30;
  wire       [4:0]    s1_outputPayload_index_31;
  wire                s1_outputPayload_last;
  wire       [4:0]    s1_outputPayload_sel_0;
  wire       [4:0]    s1_outputPayload_sel_1;
  wire       [4:0]    s1_outputPayload_sel_2;
  wire       [4:0]    s1_outputPayload_sel_3;
  wire       [4:0]    s1_outputPayload_sel_4;
  wire       [4:0]    s1_outputPayload_sel_5;
  wire       [4:0]    s1_outputPayload_sel_6;
  wire       [4:0]    s1_outputPayload_sel_7;
  wire       [4:0]    s1_outputPayload_sel_8;
  wire       [4:0]    s1_outputPayload_sel_9;
  wire       [4:0]    s1_outputPayload_sel_10;
  wire       [4:0]    s1_outputPayload_sel_11;
  wire       [4:0]    s1_outputPayload_sel_12;
  wire       [4:0]    s1_outputPayload_sel_13;
  wire       [4:0]    s1_outputPayload_sel_14;
  wire       [4:0]    s1_outputPayload_sel_15;
  wire       [4:0]    s1_outputPayload_sel_16;
  wire       [4:0]    s1_outputPayload_sel_17;
  wire       [4:0]    s1_outputPayload_sel_18;
  wire       [4:0]    s1_outputPayload_sel_19;
  wire       [4:0]    s1_outputPayload_sel_20;
  wire       [4:0]    s1_outputPayload_sel_21;
  wire       [4:0]    s1_outputPayload_sel_22;
  wire       [4:0]    s1_outputPayload_sel_23;
  wire       [4:0]    s1_outputPayload_sel_24;
  wire       [4:0]    s1_outputPayload_sel_25;
  wire       [4:0]    s1_outputPayload_sel_26;
  wire       [4:0]    s1_outputPayload_sel_27;
  wire       [4:0]    s1_outputPayload_sel_28;
  wire       [4:0]    s1_outputPayload_sel_29;
  wire       [4:0]    s1_outputPayload_sel_30;
  wire       [4:0]    s1_outputPayload_sel_31;
  reg        [31:0]   s1_outputPayload_selValid;
  wire                _zz_s1_outputPayload_selValid;
  wire                _zz_s1_outputPayload_selValid_1;
  wire                _zz_s1_outputPayload_selValid_2;
  wire                _zz_s1_outputPayload_selValid_3;
  wire                _zz_s1_outputPayload_selValid_4;
  wire                _zz_s1_outputPayload_selValid_5;
  wire                _zz_s1_outputPayload_selValid_6;
  wire                _zz_s1_outputPayload_selValid_7;
  wire                _zz_s1_outputPayload_selValid_8;
  wire                _zz_s1_outputPayload_selValid_9;
  wire                _zz_s1_outputPayload_selValid_10;
  wire                _zz_s1_outputPayload_selValid_11;
  wire                _zz_s1_outputPayload_selValid_12;
  wire                _zz_s1_outputPayload_selValid_13;
  wire                _zz_s1_outputPayload_selValid_14;
  wire                _zz_s1_outputPayload_selValid_15;
  wire                _zz_s1_outputPayload_selValid_16;
  wire                _zz_s1_outputPayload_selValid_17;
  wire                _zz_s1_outputPayload_selValid_18;
  wire                _zz_s1_outputPayload_selValid_19;
  wire                _zz_s1_outputPayload_selValid_20;
  wire                _zz_s1_outputPayload_selValid_21;
  wire                _zz_s1_outputPayload_selValid_22;
  wire                _zz_s1_outputPayload_selValid_23;
  wire                _zz_s1_outputPayload_selValid_24;
  wire                _zz_s1_outputPayload_selValid_25;
  wire                _zz_s1_outputPayload_selValid_26;
  wire                _zz_s1_outputPayload_selValid_27;
  wire                _zz_s1_outputPayload_selValid_28;
  wire                _zz_s1_outputPayload_selValid_29;
  wire                _zz_s1_outputPayload_selValid_30;
  wire                _zz_s1_outputPayload_sel_0;
  wire                _zz_s1_outputPayload_sel_0_1;
  wire                _zz_s1_outputPayload_sel_0_2;
  wire                _zz_s1_outputPayload_sel_0_3;
  wire                _zz_s1_outputPayload_sel_0_4;
  wire                _zz_s1_outputPayload_selValid_31;
  wire                _zz_s1_outputPayload_selValid_32;
  wire                _zz_s1_outputPayload_selValid_33;
  wire                _zz_s1_outputPayload_selValid_34;
  wire                _zz_s1_outputPayload_selValid_35;
  wire                _zz_s1_outputPayload_selValid_36;
  wire                _zz_s1_outputPayload_selValid_37;
  wire                _zz_s1_outputPayload_selValid_38;
  wire                _zz_s1_outputPayload_selValid_39;
  wire                _zz_s1_outputPayload_selValid_40;
  wire                _zz_s1_outputPayload_selValid_41;
  wire                _zz_s1_outputPayload_selValid_42;
  wire                _zz_s1_outputPayload_selValid_43;
  wire                _zz_s1_outputPayload_selValid_44;
  wire                _zz_s1_outputPayload_selValid_45;
  wire                _zz_s1_outputPayload_selValid_46;
  wire                _zz_s1_outputPayload_selValid_47;
  wire                _zz_s1_outputPayload_selValid_48;
  wire                _zz_s1_outputPayload_selValid_49;
  wire                _zz_s1_outputPayload_selValid_50;
  wire                _zz_s1_outputPayload_selValid_51;
  wire                _zz_s1_outputPayload_selValid_52;
  wire                _zz_s1_outputPayload_selValid_53;
  wire                _zz_s1_outputPayload_selValid_54;
  wire                _zz_s1_outputPayload_selValid_55;
  wire                _zz_s1_outputPayload_selValid_56;
  wire                _zz_s1_outputPayload_selValid_57;
  wire                _zz_s1_outputPayload_selValid_58;
  wire                _zz_s1_outputPayload_selValid_59;
  wire                _zz_s1_outputPayload_selValid_60;
  wire                _zz_s1_outputPayload_selValid_61;
  wire                _zz_s1_outputPayload_sel_1;
  wire                _zz_s1_outputPayload_sel_1_1;
  wire                _zz_s1_outputPayload_sel_1_2;
  wire                _zz_s1_outputPayload_sel_1_3;
  wire                _zz_s1_outputPayload_sel_1_4;
  wire                _zz_s1_outputPayload_selValid_62;
  wire                _zz_s1_outputPayload_selValid_63;
  wire                _zz_s1_outputPayload_selValid_64;
  wire                _zz_s1_outputPayload_selValid_65;
  wire                _zz_s1_outputPayload_selValid_66;
  wire                _zz_s1_outputPayload_selValid_67;
  wire                _zz_s1_outputPayload_selValid_68;
  wire                _zz_s1_outputPayload_selValid_69;
  wire                _zz_s1_outputPayload_selValid_70;
  wire                _zz_s1_outputPayload_selValid_71;
  wire                _zz_s1_outputPayload_selValid_72;
  wire                _zz_s1_outputPayload_selValid_73;
  wire                _zz_s1_outputPayload_selValid_74;
  wire                _zz_s1_outputPayload_selValid_75;
  wire                _zz_s1_outputPayload_selValid_76;
  wire                _zz_s1_outputPayload_selValid_77;
  wire                _zz_s1_outputPayload_selValid_78;
  wire                _zz_s1_outputPayload_selValid_79;
  wire                _zz_s1_outputPayload_selValid_80;
  wire                _zz_s1_outputPayload_selValid_81;
  wire                _zz_s1_outputPayload_selValid_82;
  wire                _zz_s1_outputPayload_selValid_83;
  wire                _zz_s1_outputPayload_selValid_84;
  wire                _zz_s1_outputPayload_selValid_85;
  wire                _zz_s1_outputPayload_selValid_86;
  wire                _zz_s1_outputPayload_selValid_87;
  wire                _zz_s1_outputPayload_selValid_88;
  wire                _zz_s1_outputPayload_selValid_89;
  wire                _zz_s1_outputPayload_selValid_90;
  wire                _zz_s1_outputPayload_selValid_91;
  wire                _zz_s1_outputPayload_selValid_92;
  wire                _zz_s1_outputPayload_sel_2;
  wire                _zz_s1_outputPayload_sel_2_1;
  wire                _zz_s1_outputPayload_sel_2_2;
  wire                _zz_s1_outputPayload_sel_2_3;
  wire                _zz_s1_outputPayload_sel_2_4;
  wire                _zz_s1_outputPayload_selValid_93;
  wire                _zz_s1_outputPayload_selValid_94;
  wire                _zz_s1_outputPayload_selValid_95;
  wire                _zz_s1_outputPayload_selValid_96;
  wire                _zz_s1_outputPayload_selValid_97;
  wire                _zz_s1_outputPayload_selValid_98;
  wire                _zz_s1_outputPayload_selValid_99;
  wire                _zz_s1_outputPayload_selValid_100;
  wire                _zz_s1_outputPayload_selValid_101;
  wire                _zz_s1_outputPayload_selValid_102;
  wire                _zz_s1_outputPayload_selValid_103;
  wire                _zz_s1_outputPayload_selValid_104;
  wire                _zz_s1_outputPayload_selValid_105;
  wire                _zz_s1_outputPayload_selValid_106;
  wire                _zz_s1_outputPayload_selValid_107;
  wire                _zz_s1_outputPayload_selValid_108;
  wire                _zz_s1_outputPayload_selValid_109;
  wire                _zz_s1_outputPayload_selValid_110;
  wire                _zz_s1_outputPayload_selValid_111;
  wire                _zz_s1_outputPayload_selValid_112;
  wire                _zz_s1_outputPayload_selValid_113;
  wire                _zz_s1_outputPayload_selValid_114;
  wire                _zz_s1_outputPayload_selValid_115;
  wire                _zz_s1_outputPayload_selValid_116;
  wire                _zz_s1_outputPayload_selValid_117;
  wire                _zz_s1_outputPayload_selValid_118;
  wire                _zz_s1_outputPayload_selValid_119;
  wire                _zz_s1_outputPayload_selValid_120;
  wire                _zz_s1_outputPayload_selValid_121;
  wire                _zz_s1_outputPayload_selValid_122;
  wire                _zz_s1_outputPayload_selValid_123;
  wire                _zz_s1_outputPayload_sel_3;
  wire                _zz_s1_outputPayload_sel_3_1;
  wire                _zz_s1_outputPayload_sel_3_2;
  wire                _zz_s1_outputPayload_sel_3_3;
  wire                _zz_s1_outputPayload_sel_3_4;
  wire                _zz_s1_outputPayload_selValid_124;
  wire                _zz_s1_outputPayload_selValid_125;
  wire                _zz_s1_outputPayload_selValid_126;
  wire                _zz_s1_outputPayload_selValid_127;
  wire                _zz_s1_outputPayload_selValid_128;
  wire                _zz_s1_outputPayload_selValid_129;
  wire                _zz_s1_outputPayload_selValid_130;
  wire                _zz_s1_outputPayload_selValid_131;
  wire                _zz_s1_outputPayload_selValid_132;
  wire                _zz_s1_outputPayload_selValid_133;
  wire                _zz_s1_outputPayload_selValid_134;
  wire                _zz_s1_outputPayload_selValid_135;
  wire                _zz_s1_outputPayload_selValid_136;
  wire                _zz_s1_outputPayload_selValid_137;
  wire                _zz_s1_outputPayload_selValid_138;
  wire                _zz_s1_outputPayload_selValid_139;
  wire                _zz_s1_outputPayload_selValid_140;
  wire                _zz_s1_outputPayload_selValid_141;
  wire                _zz_s1_outputPayload_selValid_142;
  wire                _zz_s1_outputPayload_selValid_143;
  wire                _zz_s1_outputPayload_selValid_144;
  wire                _zz_s1_outputPayload_selValid_145;
  wire                _zz_s1_outputPayload_selValid_146;
  wire                _zz_s1_outputPayload_selValid_147;
  wire                _zz_s1_outputPayload_selValid_148;
  wire                _zz_s1_outputPayload_selValid_149;
  wire                _zz_s1_outputPayload_selValid_150;
  wire                _zz_s1_outputPayload_selValid_151;
  wire                _zz_s1_outputPayload_selValid_152;
  wire                _zz_s1_outputPayload_selValid_153;
  wire                _zz_s1_outputPayload_selValid_154;
  wire                _zz_s1_outputPayload_sel_4;
  wire                _zz_s1_outputPayload_sel_4_1;
  wire                _zz_s1_outputPayload_sel_4_2;
  wire                _zz_s1_outputPayload_sel_4_3;
  wire                _zz_s1_outputPayload_sel_4_4;
  wire                _zz_s1_outputPayload_selValid_155;
  wire                _zz_s1_outputPayload_selValid_156;
  wire                _zz_s1_outputPayload_selValid_157;
  wire                _zz_s1_outputPayload_selValid_158;
  wire                _zz_s1_outputPayload_selValid_159;
  wire                _zz_s1_outputPayload_selValid_160;
  wire                _zz_s1_outputPayload_selValid_161;
  wire                _zz_s1_outputPayload_selValid_162;
  wire                _zz_s1_outputPayload_selValid_163;
  wire                _zz_s1_outputPayload_selValid_164;
  wire                _zz_s1_outputPayload_selValid_165;
  wire                _zz_s1_outputPayload_selValid_166;
  wire                _zz_s1_outputPayload_selValid_167;
  wire                _zz_s1_outputPayload_selValid_168;
  wire                _zz_s1_outputPayload_selValid_169;
  wire                _zz_s1_outputPayload_selValid_170;
  wire                _zz_s1_outputPayload_selValid_171;
  wire                _zz_s1_outputPayload_selValid_172;
  wire                _zz_s1_outputPayload_selValid_173;
  wire                _zz_s1_outputPayload_selValid_174;
  wire                _zz_s1_outputPayload_selValid_175;
  wire                _zz_s1_outputPayload_selValid_176;
  wire                _zz_s1_outputPayload_selValid_177;
  wire                _zz_s1_outputPayload_selValid_178;
  wire                _zz_s1_outputPayload_selValid_179;
  wire                _zz_s1_outputPayload_selValid_180;
  wire                _zz_s1_outputPayload_selValid_181;
  wire                _zz_s1_outputPayload_selValid_182;
  wire                _zz_s1_outputPayload_selValid_183;
  wire                _zz_s1_outputPayload_selValid_184;
  wire                _zz_s1_outputPayload_selValid_185;
  wire                _zz_s1_outputPayload_sel_5;
  wire                _zz_s1_outputPayload_sel_5_1;
  wire                _zz_s1_outputPayload_sel_5_2;
  wire                _zz_s1_outputPayload_sel_5_3;
  wire                _zz_s1_outputPayload_sel_5_4;
  wire                _zz_s1_outputPayload_selValid_186;
  wire                _zz_s1_outputPayload_selValid_187;
  wire                _zz_s1_outputPayload_selValid_188;
  wire                _zz_s1_outputPayload_selValid_189;
  wire                _zz_s1_outputPayload_selValid_190;
  wire                _zz_s1_outputPayload_selValid_191;
  wire                _zz_s1_outputPayload_selValid_192;
  wire                _zz_s1_outputPayload_selValid_193;
  wire                _zz_s1_outputPayload_selValid_194;
  wire                _zz_s1_outputPayload_selValid_195;
  wire                _zz_s1_outputPayload_selValid_196;
  wire                _zz_s1_outputPayload_selValid_197;
  wire                _zz_s1_outputPayload_selValid_198;
  wire                _zz_s1_outputPayload_selValid_199;
  wire                _zz_s1_outputPayload_selValid_200;
  wire                _zz_s1_outputPayload_selValid_201;
  wire                _zz_s1_outputPayload_selValid_202;
  wire                _zz_s1_outputPayload_selValid_203;
  wire                _zz_s1_outputPayload_selValid_204;
  wire                _zz_s1_outputPayload_selValid_205;
  wire                _zz_s1_outputPayload_selValid_206;
  wire                _zz_s1_outputPayload_selValid_207;
  wire                _zz_s1_outputPayload_selValid_208;
  wire                _zz_s1_outputPayload_selValid_209;
  wire                _zz_s1_outputPayload_selValid_210;
  wire                _zz_s1_outputPayload_selValid_211;
  wire                _zz_s1_outputPayload_selValid_212;
  wire                _zz_s1_outputPayload_selValid_213;
  wire                _zz_s1_outputPayload_selValid_214;
  wire                _zz_s1_outputPayload_selValid_215;
  wire                _zz_s1_outputPayload_selValid_216;
  wire                _zz_s1_outputPayload_sel_6;
  wire                _zz_s1_outputPayload_sel_6_1;
  wire                _zz_s1_outputPayload_sel_6_2;
  wire                _zz_s1_outputPayload_sel_6_3;
  wire                _zz_s1_outputPayload_sel_6_4;
  wire                _zz_s1_outputPayload_selValid_217;
  wire                _zz_s1_outputPayload_selValid_218;
  wire                _zz_s1_outputPayload_selValid_219;
  wire                _zz_s1_outputPayload_selValid_220;
  wire                _zz_s1_outputPayload_selValid_221;
  wire                _zz_s1_outputPayload_selValid_222;
  wire                _zz_s1_outputPayload_selValid_223;
  wire                _zz_s1_outputPayload_selValid_224;
  wire                _zz_s1_outputPayload_selValid_225;
  wire                _zz_s1_outputPayload_selValid_226;
  wire                _zz_s1_outputPayload_selValid_227;
  wire                _zz_s1_outputPayload_selValid_228;
  wire                _zz_s1_outputPayload_selValid_229;
  wire                _zz_s1_outputPayload_selValid_230;
  wire                _zz_s1_outputPayload_selValid_231;
  wire                _zz_s1_outputPayload_selValid_232;
  wire                _zz_s1_outputPayload_selValid_233;
  wire                _zz_s1_outputPayload_selValid_234;
  wire                _zz_s1_outputPayload_selValid_235;
  wire                _zz_s1_outputPayload_selValid_236;
  wire                _zz_s1_outputPayload_selValid_237;
  wire                _zz_s1_outputPayload_selValid_238;
  wire                _zz_s1_outputPayload_selValid_239;
  wire                _zz_s1_outputPayload_selValid_240;
  wire                _zz_s1_outputPayload_selValid_241;
  wire                _zz_s1_outputPayload_selValid_242;
  wire                _zz_s1_outputPayload_selValid_243;
  wire                _zz_s1_outputPayload_selValid_244;
  wire                _zz_s1_outputPayload_selValid_245;
  wire                _zz_s1_outputPayload_selValid_246;
  wire                _zz_s1_outputPayload_selValid_247;
  wire                _zz_s1_outputPayload_sel_7;
  wire                _zz_s1_outputPayload_sel_7_1;
  wire                _zz_s1_outputPayload_sel_7_2;
  wire                _zz_s1_outputPayload_sel_7_3;
  wire                _zz_s1_outputPayload_sel_7_4;
  wire                _zz_s1_outputPayload_selValid_248;
  wire                _zz_s1_outputPayload_selValid_249;
  wire                _zz_s1_outputPayload_selValid_250;
  wire                _zz_s1_outputPayload_selValid_251;
  wire                _zz_s1_outputPayload_selValid_252;
  wire                _zz_s1_outputPayload_selValid_253;
  wire                _zz_s1_outputPayload_selValid_254;
  wire                _zz_s1_outputPayload_selValid_255;
  wire                _zz_s1_outputPayload_selValid_256;
  wire                _zz_s1_outputPayload_selValid_257;
  wire                _zz_s1_outputPayload_selValid_258;
  wire                _zz_s1_outputPayload_selValid_259;
  wire                _zz_s1_outputPayload_selValid_260;
  wire                _zz_s1_outputPayload_selValid_261;
  wire                _zz_s1_outputPayload_selValid_262;
  wire                _zz_s1_outputPayload_selValid_263;
  wire                _zz_s1_outputPayload_selValid_264;
  wire                _zz_s1_outputPayload_selValid_265;
  wire                _zz_s1_outputPayload_selValid_266;
  wire                _zz_s1_outputPayload_selValid_267;
  wire                _zz_s1_outputPayload_selValid_268;
  wire                _zz_s1_outputPayload_selValid_269;
  wire                _zz_s1_outputPayload_selValid_270;
  wire                _zz_s1_outputPayload_selValid_271;
  wire                _zz_s1_outputPayload_selValid_272;
  wire                _zz_s1_outputPayload_selValid_273;
  wire                _zz_s1_outputPayload_selValid_274;
  wire                _zz_s1_outputPayload_selValid_275;
  wire                _zz_s1_outputPayload_selValid_276;
  wire                _zz_s1_outputPayload_selValid_277;
  wire                _zz_s1_outputPayload_selValid_278;
  wire                _zz_s1_outputPayload_sel_8;
  wire                _zz_s1_outputPayload_sel_8_1;
  wire                _zz_s1_outputPayload_sel_8_2;
  wire                _zz_s1_outputPayload_sel_8_3;
  wire                _zz_s1_outputPayload_sel_8_4;
  wire                _zz_s1_outputPayload_selValid_279;
  wire                _zz_s1_outputPayload_selValid_280;
  wire                _zz_s1_outputPayload_selValid_281;
  wire                _zz_s1_outputPayload_selValid_282;
  wire                _zz_s1_outputPayload_selValid_283;
  wire                _zz_s1_outputPayload_selValid_284;
  wire                _zz_s1_outputPayload_selValid_285;
  wire                _zz_s1_outputPayload_selValid_286;
  wire                _zz_s1_outputPayload_selValid_287;
  wire                _zz_s1_outputPayload_selValid_288;
  wire                _zz_s1_outputPayload_selValid_289;
  wire                _zz_s1_outputPayload_selValid_290;
  wire                _zz_s1_outputPayload_selValid_291;
  wire                _zz_s1_outputPayload_selValid_292;
  wire                _zz_s1_outputPayload_selValid_293;
  wire                _zz_s1_outputPayload_selValid_294;
  wire                _zz_s1_outputPayload_selValid_295;
  wire                _zz_s1_outputPayload_selValid_296;
  wire                _zz_s1_outputPayload_selValid_297;
  wire                _zz_s1_outputPayload_selValid_298;
  wire                _zz_s1_outputPayload_selValid_299;
  wire                _zz_s1_outputPayload_selValid_300;
  wire                _zz_s1_outputPayload_selValid_301;
  wire                _zz_s1_outputPayload_selValid_302;
  wire                _zz_s1_outputPayload_selValid_303;
  wire                _zz_s1_outputPayload_selValid_304;
  wire                _zz_s1_outputPayload_selValid_305;
  wire                _zz_s1_outputPayload_selValid_306;
  wire                _zz_s1_outputPayload_selValid_307;
  wire                _zz_s1_outputPayload_selValid_308;
  wire                _zz_s1_outputPayload_selValid_309;
  wire                _zz_s1_outputPayload_sel_9;
  wire                _zz_s1_outputPayload_sel_9_1;
  wire                _zz_s1_outputPayload_sel_9_2;
  wire                _zz_s1_outputPayload_sel_9_3;
  wire                _zz_s1_outputPayload_sel_9_4;
  wire                _zz_s1_outputPayload_selValid_310;
  wire                _zz_s1_outputPayload_selValid_311;
  wire                _zz_s1_outputPayload_selValid_312;
  wire                _zz_s1_outputPayload_selValid_313;
  wire                _zz_s1_outputPayload_selValid_314;
  wire                _zz_s1_outputPayload_selValid_315;
  wire                _zz_s1_outputPayload_selValid_316;
  wire                _zz_s1_outputPayload_selValid_317;
  wire                _zz_s1_outputPayload_selValid_318;
  wire                _zz_s1_outputPayload_selValid_319;
  wire                _zz_s1_outputPayload_selValid_320;
  wire                _zz_s1_outputPayload_selValid_321;
  wire                _zz_s1_outputPayload_selValid_322;
  wire                _zz_s1_outputPayload_selValid_323;
  wire                _zz_s1_outputPayload_selValid_324;
  wire                _zz_s1_outputPayload_selValid_325;
  wire                _zz_s1_outputPayload_selValid_326;
  wire                _zz_s1_outputPayload_selValid_327;
  wire                _zz_s1_outputPayload_selValid_328;
  wire                _zz_s1_outputPayload_selValid_329;
  wire                _zz_s1_outputPayload_selValid_330;
  wire                _zz_s1_outputPayload_selValid_331;
  wire                _zz_s1_outputPayload_selValid_332;
  wire                _zz_s1_outputPayload_selValid_333;
  wire                _zz_s1_outputPayload_selValid_334;
  wire                _zz_s1_outputPayload_selValid_335;
  wire                _zz_s1_outputPayload_selValid_336;
  wire                _zz_s1_outputPayload_selValid_337;
  wire                _zz_s1_outputPayload_selValid_338;
  wire                _zz_s1_outputPayload_selValid_339;
  wire                _zz_s1_outputPayload_selValid_340;
  wire                _zz_s1_outputPayload_sel_10;
  wire                _zz_s1_outputPayload_sel_10_1;
  wire                _zz_s1_outputPayload_sel_10_2;
  wire                _zz_s1_outputPayload_sel_10_3;
  wire                _zz_s1_outputPayload_sel_10_4;
  wire                _zz_s1_outputPayload_selValid_341;
  wire                _zz_s1_outputPayload_selValid_342;
  wire                _zz_s1_outputPayload_selValid_343;
  wire                _zz_s1_outputPayload_selValid_344;
  wire                _zz_s1_outputPayload_selValid_345;
  wire                _zz_s1_outputPayload_selValid_346;
  wire                _zz_s1_outputPayload_selValid_347;
  wire                _zz_s1_outputPayload_selValid_348;
  wire                _zz_s1_outputPayload_selValid_349;
  wire                _zz_s1_outputPayload_selValid_350;
  wire                _zz_s1_outputPayload_selValid_351;
  wire                _zz_s1_outputPayload_selValid_352;
  wire                _zz_s1_outputPayload_selValid_353;
  wire                _zz_s1_outputPayload_selValid_354;
  wire                _zz_s1_outputPayload_selValid_355;
  wire                _zz_s1_outputPayload_selValid_356;
  wire                _zz_s1_outputPayload_selValid_357;
  wire                _zz_s1_outputPayload_selValid_358;
  wire                _zz_s1_outputPayload_selValid_359;
  wire                _zz_s1_outputPayload_selValid_360;
  wire                _zz_s1_outputPayload_selValid_361;
  wire                _zz_s1_outputPayload_selValid_362;
  wire                _zz_s1_outputPayload_selValid_363;
  wire                _zz_s1_outputPayload_selValid_364;
  wire                _zz_s1_outputPayload_selValid_365;
  wire                _zz_s1_outputPayload_selValid_366;
  wire                _zz_s1_outputPayload_selValid_367;
  wire                _zz_s1_outputPayload_selValid_368;
  wire                _zz_s1_outputPayload_selValid_369;
  wire                _zz_s1_outputPayload_selValid_370;
  wire                _zz_s1_outputPayload_selValid_371;
  wire                _zz_s1_outputPayload_sel_11;
  wire                _zz_s1_outputPayload_sel_11_1;
  wire                _zz_s1_outputPayload_sel_11_2;
  wire                _zz_s1_outputPayload_sel_11_3;
  wire                _zz_s1_outputPayload_sel_11_4;
  wire                _zz_s1_outputPayload_selValid_372;
  wire                _zz_s1_outputPayload_selValid_373;
  wire                _zz_s1_outputPayload_selValid_374;
  wire                _zz_s1_outputPayload_selValid_375;
  wire                _zz_s1_outputPayload_selValid_376;
  wire                _zz_s1_outputPayload_selValid_377;
  wire                _zz_s1_outputPayload_selValid_378;
  wire                _zz_s1_outputPayload_selValid_379;
  wire                _zz_s1_outputPayload_selValid_380;
  wire                _zz_s1_outputPayload_selValid_381;
  wire                _zz_s1_outputPayload_selValid_382;
  wire                _zz_s1_outputPayload_selValid_383;
  wire                _zz_s1_outputPayload_selValid_384;
  wire                _zz_s1_outputPayload_selValid_385;
  wire                _zz_s1_outputPayload_selValid_386;
  wire                _zz_s1_outputPayload_selValid_387;
  wire                _zz_s1_outputPayload_selValid_388;
  wire                _zz_s1_outputPayload_selValid_389;
  wire                _zz_s1_outputPayload_selValid_390;
  wire                _zz_s1_outputPayload_selValid_391;
  wire                _zz_s1_outputPayload_selValid_392;
  wire                _zz_s1_outputPayload_selValid_393;
  wire                _zz_s1_outputPayload_selValid_394;
  wire                _zz_s1_outputPayload_selValid_395;
  wire                _zz_s1_outputPayload_selValid_396;
  wire                _zz_s1_outputPayload_selValid_397;
  wire                _zz_s1_outputPayload_selValid_398;
  wire                _zz_s1_outputPayload_selValid_399;
  wire                _zz_s1_outputPayload_selValid_400;
  wire                _zz_s1_outputPayload_selValid_401;
  wire                _zz_s1_outputPayload_selValid_402;
  wire                _zz_s1_outputPayload_sel_12;
  wire                _zz_s1_outputPayload_sel_12_1;
  wire                _zz_s1_outputPayload_sel_12_2;
  wire                _zz_s1_outputPayload_sel_12_3;
  wire                _zz_s1_outputPayload_sel_12_4;
  wire                _zz_s1_outputPayload_selValid_403;
  wire                _zz_s1_outputPayload_selValid_404;
  wire                _zz_s1_outputPayload_selValid_405;
  wire                _zz_s1_outputPayload_selValid_406;
  wire                _zz_s1_outputPayload_selValid_407;
  wire                _zz_s1_outputPayload_selValid_408;
  wire                _zz_s1_outputPayload_selValid_409;
  wire                _zz_s1_outputPayload_selValid_410;
  wire                _zz_s1_outputPayload_selValid_411;
  wire                _zz_s1_outputPayload_selValid_412;
  wire                _zz_s1_outputPayload_selValid_413;
  wire                _zz_s1_outputPayload_selValid_414;
  wire                _zz_s1_outputPayload_selValid_415;
  wire                _zz_s1_outputPayload_selValid_416;
  wire                _zz_s1_outputPayload_selValid_417;
  wire                _zz_s1_outputPayload_selValid_418;
  wire                _zz_s1_outputPayload_selValid_419;
  wire                _zz_s1_outputPayload_selValid_420;
  wire                _zz_s1_outputPayload_selValid_421;
  wire                _zz_s1_outputPayload_selValid_422;
  wire                _zz_s1_outputPayload_selValid_423;
  wire                _zz_s1_outputPayload_selValid_424;
  wire                _zz_s1_outputPayload_selValid_425;
  wire                _zz_s1_outputPayload_selValid_426;
  wire                _zz_s1_outputPayload_selValid_427;
  wire                _zz_s1_outputPayload_selValid_428;
  wire                _zz_s1_outputPayload_selValid_429;
  wire                _zz_s1_outputPayload_selValid_430;
  wire                _zz_s1_outputPayload_selValid_431;
  wire                _zz_s1_outputPayload_selValid_432;
  wire                _zz_s1_outputPayload_selValid_433;
  wire                _zz_s1_outputPayload_sel_13;
  wire                _zz_s1_outputPayload_sel_13_1;
  wire                _zz_s1_outputPayload_sel_13_2;
  wire                _zz_s1_outputPayload_sel_13_3;
  wire                _zz_s1_outputPayload_sel_13_4;
  wire                _zz_s1_outputPayload_selValid_434;
  wire                _zz_s1_outputPayload_selValid_435;
  wire                _zz_s1_outputPayload_selValid_436;
  wire                _zz_s1_outputPayload_selValid_437;
  wire                _zz_s1_outputPayload_selValid_438;
  wire                _zz_s1_outputPayload_selValid_439;
  wire                _zz_s1_outputPayload_selValid_440;
  wire                _zz_s1_outputPayload_selValid_441;
  wire                _zz_s1_outputPayload_selValid_442;
  wire                _zz_s1_outputPayload_selValid_443;
  wire                _zz_s1_outputPayload_selValid_444;
  wire                _zz_s1_outputPayload_selValid_445;
  wire                _zz_s1_outputPayload_selValid_446;
  wire                _zz_s1_outputPayload_selValid_447;
  wire                _zz_s1_outputPayload_selValid_448;
  wire                _zz_s1_outputPayload_selValid_449;
  wire                _zz_s1_outputPayload_selValid_450;
  wire                _zz_s1_outputPayload_selValid_451;
  wire                _zz_s1_outputPayload_selValid_452;
  wire                _zz_s1_outputPayload_selValid_453;
  wire                _zz_s1_outputPayload_selValid_454;
  wire                _zz_s1_outputPayload_selValid_455;
  wire                _zz_s1_outputPayload_selValid_456;
  wire                _zz_s1_outputPayload_selValid_457;
  wire                _zz_s1_outputPayload_selValid_458;
  wire                _zz_s1_outputPayload_selValid_459;
  wire                _zz_s1_outputPayload_selValid_460;
  wire                _zz_s1_outputPayload_selValid_461;
  wire                _zz_s1_outputPayload_selValid_462;
  wire                _zz_s1_outputPayload_selValid_463;
  wire                _zz_s1_outputPayload_selValid_464;
  wire                _zz_s1_outputPayload_sel_14;
  wire                _zz_s1_outputPayload_sel_14_1;
  wire                _zz_s1_outputPayload_sel_14_2;
  wire                _zz_s1_outputPayload_sel_14_3;
  wire                _zz_s1_outputPayload_sel_14_4;
  wire                _zz_s1_outputPayload_selValid_465;
  wire                _zz_s1_outputPayload_selValid_466;
  wire                _zz_s1_outputPayload_selValid_467;
  wire                _zz_s1_outputPayload_selValid_468;
  wire                _zz_s1_outputPayload_selValid_469;
  wire                _zz_s1_outputPayload_selValid_470;
  wire                _zz_s1_outputPayload_selValid_471;
  wire                _zz_s1_outputPayload_selValid_472;
  wire                _zz_s1_outputPayload_selValid_473;
  wire                _zz_s1_outputPayload_selValid_474;
  wire                _zz_s1_outputPayload_selValid_475;
  wire                _zz_s1_outputPayload_selValid_476;
  wire                _zz_s1_outputPayload_selValid_477;
  wire                _zz_s1_outputPayload_selValid_478;
  wire                _zz_s1_outputPayload_selValid_479;
  wire                _zz_s1_outputPayload_selValid_480;
  wire                _zz_s1_outputPayload_selValid_481;
  wire                _zz_s1_outputPayload_selValid_482;
  wire                _zz_s1_outputPayload_selValid_483;
  wire                _zz_s1_outputPayload_selValid_484;
  wire                _zz_s1_outputPayload_selValid_485;
  wire                _zz_s1_outputPayload_selValid_486;
  wire                _zz_s1_outputPayload_selValid_487;
  wire                _zz_s1_outputPayload_selValid_488;
  wire                _zz_s1_outputPayload_selValid_489;
  wire                _zz_s1_outputPayload_selValid_490;
  wire                _zz_s1_outputPayload_selValid_491;
  wire                _zz_s1_outputPayload_selValid_492;
  wire                _zz_s1_outputPayload_selValid_493;
  wire                _zz_s1_outputPayload_selValid_494;
  wire                _zz_s1_outputPayload_selValid_495;
  wire                _zz_s1_outputPayload_sel_15;
  wire                _zz_s1_outputPayload_sel_15_1;
  wire                _zz_s1_outputPayload_sel_15_2;
  wire                _zz_s1_outputPayload_sel_15_3;
  wire                _zz_s1_outputPayload_sel_15_4;
  wire                _zz_s1_outputPayload_selValid_496;
  wire                _zz_s1_outputPayload_selValid_497;
  wire                _zz_s1_outputPayload_selValid_498;
  wire                _zz_s1_outputPayload_selValid_499;
  wire                _zz_s1_outputPayload_selValid_500;
  wire                _zz_s1_outputPayload_selValid_501;
  wire                _zz_s1_outputPayload_selValid_502;
  wire                _zz_s1_outputPayload_selValid_503;
  wire                _zz_s1_outputPayload_selValid_504;
  wire                _zz_s1_outputPayload_selValid_505;
  wire                _zz_s1_outputPayload_selValid_506;
  wire                _zz_s1_outputPayload_selValid_507;
  wire                _zz_s1_outputPayload_selValid_508;
  wire                _zz_s1_outputPayload_selValid_509;
  wire                _zz_s1_outputPayload_selValid_510;
  wire                _zz_s1_outputPayload_selValid_511;
  wire                _zz_s1_outputPayload_selValid_512;
  wire                _zz_s1_outputPayload_selValid_513;
  wire                _zz_s1_outputPayload_selValid_514;
  wire                _zz_s1_outputPayload_selValid_515;
  wire                _zz_s1_outputPayload_selValid_516;
  wire                _zz_s1_outputPayload_selValid_517;
  wire                _zz_s1_outputPayload_selValid_518;
  wire                _zz_s1_outputPayload_selValid_519;
  wire                _zz_s1_outputPayload_selValid_520;
  wire                _zz_s1_outputPayload_selValid_521;
  wire                _zz_s1_outputPayload_selValid_522;
  wire                _zz_s1_outputPayload_selValid_523;
  wire                _zz_s1_outputPayload_selValid_524;
  wire                _zz_s1_outputPayload_selValid_525;
  wire                _zz_s1_outputPayload_selValid_526;
  wire                _zz_s1_outputPayload_sel_16;
  wire                _zz_s1_outputPayload_sel_16_1;
  wire                _zz_s1_outputPayload_sel_16_2;
  wire                _zz_s1_outputPayload_sel_16_3;
  wire                _zz_s1_outputPayload_sel_16_4;
  wire                _zz_s1_outputPayload_selValid_527;
  wire                _zz_s1_outputPayload_selValid_528;
  wire                _zz_s1_outputPayload_selValid_529;
  wire                _zz_s1_outputPayload_selValid_530;
  wire                _zz_s1_outputPayload_selValid_531;
  wire                _zz_s1_outputPayload_selValid_532;
  wire                _zz_s1_outputPayload_selValid_533;
  wire                _zz_s1_outputPayload_selValid_534;
  wire                _zz_s1_outputPayload_selValid_535;
  wire                _zz_s1_outputPayload_selValid_536;
  wire                _zz_s1_outputPayload_selValid_537;
  wire                _zz_s1_outputPayload_selValid_538;
  wire                _zz_s1_outputPayload_selValid_539;
  wire                _zz_s1_outputPayload_selValid_540;
  wire                _zz_s1_outputPayload_selValid_541;
  wire                _zz_s1_outputPayload_selValid_542;
  wire                _zz_s1_outputPayload_selValid_543;
  wire                _zz_s1_outputPayload_selValid_544;
  wire                _zz_s1_outputPayload_selValid_545;
  wire                _zz_s1_outputPayload_selValid_546;
  wire                _zz_s1_outputPayload_selValid_547;
  wire                _zz_s1_outputPayload_selValid_548;
  wire                _zz_s1_outputPayload_selValid_549;
  wire                _zz_s1_outputPayload_selValid_550;
  wire                _zz_s1_outputPayload_selValid_551;
  wire                _zz_s1_outputPayload_selValid_552;
  wire                _zz_s1_outputPayload_selValid_553;
  wire                _zz_s1_outputPayload_selValid_554;
  wire                _zz_s1_outputPayload_selValid_555;
  wire                _zz_s1_outputPayload_selValid_556;
  wire                _zz_s1_outputPayload_selValid_557;
  wire                _zz_s1_outputPayload_sel_17;
  wire                _zz_s1_outputPayload_sel_17_1;
  wire                _zz_s1_outputPayload_sel_17_2;
  wire                _zz_s1_outputPayload_sel_17_3;
  wire                _zz_s1_outputPayload_sel_17_4;
  wire                _zz_s1_outputPayload_selValid_558;
  wire                _zz_s1_outputPayload_selValid_559;
  wire                _zz_s1_outputPayload_selValid_560;
  wire                _zz_s1_outputPayload_selValid_561;
  wire                _zz_s1_outputPayload_selValid_562;
  wire                _zz_s1_outputPayload_selValid_563;
  wire                _zz_s1_outputPayload_selValid_564;
  wire                _zz_s1_outputPayload_selValid_565;
  wire                _zz_s1_outputPayload_selValid_566;
  wire                _zz_s1_outputPayload_selValid_567;
  wire                _zz_s1_outputPayload_selValid_568;
  wire                _zz_s1_outputPayload_selValid_569;
  wire                _zz_s1_outputPayload_selValid_570;
  wire                _zz_s1_outputPayload_selValid_571;
  wire                _zz_s1_outputPayload_selValid_572;
  wire                _zz_s1_outputPayload_selValid_573;
  wire                _zz_s1_outputPayload_selValid_574;
  wire                _zz_s1_outputPayload_selValid_575;
  wire                _zz_s1_outputPayload_selValid_576;
  wire                _zz_s1_outputPayload_selValid_577;
  wire                _zz_s1_outputPayload_selValid_578;
  wire                _zz_s1_outputPayload_selValid_579;
  wire                _zz_s1_outputPayload_selValid_580;
  wire                _zz_s1_outputPayload_selValid_581;
  wire                _zz_s1_outputPayload_selValid_582;
  wire                _zz_s1_outputPayload_selValid_583;
  wire                _zz_s1_outputPayload_selValid_584;
  wire                _zz_s1_outputPayload_selValid_585;
  wire                _zz_s1_outputPayload_selValid_586;
  wire                _zz_s1_outputPayload_selValid_587;
  wire                _zz_s1_outputPayload_selValid_588;
  wire                _zz_s1_outputPayload_sel_18;
  wire                _zz_s1_outputPayload_sel_18_1;
  wire                _zz_s1_outputPayload_sel_18_2;
  wire                _zz_s1_outputPayload_sel_18_3;
  wire                _zz_s1_outputPayload_sel_18_4;
  wire                _zz_s1_outputPayload_selValid_589;
  wire                _zz_s1_outputPayload_selValid_590;
  wire                _zz_s1_outputPayload_selValid_591;
  wire                _zz_s1_outputPayload_selValid_592;
  wire                _zz_s1_outputPayload_selValid_593;
  wire                _zz_s1_outputPayload_selValid_594;
  wire                _zz_s1_outputPayload_selValid_595;
  wire                _zz_s1_outputPayload_selValid_596;
  wire                _zz_s1_outputPayload_selValid_597;
  wire                _zz_s1_outputPayload_selValid_598;
  wire                _zz_s1_outputPayload_selValid_599;
  wire                _zz_s1_outputPayload_selValid_600;
  wire                _zz_s1_outputPayload_selValid_601;
  wire                _zz_s1_outputPayload_selValid_602;
  wire                _zz_s1_outputPayload_selValid_603;
  wire                _zz_s1_outputPayload_selValid_604;
  wire                _zz_s1_outputPayload_selValid_605;
  wire                _zz_s1_outputPayload_selValid_606;
  wire                _zz_s1_outputPayload_selValid_607;
  wire                _zz_s1_outputPayload_selValid_608;
  wire                _zz_s1_outputPayload_selValid_609;
  wire                _zz_s1_outputPayload_selValid_610;
  wire                _zz_s1_outputPayload_selValid_611;
  wire                _zz_s1_outputPayload_selValid_612;
  wire                _zz_s1_outputPayload_selValid_613;
  wire                _zz_s1_outputPayload_selValid_614;
  wire                _zz_s1_outputPayload_selValid_615;
  wire                _zz_s1_outputPayload_selValid_616;
  wire                _zz_s1_outputPayload_selValid_617;
  wire                _zz_s1_outputPayload_selValid_618;
  wire                _zz_s1_outputPayload_selValid_619;
  wire                _zz_s1_outputPayload_sel_19;
  wire                _zz_s1_outputPayload_sel_19_1;
  wire                _zz_s1_outputPayload_sel_19_2;
  wire                _zz_s1_outputPayload_sel_19_3;
  wire                _zz_s1_outputPayload_sel_19_4;
  wire                _zz_s1_outputPayload_selValid_620;
  wire                _zz_s1_outputPayload_selValid_621;
  wire                _zz_s1_outputPayload_selValid_622;
  wire                _zz_s1_outputPayload_selValid_623;
  wire                _zz_s1_outputPayload_selValid_624;
  wire                _zz_s1_outputPayload_selValid_625;
  wire                _zz_s1_outputPayload_selValid_626;
  wire                _zz_s1_outputPayload_selValid_627;
  wire                _zz_s1_outputPayload_selValid_628;
  wire                _zz_s1_outputPayload_selValid_629;
  wire                _zz_s1_outputPayload_selValid_630;
  wire                _zz_s1_outputPayload_selValid_631;
  wire                _zz_s1_outputPayload_selValid_632;
  wire                _zz_s1_outputPayload_selValid_633;
  wire                _zz_s1_outputPayload_selValid_634;
  wire                _zz_s1_outputPayload_selValid_635;
  wire                _zz_s1_outputPayload_selValid_636;
  wire                _zz_s1_outputPayload_selValid_637;
  wire                _zz_s1_outputPayload_selValid_638;
  wire                _zz_s1_outputPayload_selValid_639;
  wire                _zz_s1_outputPayload_selValid_640;
  wire                _zz_s1_outputPayload_selValid_641;
  wire                _zz_s1_outputPayload_selValid_642;
  wire                _zz_s1_outputPayload_selValid_643;
  wire                _zz_s1_outputPayload_selValid_644;
  wire                _zz_s1_outputPayload_selValid_645;
  wire                _zz_s1_outputPayload_selValid_646;
  wire                _zz_s1_outputPayload_selValid_647;
  wire                _zz_s1_outputPayload_selValid_648;
  wire                _zz_s1_outputPayload_selValid_649;
  wire                _zz_s1_outputPayload_selValid_650;
  wire                _zz_s1_outputPayload_sel_20;
  wire                _zz_s1_outputPayload_sel_20_1;
  wire                _zz_s1_outputPayload_sel_20_2;
  wire                _zz_s1_outputPayload_sel_20_3;
  wire                _zz_s1_outputPayload_sel_20_4;
  wire                _zz_s1_outputPayload_selValid_651;
  wire                _zz_s1_outputPayload_selValid_652;
  wire                _zz_s1_outputPayload_selValid_653;
  wire                _zz_s1_outputPayload_selValid_654;
  wire                _zz_s1_outputPayload_selValid_655;
  wire                _zz_s1_outputPayload_selValid_656;
  wire                _zz_s1_outputPayload_selValid_657;
  wire                _zz_s1_outputPayload_selValid_658;
  wire                _zz_s1_outputPayload_selValid_659;
  wire                _zz_s1_outputPayload_selValid_660;
  wire                _zz_s1_outputPayload_selValid_661;
  wire                _zz_s1_outputPayload_selValid_662;
  wire                _zz_s1_outputPayload_selValid_663;
  wire                _zz_s1_outputPayload_selValid_664;
  wire                _zz_s1_outputPayload_selValid_665;
  wire                _zz_s1_outputPayload_selValid_666;
  wire                _zz_s1_outputPayload_selValid_667;
  wire                _zz_s1_outputPayload_selValid_668;
  wire                _zz_s1_outputPayload_selValid_669;
  wire                _zz_s1_outputPayload_selValid_670;
  wire                _zz_s1_outputPayload_selValid_671;
  wire                _zz_s1_outputPayload_selValid_672;
  wire                _zz_s1_outputPayload_selValid_673;
  wire                _zz_s1_outputPayload_selValid_674;
  wire                _zz_s1_outputPayload_selValid_675;
  wire                _zz_s1_outputPayload_selValid_676;
  wire                _zz_s1_outputPayload_selValid_677;
  wire                _zz_s1_outputPayload_selValid_678;
  wire                _zz_s1_outputPayload_selValid_679;
  wire                _zz_s1_outputPayload_selValid_680;
  wire                _zz_s1_outputPayload_selValid_681;
  wire                _zz_s1_outputPayload_sel_21;
  wire                _zz_s1_outputPayload_sel_21_1;
  wire                _zz_s1_outputPayload_sel_21_2;
  wire                _zz_s1_outputPayload_sel_21_3;
  wire                _zz_s1_outputPayload_sel_21_4;
  wire                _zz_s1_outputPayload_selValid_682;
  wire                _zz_s1_outputPayload_selValid_683;
  wire                _zz_s1_outputPayload_selValid_684;
  wire                _zz_s1_outputPayload_selValid_685;
  wire                _zz_s1_outputPayload_selValid_686;
  wire                _zz_s1_outputPayload_selValid_687;
  wire                _zz_s1_outputPayload_selValid_688;
  wire                _zz_s1_outputPayload_selValid_689;
  wire                _zz_s1_outputPayload_selValid_690;
  wire                _zz_s1_outputPayload_selValid_691;
  wire                _zz_s1_outputPayload_selValid_692;
  wire                _zz_s1_outputPayload_selValid_693;
  wire                _zz_s1_outputPayload_selValid_694;
  wire                _zz_s1_outputPayload_selValid_695;
  wire                _zz_s1_outputPayload_selValid_696;
  wire                _zz_s1_outputPayload_selValid_697;
  wire                _zz_s1_outputPayload_selValid_698;
  wire                _zz_s1_outputPayload_selValid_699;
  wire                _zz_s1_outputPayload_selValid_700;
  wire                _zz_s1_outputPayload_selValid_701;
  wire                _zz_s1_outputPayload_selValid_702;
  wire                _zz_s1_outputPayload_selValid_703;
  wire                _zz_s1_outputPayload_selValid_704;
  wire                _zz_s1_outputPayload_selValid_705;
  wire                _zz_s1_outputPayload_selValid_706;
  wire                _zz_s1_outputPayload_selValid_707;
  wire                _zz_s1_outputPayload_selValid_708;
  wire                _zz_s1_outputPayload_selValid_709;
  wire                _zz_s1_outputPayload_selValid_710;
  wire                _zz_s1_outputPayload_selValid_711;
  wire                _zz_s1_outputPayload_selValid_712;
  wire                _zz_s1_outputPayload_sel_22;
  wire                _zz_s1_outputPayload_sel_22_1;
  wire                _zz_s1_outputPayload_sel_22_2;
  wire                _zz_s1_outputPayload_sel_22_3;
  wire                _zz_s1_outputPayload_sel_22_4;
  wire                _zz_s1_outputPayload_selValid_713;
  wire                _zz_s1_outputPayload_selValid_714;
  wire                _zz_s1_outputPayload_selValid_715;
  wire                _zz_s1_outputPayload_selValid_716;
  wire                _zz_s1_outputPayload_selValid_717;
  wire                _zz_s1_outputPayload_selValid_718;
  wire                _zz_s1_outputPayload_selValid_719;
  wire                _zz_s1_outputPayload_selValid_720;
  wire                _zz_s1_outputPayload_selValid_721;
  wire                _zz_s1_outputPayload_selValid_722;
  wire                _zz_s1_outputPayload_selValid_723;
  wire                _zz_s1_outputPayload_selValid_724;
  wire                _zz_s1_outputPayload_selValid_725;
  wire                _zz_s1_outputPayload_selValid_726;
  wire                _zz_s1_outputPayload_selValid_727;
  wire                _zz_s1_outputPayload_selValid_728;
  wire                _zz_s1_outputPayload_selValid_729;
  wire                _zz_s1_outputPayload_selValid_730;
  wire                _zz_s1_outputPayload_selValid_731;
  wire                _zz_s1_outputPayload_selValid_732;
  wire                _zz_s1_outputPayload_selValid_733;
  wire                _zz_s1_outputPayload_selValid_734;
  wire                _zz_s1_outputPayload_selValid_735;
  wire                _zz_s1_outputPayload_selValid_736;
  wire                _zz_s1_outputPayload_selValid_737;
  wire                _zz_s1_outputPayload_selValid_738;
  wire                _zz_s1_outputPayload_selValid_739;
  wire                _zz_s1_outputPayload_selValid_740;
  wire                _zz_s1_outputPayload_selValid_741;
  wire                _zz_s1_outputPayload_selValid_742;
  wire                _zz_s1_outputPayload_selValid_743;
  wire                _zz_s1_outputPayload_sel_23;
  wire                _zz_s1_outputPayload_sel_23_1;
  wire                _zz_s1_outputPayload_sel_23_2;
  wire                _zz_s1_outputPayload_sel_23_3;
  wire                _zz_s1_outputPayload_sel_23_4;
  wire                _zz_s1_outputPayload_selValid_744;
  wire                _zz_s1_outputPayload_selValid_745;
  wire                _zz_s1_outputPayload_selValid_746;
  wire                _zz_s1_outputPayload_selValid_747;
  wire                _zz_s1_outputPayload_selValid_748;
  wire                _zz_s1_outputPayload_selValid_749;
  wire                _zz_s1_outputPayload_selValid_750;
  wire                _zz_s1_outputPayload_selValid_751;
  wire                _zz_s1_outputPayload_selValid_752;
  wire                _zz_s1_outputPayload_selValid_753;
  wire                _zz_s1_outputPayload_selValid_754;
  wire                _zz_s1_outputPayload_selValid_755;
  wire                _zz_s1_outputPayload_selValid_756;
  wire                _zz_s1_outputPayload_selValid_757;
  wire                _zz_s1_outputPayload_selValid_758;
  wire                _zz_s1_outputPayload_selValid_759;
  wire                _zz_s1_outputPayload_selValid_760;
  wire                _zz_s1_outputPayload_selValid_761;
  wire                _zz_s1_outputPayload_selValid_762;
  wire                _zz_s1_outputPayload_selValid_763;
  wire                _zz_s1_outputPayload_selValid_764;
  wire                _zz_s1_outputPayload_selValid_765;
  wire                _zz_s1_outputPayload_selValid_766;
  wire                _zz_s1_outputPayload_selValid_767;
  wire                _zz_s1_outputPayload_selValid_768;
  wire                _zz_s1_outputPayload_selValid_769;
  wire                _zz_s1_outputPayload_selValid_770;
  wire                _zz_s1_outputPayload_selValid_771;
  wire                _zz_s1_outputPayload_selValid_772;
  wire                _zz_s1_outputPayload_selValid_773;
  wire                _zz_s1_outputPayload_selValid_774;
  wire                _zz_s1_outputPayload_sel_24;
  wire                _zz_s1_outputPayload_sel_24_1;
  wire                _zz_s1_outputPayload_sel_24_2;
  wire                _zz_s1_outputPayload_sel_24_3;
  wire                _zz_s1_outputPayload_sel_24_4;
  wire                _zz_s1_outputPayload_selValid_775;
  wire                _zz_s1_outputPayload_selValid_776;
  wire                _zz_s1_outputPayload_selValid_777;
  wire                _zz_s1_outputPayload_selValid_778;
  wire                _zz_s1_outputPayload_selValid_779;
  wire                _zz_s1_outputPayload_selValid_780;
  wire                _zz_s1_outputPayload_selValid_781;
  wire                _zz_s1_outputPayload_selValid_782;
  wire                _zz_s1_outputPayload_selValid_783;
  wire                _zz_s1_outputPayload_selValid_784;
  wire                _zz_s1_outputPayload_selValid_785;
  wire                _zz_s1_outputPayload_selValid_786;
  wire                _zz_s1_outputPayload_selValid_787;
  wire                _zz_s1_outputPayload_selValid_788;
  wire                _zz_s1_outputPayload_selValid_789;
  wire                _zz_s1_outputPayload_selValid_790;
  wire                _zz_s1_outputPayload_selValid_791;
  wire                _zz_s1_outputPayload_selValid_792;
  wire                _zz_s1_outputPayload_selValid_793;
  wire                _zz_s1_outputPayload_selValid_794;
  wire                _zz_s1_outputPayload_selValid_795;
  wire                _zz_s1_outputPayload_selValid_796;
  wire                _zz_s1_outputPayload_selValid_797;
  wire                _zz_s1_outputPayload_selValid_798;
  wire                _zz_s1_outputPayload_selValid_799;
  wire                _zz_s1_outputPayload_selValid_800;
  wire                _zz_s1_outputPayload_selValid_801;
  wire                _zz_s1_outputPayload_selValid_802;
  wire                _zz_s1_outputPayload_selValid_803;
  wire                _zz_s1_outputPayload_selValid_804;
  wire                _zz_s1_outputPayload_selValid_805;
  wire                _zz_s1_outputPayload_sel_25;
  wire                _zz_s1_outputPayload_sel_25_1;
  wire                _zz_s1_outputPayload_sel_25_2;
  wire                _zz_s1_outputPayload_sel_25_3;
  wire                _zz_s1_outputPayload_sel_25_4;
  wire                _zz_s1_outputPayload_selValid_806;
  wire                _zz_s1_outputPayload_selValid_807;
  wire                _zz_s1_outputPayload_selValid_808;
  wire                _zz_s1_outputPayload_selValid_809;
  wire                _zz_s1_outputPayload_selValid_810;
  wire                _zz_s1_outputPayload_selValid_811;
  wire                _zz_s1_outputPayload_selValid_812;
  wire                _zz_s1_outputPayload_selValid_813;
  wire                _zz_s1_outputPayload_selValid_814;
  wire                _zz_s1_outputPayload_selValid_815;
  wire                _zz_s1_outputPayload_selValid_816;
  wire                _zz_s1_outputPayload_selValid_817;
  wire                _zz_s1_outputPayload_selValid_818;
  wire                _zz_s1_outputPayload_selValid_819;
  wire                _zz_s1_outputPayload_selValid_820;
  wire                _zz_s1_outputPayload_selValid_821;
  wire                _zz_s1_outputPayload_selValid_822;
  wire                _zz_s1_outputPayload_selValid_823;
  wire                _zz_s1_outputPayload_selValid_824;
  wire                _zz_s1_outputPayload_selValid_825;
  wire                _zz_s1_outputPayload_selValid_826;
  wire                _zz_s1_outputPayload_selValid_827;
  wire                _zz_s1_outputPayload_selValid_828;
  wire                _zz_s1_outputPayload_selValid_829;
  wire                _zz_s1_outputPayload_selValid_830;
  wire                _zz_s1_outputPayload_selValid_831;
  wire                _zz_s1_outputPayload_selValid_832;
  wire                _zz_s1_outputPayload_selValid_833;
  wire                _zz_s1_outputPayload_selValid_834;
  wire                _zz_s1_outputPayload_selValid_835;
  wire                _zz_s1_outputPayload_selValid_836;
  wire                _zz_s1_outputPayload_sel_26;
  wire                _zz_s1_outputPayload_sel_26_1;
  wire                _zz_s1_outputPayload_sel_26_2;
  wire                _zz_s1_outputPayload_sel_26_3;
  wire                _zz_s1_outputPayload_sel_26_4;
  wire                _zz_s1_outputPayload_selValid_837;
  wire                _zz_s1_outputPayload_selValid_838;
  wire                _zz_s1_outputPayload_selValid_839;
  wire                _zz_s1_outputPayload_selValid_840;
  wire                _zz_s1_outputPayload_selValid_841;
  wire                _zz_s1_outputPayload_selValid_842;
  wire                _zz_s1_outputPayload_selValid_843;
  wire                _zz_s1_outputPayload_selValid_844;
  wire                _zz_s1_outputPayload_selValid_845;
  wire                _zz_s1_outputPayload_selValid_846;
  wire                _zz_s1_outputPayload_selValid_847;
  wire                _zz_s1_outputPayload_selValid_848;
  wire                _zz_s1_outputPayload_selValid_849;
  wire                _zz_s1_outputPayload_selValid_850;
  wire                _zz_s1_outputPayload_selValid_851;
  wire                _zz_s1_outputPayload_selValid_852;
  wire                _zz_s1_outputPayload_selValid_853;
  wire                _zz_s1_outputPayload_selValid_854;
  wire                _zz_s1_outputPayload_selValid_855;
  wire                _zz_s1_outputPayload_selValid_856;
  wire                _zz_s1_outputPayload_selValid_857;
  wire                _zz_s1_outputPayload_selValid_858;
  wire                _zz_s1_outputPayload_selValid_859;
  wire                _zz_s1_outputPayload_selValid_860;
  wire                _zz_s1_outputPayload_selValid_861;
  wire                _zz_s1_outputPayload_selValid_862;
  wire                _zz_s1_outputPayload_selValid_863;
  wire                _zz_s1_outputPayload_selValid_864;
  wire                _zz_s1_outputPayload_selValid_865;
  wire                _zz_s1_outputPayload_selValid_866;
  wire                _zz_s1_outputPayload_selValid_867;
  wire                _zz_s1_outputPayload_sel_27;
  wire                _zz_s1_outputPayload_sel_27_1;
  wire                _zz_s1_outputPayload_sel_27_2;
  wire                _zz_s1_outputPayload_sel_27_3;
  wire                _zz_s1_outputPayload_sel_27_4;
  wire                _zz_s1_outputPayload_selValid_868;
  wire                _zz_s1_outputPayload_selValid_869;
  wire                _zz_s1_outputPayload_selValid_870;
  wire                _zz_s1_outputPayload_selValid_871;
  wire                _zz_s1_outputPayload_selValid_872;
  wire                _zz_s1_outputPayload_selValid_873;
  wire                _zz_s1_outputPayload_selValid_874;
  wire                _zz_s1_outputPayload_selValid_875;
  wire                _zz_s1_outputPayload_selValid_876;
  wire                _zz_s1_outputPayload_selValid_877;
  wire                _zz_s1_outputPayload_selValid_878;
  wire                _zz_s1_outputPayload_selValid_879;
  wire                _zz_s1_outputPayload_selValid_880;
  wire                _zz_s1_outputPayload_selValid_881;
  wire                _zz_s1_outputPayload_selValid_882;
  wire                _zz_s1_outputPayload_selValid_883;
  wire                _zz_s1_outputPayload_selValid_884;
  wire                _zz_s1_outputPayload_selValid_885;
  wire                _zz_s1_outputPayload_selValid_886;
  wire                _zz_s1_outputPayload_selValid_887;
  wire                _zz_s1_outputPayload_selValid_888;
  wire                _zz_s1_outputPayload_selValid_889;
  wire                _zz_s1_outputPayload_selValid_890;
  wire                _zz_s1_outputPayload_selValid_891;
  wire                _zz_s1_outputPayload_selValid_892;
  wire                _zz_s1_outputPayload_selValid_893;
  wire                _zz_s1_outputPayload_selValid_894;
  wire                _zz_s1_outputPayload_selValid_895;
  wire                _zz_s1_outputPayload_selValid_896;
  wire                _zz_s1_outputPayload_selValid_897;
  wire                _zz_s1_outputPayload_selValid_898;
  wire                _zz_s1_outputPayload_sel_28;
  wire                _zz_s1_outputPayload_sel_28_1;
  wire                _zz_s1_outputPayload_sel_28_2;
  wire                _zz_s1_outputPayload_sel_28_3;
  wire                _zz_s1_outputPayload_sel_28_4;
  wire                _zz_s1_outputPayload_selValid_899;
  wire                _zz_s1_outputPayload_selValid_900;
  wire                _zz_s1_outputPayload_selValid_901;
  wire                _zz_s1_outputPayload_selValid_902;
  wire                _zz_s1_outputPayload_selValid_903;
  wire                _zz_s1_outputPayload_selValid_904;
  wire                _zz_s1_outputPayload_selValid_905;
  wire                _zz_s1_outputPayload_selValid_906;
  wire                _zz_s1_outputPayload_selValid_907;
  wire                _zz_s1_outputPayload_selValid_908;
  wire                _zz_s1_outputPayload_selValid_909;
  wire                _zz_s1_outputPayload_selValid_910;
  wire                _zz_s1_outputPayload_selValid_911;
  wire                _zz_s1_outputPayload_selValid_912;
  wire                _zz_s1_outputPayload_selValid_913;
  wire                _zz_s1_outputPayload_selValid_914;
  wire                _zz_s1_outputPayload_selValid_915;
  wire                _zz_s1_outputPayload_selValid_916;
  wire                _zz_s1_outputPayload_selValid_917;
  wire                _zz_s1_outputPayload_selValid_918;
  wire                _zz_s1_outputPayload_selValid_919;
  wire                _zz_s1_outputPayload_selValid_920;
  wire                _zz_s1_outputPayload_selValid_921;
  wire                _zz_s1_outputPayload_selValid_922;
  wire                _zz_s1_outputPayload_selValid_923;
  wire                _zz_s1_outputPayload_selValid_924;
  wire                _zz_s1_outputPayload_selValid_925;
  wire                _zz_s1_outputPayload_selValid_926;
  wire                _zz_s1_outputPayload_selValid_927;
  wire                _zz_s1_outputPayload_selValid_928;
  wire                _zz_s1_outputPayload_selValid_929;
  wire                _zz_s1_outputPayload_sel_29;
  wire                _zz_s1_outputPayload_sel_29_1;
  wire                _zz_s1_outputPayload_sel_29_2;
  wire                _zz_s1_outputPayload_sel_29_3;
  wire                _zz_s1_outputPayload_sel_29_4;
  wire                _zz_s1_outputPayload_selValid_930;
  wire                _zz_s1_outputPayload_selValid_931;
  wire                _zz_s1_outputPayload_selValid_932;
  wire                _zz_s1_outputPayload_selValid_933;
  wire                _zz_s1_outputPayload_selValid_934;
  wire                _zz_s1_outputPayload_selValid_935;
  wire                _zz_s1_outputPayload_selValid_936;
  wire                _zz_s1_outputPayload_selValid_937;
  wire                _zz_s1_outputPayload_selValid_938;
  wire                _zz_s1_outputPayload_selValid_939;
  wire                _zz_s1_outputPayload_selValid_940;
  wire                _zz_s1_outputPayload_selValid_941;
  wire                _zz_s1_outputPayload_selValid_942;
  wire                _zz_s1_outputPayload_selValid_943;
  wire                _zz_s1_outputPayload_selValid_944;
  wire                _zz_s1_outputPayload_selValid_945;
  wire                _zz_s1_outputPayload_selValid_946;
  wire                _zz_s1_outputPayload_selValid_947;
  wire                _zz_s1_outputPayload_selValid_948;
  wire                _zz_s1_outputPayload_selValid_949;
  wire                _zz_s1_outputPayload_selValid_950;
  wire                _zz_s1_outputPayload_selValid_951;
  wire                _zz_s1_outputPayload_selValid_952;
  wire                _zz_s1_outputPayload_selValid_953;
  wire                _zz_s1_outputPayload_selValid_954;
  wire                _zz_s1_outputPayload_selValid_955;
  wire                _zz_s1_outputPayload_selValid_956;
  wire                _zz_s1_outputPayload_selValid_957;
  wire                _zz_s1_outputPayload_selValid_958;
  wire                _zz_s1_outputPayload_selValid_959;
  wire                _zz_s1_outputPayload_selValid_960;
  wire                _zz_s1_outputPayload_sel_30;
  wire                _zz_s1_outputPayload_sel_30_1;
  wire                _zz_s1_outputPayload_sel_30_2;
  wire                _zz_s1_outputPayload_sel_30_3;
  wire                _zz_s1_outputPayload_sel_30_4;
  wire                _zz_s1_outputPayload_selValid_961;
  wire                _zz_s1_outputPayload_selValid_962;
  wire                _zz_s1_outputPayload_selValid_963;
  wire                _zz_s1_outputPayload_selValid_964;
  wire                _zz_s1_outputPayload_selValid_965;
  wire                _zz_s1_outputPayload_selValid_966;
  wire                _zz_s1_outputPayload_selValid_967;
  wire                _zz_s1_outputPayload_selValid_968;
  wire                _zz_s1_outputPayload_selValid_969;
  wire                _zz_s1_outputPayload_selValid_970;
  wire                _zz_s1_outputPayload_selValid_971;
  wire                _zz_s1_outputPayload_selValid_972;
  wire                _zz_s1_outputPayload_selValid_973;
  wire                _zz_s1_outputPayload_selValid_974;
  wire                _zz_s1_outputPayload_selValid_975;
  wire                _zz_s1_outputPayload_selValid_976;
  wire                _zz_s1_outputPayload_selValid_977;
  wire                _zz_s1_outputPayload_selValid_978;
  wire                _zz_s1_outputPayload_selValid_979;
  wire                _zz_s1_outputPayload_selValid_980;
  wire                _zz_s1_outputPayload_selValid_981;
  wire                _zz_s1_outputPayload_selValid_982;
  wire                _zz_s1_outputPayload_selValid_983;
  wire                _zz_s1_outputPayload_selValid_984;
  wire                _zz_s1_outputPayload_selValid_985;
  wire                _zz_s1_outputPayload_selValid_986;
  wire                _zz_s1_outputPayload_selValid_987;
  wire                _zz_s1_outputPayload_selValid_988;
  wire                _zz_s1_outputPayload_selValid_989;
  wire                _zz_s1_outputPayload_selValid_990;
  wire                _zz_s1_outputPayload_selValid_991;
  wire                _zz_s1_outputPayload_sel_31;
  wire                _zz_s1_outputPayload_sel_31_1;
  wire                _zz_s1_outputPayload_sel_31_2;
  wire                _zz_s1_outputPayload_sel_31_3;
  wire                _zz_s1_outputPayload_sel_31_4;
  wire                s1_output_valid;
  reg                 s1_output_ready;
  wire       [255:0]  s1_output_payload_cmd_data;
  wire       [31:0]   s1_output_payload_cmd_mask;
  wire       [4:0]    s1_output_payload_index_0;
  wire       [4:0]    s1_output_payload_index_1;
  wire       [4:0]    s1_output_payload_index_2;
  wire       [4:0]    s1_output_payload_index_3;
  wire       [4:0]    s1_output_payload_index_4;
  wire       [4:0]    s1_output_payload_index_5;
  wire       [4:0]    s1_output_payload_index_6;
  wire       [4:0]    s1_output_payload_index_7;
  wire       [4:0]    s1_output_payload_index_8;
  wire       [4:0]    s1_output_payload_index_9;
  wire       [4:0]    s1_output_payload_index_10;
  wire       [4:0]    s1_output_payload_index_11;
  wire       [4:0]    s1_output_payload_index_12;
  wire       [4:0]    s1_output_payload_index_13;
  wire       [4:0]    s1_output_payload_index_14;
  wire       [4:0]    s1_output_payload_index_15;
  wire       [4:0]    s1_output_payload_index_16;
  wire       [4:0]    s1_output_payload_index_17;
  wire       [4:0]    s1_output_payload_index_18;
  wire       [4:0]    s1_output_payload_index_19;
  wire       [4:0]    s1_output_payload_index_20;
  wire       [4:0]    s1_output_payload_index_21;
  wire       [4:0]    s1_output_payload_index_22;
  wire       [4:0]    s1_output_payload_index_23;
  wire       [4:0]    s1_output_payload_index_24;
  wire       [4:0]    s1_output_payload_index_25;
  wire       [4:0]    s1_output_payload_index_26;
  wire       [4:0]    s1_output_payload_index_27;
  wire       [4:0]    s1_output_payload_index_28;
  wire       [4:0]    s1_output_payload_index_29;
  wire       [4:0]    s1_output_payload_index_30;
  wire       [4:0]    s1_output_payload_index_31;
  wire                s1_output_payload_last;
  wire       [4:0]    s1_output_payload_sel_0;
  wire       [4:0]    s1_output_payload_sel_1;
  wire       [4:0]    s1_output_payload_sel_2;
  wire       [4:0]    s1_output_payload_sel_3;
  wire       [4:0]    s1_output_payload_sel_4;
  wire       [4:0]    s1_output_payload_sel_5;
  wire       [4:0]    s1_output_payload_sel_6;
  wire       [4:0]    s1_output_payload_sel_7;
  wire       [4:0]    s1_output_payload_sel_8;
  wire       [4:0]    s1_output_payload_sel_9;
  wire       [4:0]    s1_output_payload_sel_10;
  wire       [4:0]    s1_output_payload_sel_11;
  wire       [4:0]    s1_output_payload_sel_12;
  wire       [4:0]    s1_output_payload_sel_13;
  wire       [4:0]    s1_output_payload_sel_14;
  wire       [4:0]    s1_output_payload_sel_15;
  wire       [4:0]    s1_output_payload_sel_16;
  wire       [4:0]    s1_output_payload_sel_17;
  wire       [4:0]    s1_output_payload_sel_18;
  wire       [4:0]    s1_output_payload_sel_19;
  wire       [4:0]    s1_output_payload_sel_20;
  wire       [4:0]    s1_output_payload_sel_21;
  wire       [4:0]    s1_output_payload_sel_22;
  wire       [4:0]    s1_output_payload_sel_23;
  wire       [4:0]    s1_output_payload_sel_24;
  wire       [4:0]    s1_output_payload_sel_25;
  wire       [4:0]    s1_output_payload_sel_26;
  wire       [4:0]    s1_output_payload_sel_27;
  wire       [4:0]    s1_output_payload_sel_28;
  wire       [4:0]    s1_output_payload_sel_29;
  wire       [4:0]    s1_output_payload_sel_30;
  wire       [4:0]    s1_output_payload_sel_31;
  wire       [31:0]   s1_output_payload_selValid;
  wire                s2_input_valid;
  reg                 s2_input_ready;
  wire       [255:0]  s2_input_payload_cmd_data;
  wire       [31:0]   s2_input_payload_cmd_mask;
  wire       [4:0]    s2_input_payload_index_0;
  wire       [4:0]    s2_input_payload_index_1;
  wire       [4:0]    s2_input_payload_index_2;
  wire       [4:0]    s2_input_payload_index_3;
  wire       [4:0]    s2_input_payload_index_4;
  wire       [4:0]    s2_input_payload_index_5;
  wire       [4:0]    s2_input_payload_index_6;
  wire       [4:0]    s2_input_payload_index_7;
  wire       [4:0]    s2_input_payload_index_8;
  wire       [4:0]    s2_input_payload_index_9;
  wire       [4:0]    s2_input_payload_index_10;
  wire       [4:0]    s2_input_payload_index_11;
  wire       [4:0]    s2_input_payload_index_12;
  wire       [4:0]    s2_input_payload_index_13;
  wire       [4:0]    s2_input_payload_index_14;
  wire       [4:0]    s2_input_payload_index_15;
  wire       [4:0]    s2_input_payload_index_16;
  wire       [4:0]    s2_input_payload_index_17;
  wire       [4:0]    s2_input_payload_index_18;
  wire       [4:0]    s2_input_payload_index_19;
  wire       [4:0]    s2_input_payload_index_20;
  wire       [4:0]    s2_input_payload_index_21;
  wire       [4:0]    s2_input_payload_index_22;
  wire       [4:0]    s2_input_payload_index_23;
  wire       [4:0]    s2_input_payload_index_24;
  wire       [4:0]    s2_input_payload_index_25;
  wire       [4:0]    s2_input_payload_index_26;
  wire       [4:0]    s2_input_payload_index_27;
  wire       [4:0]    s2_input_payload_index_28;
  wire       [4:0]    s2_input_payload_index_29;
  wire       [4:0]    s2_input_payload_index_30;
  wire       [4:0]    s2_input_payload_index_31;
  wire                s2_input_payload_last;
  wire       [4:0]    s2_input_payload_sel_0;
  wire       [4:0]    s2_input_payload_sel_1;
  wire       [4:0]    s2_input_payload_sel_2;
  wire       [4:0]    s2_input_payload_sel_3;
  wire       [4:0]    s2_input_payload_sel_4;
  wire       [4:0]    s2_input_payload_sel_5;
  wire       [4:0]    s2_input_payload_sel_6;
  wire       [4:0]    s2_input_payload_sel_7;
  wire       [4:0]    s2_input_payload_sel_8;
  wire       [4:0]    s2_input_payload_sel_9;
  wire       [4:0]    s2_input_payload_sel_10;
  wire       [4:0]    s2_input_payload_sel_11;
  wire       [4:0]    s2_input_payload_sel_12;
  wire       [4:0]    s2_input_payload_sel_13;
  wire       [4:0]    s2_input_payload_sel_14;
  wire       [4:0]    s2_input_payload_sel_15;
  wire       [4:0]    s2_input_payload_sel_16;
  wire       [4:0]    s2_input_payload_sel_17;
  wire       [4:0]    s2_input_payload_sel_18;
  wire       [4:0]    s2_input_payload_sel_19;
  wire       [4:0]    s2_input_payload_sel_20;
  wire       [4:0]    s2_input_payload_sel_21;
  wire       [4:0]    s2_input_payload_sel_22;
  wire       [4:0]    s2_input_payload_sel_23;
  wire       [4:0]    s2_input_payload_sel_24;
  wire       [4:0]    s2_input_payload_sel_25;
  wire       [4:0]    s2_input_payload_sel_26;
  wire       [4:0]    s2_input_payload_sel_27;
  wire       [4:0]    s2_input_payload_sel_28;
  wire       [4:0]    s2_input_payload_sel_29;
  wire       [4:0]    s2_input_payload_sel_30;
  wire       [4:0]    s2_input_payload_sel_31;
  wire       [31:0]   s2_input_payload_selValid;
  reg                 s1_output_rValid;
  reg        [255:0]  s1_output_rData_cmd_data;
  reg        [31:0]   s1_output_rData_cmd_mask;
  reg        [4:0]    s1_output_rData_index_0;
  reg        [4:0]    s1_output_rData_index_1;
  reg        [4:0]    s1_output_rData_index_2;
  reg        [4:0]    s1_output_rData_index_3;
  reg        [4:0]    s1_output_rData_index_4;
  reg        [4:0]    s1_output_rData_index_5;
  reg        [4:0]    s1_output_rData_index_6;
  reg        [4:0]    s1_output_rData_index_7;
  reg        [4:0]    s1_output_rData_index_8;
  reg        [4:0]    s1_output_rData_index_9;
  reg        [4:0]    s1_output_rData_index_10;
  reg        [4:0]    s1_output_rData_index_11;
  reg        [4:0]    s1_output_rData_index_12;
  reg        [4:0]    s1_output_rData_index_13;
  reg        [4:0]    s1_output_rData_index_14;
  reg        [4:0]    s1_output_rData_index_15;
  reg        [4:0]    s1_output_rData_index_16;
  reg        [4:0]    s1_output_rData_index_17;
  reg        [4:0]    s1_output_rData_index_18;
  reg        [4:0]    s1_output_rData_index_19;
  reg        [4:0]    s1_output_rData_index_20;
  reg        [4:0]    s1_output_rData_index_21;
  reg        [4:0]    s1_output_rData_index_22;
  reg        [4:0]    s1_output_rData_index_23;
  reg        [4:0]    s1_output_rData_index_24;
  reg        [4:0]    s1_output_rData_index_25;
  reg        [4:0]    s1_output_rData_index_26;
  reg        [4:0]    s1_output_rData_index_27;
  reg        [4:0]    s1_output_rData_index_28;
  reg        [4:0]    s1_output_rData_index_29;
  reg        [4:0]    s1_output_rData_index_30;
  reg        [4:0]    s1_output_rData_index_31;
  reg                 s1_output_rData_last;
  reg        [4:0]    s1_output_rData_sel_0;
  reg        [4:0]    s1_output_rData_sel_1;
  reg        [4:0]    s1_output_rData_sel_2;
  reg        [4:0]    s1_output_rData_sel_3;
  reg        [4:0]    s1_output_rData_sel_4;
  reg        [4:0]    s1_output_rData_sel_5;
  reg        [4:0]    s1_output_rData_sel_6;
  reg        [4:0]    s1_output_rData_sel_7;
  reg        [4:0]    s1_output_rData_sel_8;
  reg        [4:0]    s1_output_rData_sel_9;
  reg        [4:0]    s1_output_rData_sel_10;
  reg        [4:0]    s1_output_rData_sel_11;
  reg        [4:0]    s1_output_rData_sel_12;
  reg        [4:0]    s1_output_rData_sel_13;
  reg        [4:0]    s1_output_rData_sel_14;
  reg        [4:0]    s1_output_rData_sel_15;
  reg        [4:0]    s1_output_rData_sel_16;
  reg        [4:0]    s1_output_rData_sel_17;
  reg        [4:0]    s1_output_rData_sel_18;
  reg        [4:0]    s1_output_rData_sel_19;
  reg        [4:0]    s1_output_rData_sel_20;
  reg        [4:0]    s1_output_rData_sel_21;
  reg        [4:0]    s1_output_rData_sel_22;
  reg        [4:0]    s1_output_rData_sel_23;
  reg        [4:0]    s1_output_rData_sel_24;
  reg        [4:0]    s1_output_rData_sel_25;
  reg        [4:0]    s1_output_rData_sel_26;
  reg        [4:0]    s1_output_rData_sel_27;
  reg        [4:0]    s1_output_rData_sel_28;
  reg        [4:0]    s1_output_rData_sel_29;
  reg        [4:0]    s1_output_rData_sel_30;
  reg        [4:0]    s1_output_rData_sel_31;
  reg        [31:0]   s1_output_rData_selValid;
  wire                when_Stream_l375_2;
  wire                when_DmaSg_l1464;
  wire                s2_input_fire;
  wire       [7:0]    s2_inputDataBytes_0;
  wire       [7:0]    s2_inputDataBytes_1;
  wire       [7:0]    s2_inputDataBytes_2;
  wire       [7:0]    s2_inputDataBytes_3;
  wire       [7:0]    s2_inputDataBytes_4;
  wire       [7:0]    s2_inputDataBytes_5;
  wire       [7:0]    s2_inputDataBytes_6;
  wire       [7:0]    s2_inputDataBytes_7;
  wire       [7:0]    s2_inputDataBytes_8;
  wire       [7:0]    s2_inputDataBytes_9;
  wire       [7:0]    s2_inputDataBytes_10;
  wire       [7:0]    s2_inputDataBytes_11;
  wire       [7:0]    s2_inputDataBytes_12;
  wire       [7:0]    s2_inputDataBytes_13;
  wire       [7:0]    s2_inputDataBytes_14;
  wire       [7:0]    s2_inputDataBytes_15;
  wire       [7:0]    s2_inputDataBytes_16;
  wire       [7:0]    s2_inputDataBytes_17;
  wire       [7:0]    s2_inputDataBytes_18;
  wire       [7:0]    s2_inputDataBytes_19;
  wire       [7:0]    s2_inputDataBytes_20;
  wire       [7:0]    s2_inputDataBytes_21;
  wire       [7:0]    s2_inputDataBytes_22;
  wire       [7:0]    s2_inputDataBytes_23;
  wire       [7:0]    s2_inputDataBytes_24;
  wire       [7:0]    s2_inputDataBytes_25;
  wire       [7:0]    s2_inputDataBytes_26;
  wire       [7:0]    s2_inputDataBytes_27;
  wire       [7:0]    s2_inputDataBytes_28;
  wire       [7:0]    s2_inputDataBytes_29;
  wire       [7:0]    s2_inputDataBytes_30;
  wire       [7:0]    s2_inputDataBytes_31;
  reg                 s2_byteLogic_0_buffer_valid;
  reg        [7:0]    s2_byteLogic_0_buffer_data;
  wire                s2_byteLogic_0_lastUsed;
  wire                s2_byteLogic_0_inputMask;
  wire       [7:0]    s2_byteLogic_0_inputData;
  wire                s2_byteLogic_0_outputMask;
  wire       [7:0]    s2_byteLogic_0_outputData;
  wire                when_DmaSg_l1493;
  reg                 s2_byteLogic_1_buffer_valid;
  reg        [7:0]    s2_byteLogic_1_buffer_data;
  wire                s2_byteLogic_1_lastUsed;
  wire                s2_byteLogic_1_inputMask;
  wire       [7:0]    s2_byteLogic_1_inputData;
  wire                s2_byteLogic_1_outputMask;
  wire       [7:0]    s2_byteLogic_1_outputData;
  wire                when_DmaSg_l1493_1;
  reg                 s2_byteLogic_2_buffer_valid;
  reg        [7:0]    s2_byteLogic_2_buffer_data;
  wire                s2_byteLogic_2_lastUsed;
  wire                s2_byteLogic_2_inputMask;
  wire       [7:0]    s2_byteLogic_2_inputData;
  wire                s2_byteLogic_2_outputMask;
  wire       [7:0]    s2_byteLogic_2_outputData;
  wire                when_DmaSg_l1493_2;
  reg                 s2_byteLogic_3_buffer_valid;
  reg        [7:0]    s2_byteLogic_3_buffer_data;
  wire                s2_byteLogic_3_lastUsed;
  wire                s2_byteLogic_3_inputMask;
  wire       [7:0]    s2_byteLogic_3_inputData;
  wire                s2_byteLogic_3_outputMask;
  wire       [7:0]    s2_byteLogic_3_outputData;
  wire                when_DmaSg_l1493_3;
  reg                 s2_byteLogic_4_buffer_valid;
  reg        [7:0]    s2_byteLogic_4_buffer_data;
  wire                s2_byteLogic_4_lastUsed;
  wire                s2_byteLogic_4_inputMask;
  wire       [7:0]    s2_byteLogic_4_inputData;
  wire                s2_byteLogic_4_outputMask;
  wire       [7:0]    s2_byteLogic_4_outputData;
  wire                when_DmaSg_l1493_4;
  reg                 s2_byteLogic_5_buffer_valid;
  reg        [7:0]    s2_byteLogic_5_buffer_data;
  wire                s2_byteLogic_5_lastUsed;
  wire                s2_byteLogic_5_inputMask;
  wire       [7:0]    s2_byteLogic_5_inputData;
  wire                s2_byteLogic_5_outputMask;
  wire       [7:0]    s2_byteLogic_5_outputData;
  wire                when_DmaSg_l1493_5;
  reg                 s2_byteLogic_6_buffer_valid;
  reg        [7:0]    s2_byteLogic_6_buffer_data;
  wire                s2_byteLogic_6_lastUsed;
  wire                s2_byteLogic_6_inputMask;
  wire       [7:0]    s2_byteLogic_6_inputData;
  wire                s2_byteLogic_6_outputMask;
  wire       [7:0]    s2_byteLogic_6_outputData;
  wire                when_DmaSg_l1493_6;
  reg                 s2_byteLogic_7_buffer_valid;
  reg        [7:0]    s2_byteLogic_7_buffer_data;
  wire                s2_byteLogic_7_lastUsed;
  wire                s2_byteLogic_7_inputMask;
  wire       [7:0]    s2_byteLogic_7_inputData;
  wire                s2_byteLogic_7_outputMask;
  wire       [7:0]    s2_byteLogic_7_outputData;
  wire                when_DmaSg_l1493_7;
  reg                 s2_byteLogic_8_buffer_valid;
  reg        [7:0]    s2_byteLogic_8_buffer_data;
  wire                s2_byteLogic_8_lastUsed;
  wire                s2_byteLogic_8_inputMask;
  wire       [7:0]    s2_byteLogic_8_inputData;
  wire                s2_byteLogic_8_outputMask;
  wire       [7:0]    s2_byteLogic_8_outputData;
  wire                when_DmaSg_l1493_8;
  reg                 s2_byteLogic_9_buffer_valid;
  reg        [7:0]    s2_byteLogic_9_buffer_data;
  wire                s2_byteLogic_9_lastUsed;
  wire                s2_byteLogic_9_inputMask;
  wire       [7:0]    s2_byteLogic_9_inputData;
  wire                s2_byteLogic_9_outputMask;
  wire       [7:0]    s2_byteLogic_9_outputData;
  wire                when_DmaSg_l1493_9;
  reg                 s2_byteLogic_10_buffer_valid;
  reg        [7:0]    s2_byteLogic_10_buffer_data;
  wire                s2_byteLogic_10_lastUsed;
  wire                s2_byteLogic_10_inputMask;
  wire       [7:0]    s2_byteLogic_10_inputData;
  wire                s2_byteLogic_10_outputMask;
  wire       [7:0]    s2_byteLogic_10_outputData;
  wire                when_DmaSg_l1493_10;
  reg                 s2_byteLogic_11_buffer_valid;
  reg        [7:0]    s2_byteLogic_11_buffer_data;
  wire                s2_byteLogic_11_lastUsed;
  wire                s2_byteLogic_11_inputMask;
  wire       [7:0]    s2_byteLogic_11_inputData;
  wire                s2_byteLogic_11_outputMask;
  wire       [7:0]    s2_byteLogic_11_outputData;
  wire                when_DmaSg_l1493_11;
  reg                 s2_byteLogic_12_buffer_valid;
  reg        [7:0]    s2_byteLogic_12_buffer_data;
  wire                s2_byteLogic_12_lastUsed;
  wire                s2_byteLogic_12_inputMask;
  wire       [7:0]    s2_byteLogic_12_inputData;
  wire                s2_byteLogic_12_outputMask;
  wire       [7:0]    s2_byteLogic_12_outputData;
  wire                when_DmaSg_l1493_12;
  reg                 s2_byteLogic_13_buffer_valid;
  reg        [7:0]    s2_byteLogic_13_buffer_data;
  wire                s2_byteLogic_13_lastUsed;
  wire                s2_byteLogic_13_inputMask;
  wire       [7:0]    s2_byteLogic_13_inputData;
  wire                s2_byteLogic_13_outputMask;
  wire       [7:0]    s2_byteLogic_13_outputData;
  wire                when_DmaSg_l1493_13;
  reg                 s2_byteLogic_14_buffer_valid;
  reg        [7:0]    s2_byteLogic_14_buffer_data;
  wire                s2_byteLogic_14_lastUsed;
  wire                s2_byteLogic_14_inputMask;
  wire       [7:0]    s2_byteLogic_14_inputData;
  wire                s2_byteLogic_14_outputMask;
  wire       [7:0]    s2_byteLogic_14_outputData;
  wire                when_DmaSg_l1493_14;
  reg                 s2_byteLogic_15_buffer_valid;
  reg        [7:0]    s2_byteLogic_15_buffer_data;
  wire                s2_byteLogic_15_lastUsed;
  wire                s2_byteLogic_15_inputMask;
  wire       [7:0]    s2_byteLogic_15_inputData;
  wire                s2_byteLogic_15_outputMask;
  wire       [7:0]    s2_byteLogic_15_outputData;
  wire                when_DmaSg_l1493_15;
  reg                 s2_byteLogic_16_buffer_valid;
  reg        [7:0]    s2_byteLogic_16_buffer_data;
  wire                s2_byteLogic_16_lastUsed;
  wire                s2_byteLogic_16_inputMask;
  wire       [7:0]    s2_byteLogic_16_inputData;
  wire                s2_byteLogic_16_outputMask;
  wire       [7:0]    s2_byteLogic_16_outputData;
  wire                when_DmaSg_l1493_16;
  reg                 s2_byteLogic_17_buffer_valid;
  reg        [7:0]    s2_byteLogic_17_buffer_data;
  wire                s2_byteLogic_17_lastUsed;
  wire                s2_byteLogic_17_inputMask;
  wire       [7:0]    s2_byteLogic_17_inputData;
  wire                s2_byteLogic_17_outputMask;
  wire       [7:0]    s2_byteLogic_17_outputData;
  wire                when_DmaSg_l1493_17;
  reg                 s2_byteLogic_18_buffer_valid;
  reg        [7:0]    s2_byteLogic_18_buffer_data;
  wire                s2_byteLogic_18_lastUsed;
  wire                s2_byteLogic_18_inputMask;
  wire       [7:0]    s2_byteLogic_18_inputData;
  wire                s2_byteLogic_18_outputMask;
  wire       [7:0]    s2_byteLogic_18_outputData;
  wire                when_DmaSg_l1493_18;
  reg                 s2_byteLogic_19_buffer_valid;
  reg        [7:0]    s2_byteLogic_19_buffer_data;
  wire                s2_byteLogic_19_lastUsed;
  wire                s2_byteLogic_19_inputMask;
  wire       [7:0]    s2_byteLogic_19_inputData;
  wire                s2_byteLogic_19_outputMask;
  wire       [7:0]    s2_byteLogic_19_outputData;
  wire                when_DmaSg_l1493_19;
  reg                 s2_byteLogic_20_buffer_valid;
  reg        [7:0]    s2_byteLogic_20_buffer_data;
  wire                s2_byteLogic_20_lastUsed;
  wire                s2_byteLogic_20_inputMask;
  wire       [7:0]    s2_byteLogic_20_inputData;
  wire                s2_byteLogic_20_outputMask;
  wire       [7:0]    s2_byteLogic_20_outputData;
  wire                when_DmaSg_l1493_20;
  reg                 s2_byteLogic_21_buffer_valid;
  reg        [7:0]    s2_byteLogic_21_buffer_data;
  wire                s2_byteLogic_21_lastUsed;
  wire                s2_byteLogic_21_inputMask;
  wire       [7:0]    s2_byteLogic_21_inputData;
  wire                s2_byteLogic_21_outputMask;
  wire       [7:0]    s2_byteLogic_21_outputData;
  wire                when_DmaSg_l1493_21;
  reg                 s2_byteLogic_22_buffer_valid;
  reg        [7:0]    s2_byteLogic_22_buffer_data;
  wire                s2_byteLogic_22_lastUsed;
  wire                s2_byteLogic_22_inputMask;
  wire       [7:0]    s2_byteLogic_22_inputData;
  wire                s2_byteLogic_22_outputMask;
  wire       [7:0]    s2_byteLogic_22_outputData;
  wire                when_DmaSg_l1493_22;
  reg                 s2_byteLogic_23_buffer_valid;
  reg        [7:0]    s2_byteLogic_23_buffer_data;
  wire                s2_byteLogic_23_lastUsed;
  wire                s2_byteLogic_23_inputMask;
  wire       [7:0]    s2_byteLogic_23_inputData;
  wire                s2_byteLogic_23_outputMask;
  wire       [7:0]    s2_byteLogic_23_outputData;
  wire                when_DmaSg_l1493_23;
  reg                 s2_byteLogic_24_buffer_valid;
  reg        [7:0]    s2_byteLogic_24_buffer_data;
  wire                s2_byteLogic_24_lastUsed;
  wire                s2_byteLogic_24_inputMask;
  wire       [7:0]    s2_byteLogic_24_inputData;
  wire                s2_byteLogic_24_outputMask;
  wire       [7:0]    s2_byteLogic_24_outputData;
  wire                when_DmaSg_l1493_24;
  reg                 s2_byteLogic_25_buffer_valid;
  reg        [7:0]    s2_byteLogic_25_buffer_data;
  wire                s2_byteLogic_25_lastUsed;
  wire                s2_byteLogic_25_inputMask;
  wire       [7:0]    s2_byteLogic_25_inputData;
  wire                s2_byteLogic_25_outputMask;
  wire       [7:0]    s2_byteLogic_25_outputData;
  wire                when_DmaSg_l1493_25;
  reg                 s2_byteLogic_26_buffer_valid;
  reg        [7:0]    s2_byteLogic_26_buffer_data;
  wire                s2_byteLogic_26_lastUsed;
  wire                s2_byteLogic_26_inputMask;
  wire       [7:0]    s2_byteLogic_26_inputData;
  wire                s2_byteLogic_26_outputMask;
  wire       [7:0]    s2_byteLogic_26_outputData;
  wire                when_DmaSg_l1493_26;
  reg                 s2_byteLogic_27_buffer_valid;
  reg        [7:0]    s2_byteLogic_27_buffer_data;
  wire                s2_byteLogic_27_lastUsed;
  wire                s2_byteLogic_27_inputMask;
  wire       [7:0]    s2_byteLogic_27_inputData;
  wire                s2_byteLogic_27_outputMask;
  wire       [7:0]    s2_byteLogic_27_outputData;
  wire                when_DmaSg_l1493_27;
  reg                 s2_byteLogic_28_buffer_valid;
  reg        [7:0]    s2_byteLogic_28_buffer_data;
  wire                s2_byteLogic_28_lastUsed;
  wire                s2_byteLogic_28_inputMask;
  wire       [7:0]    s2_byteLogic_28_inputData;
  wire                s2_byteLogic_28_outputMask;
  wire       [7:0]    s2_byteLogic_28_outputData;
  wire                when_DmaSg_l1493_28;
  reg                 s2_byteLogic_29_buffer_valid;
  reg        [7:0]    s2_byteLogic_29_buffer_data;
  wire                s2_byteLogic_29_lastUsed;
  wire                s2_byteLogic_29_inputMask;
  wire       [7:0]    s2_byteLogic_29_inputData;
  wire                s2_byteLogic_29_outputMask;
  wire       [7:0]    s2_byteLogic_29_outputData;
  wire                when_DmaSg_l1493_29;
  reg                 s2_byteLogic_30_buffer_valid;
  reg        [7:0]    s2_byteLogic_30_buffer_data;
  wire                s2_byteLogic_30_lastUsed;
  wire                s2_byteLogic_30_inputMask;
  wire       [7:0]    s2_byteLogic_30_inputData;
  wire                s2_byteLogic_30_outputMask;
  wire       [7:0]    s2_byteLogic_30_outputData;
  wire                when_DmaSg_l1493_30;
  reg                 s2_byteLogic_31_buffer_valid;
  reg        [7:0]    s2_byteLogic_31_buffer_data;
  wire                s2_byteLogic_31_lastUsed;
  wire                s2_byteLogic_31_inputMask;
  wire       [7:0]    s2_byteLogic_31_inputData;
  wire                s2_byteLogic_31_outputMask;
  wire       [7:0]    s2_byteLogic_31_outputData;
  wire                when_DmaSg_l1493_31;
  wire                _zz_io_output_usedUntil;
  wire                _zz_io_output_usedUntil_1;
  wire                _zz_io_output_usedUntil_2;
  wire                _zz_io_output_usedUntil_3;
  wire                _zz_io_output_usedUntil_4;

  assign _zz_s0_countOnesLogic_3_13 = _zz_s0_countOnesLogic_3;
  assign _zz_s0_countOnesLogic_3_12 = {2'd0, _zz_s0_countOnesLogic_3_13};
  assign _zz_s0_countOnesLogic_4_13 = {_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3};
  assign _zz_s0_countOnesLogic_4_12 = {1'd0, _zz_s0_countOnesLogic_4_13};
  assign _zz_s0_countOnesLogic_6_9 = (_zz_s0_countOnesLogic_6_10 + _zz_s0_countOnesLogic_6_12);
  assign _zz_s0_countOnesLogic_6_16 = _zz_s0_countOnesLogic_6;
  assign _zz_s0_countOnesLogic_6_15 = {2'd0, _zz_s0_countOnesLogic_6_16};
  assign _zz_s0_countOnesLogic_7_9 = (_zz_s0_countOnesLogic_7_10 + _zz_s0_countOnesLogic_7_12);
  assign _zz_s0_countOnesLogic_7_16 = {_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6};
  assign _zz_s0_countOnesLogic_7_15 = {1'd0, _zz_s0_countOnesLogic_7_16};
  assign _zz_s0_countOnesLogic_8_9 = (_zz_s0_countOnesLogic_8_10 + _zz_s0_countOnesLogic_8_12);
  assign _zz_s0_countOnesLogic_9_9 = (_zz_s0_countOnesLogic_9_10 + _zz_s0_countOnesLogic_9_12);
  assign _zz_s0_countOnesLogic_9_14 = (_zz_s0_countOnesLogic_9_15 + _zz_s0_countOnesLogic_9_17);
  assign _zz_s0_countOnesLogic_9_19 = _zz_s0_countOnesLogic_9;
  assign _zz_s0_countOnesLogic_9_18 = {2'd0, _zz_s0_countOnesLogic_9_19};
  assign _zz_s0_countOnesLogic_10_9 = (_zz_s0_countOnesLogic_10_10 + _zz_s0_countOnesLogic_10_12);
  assign _zz_s0_countOnesLogic_10_14 = (_zz_s0_countOnesLogic_10_15 + _zz_s0_countOnesLogic_10_17);
  assign _zz_s0_countOnesLogic_10_19 = {_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9};
  assign _zz_s0_countOnesLogic_10_18 = {1'd0, _zz_s0_countOnesLogic_10_19};
  assign _zz_s0_countOnesLogic_11_9 = (_zz_s0_countOnesLogic_11_10 + _zz_s0_countOnesLogic_11_12);
  assign _zz_s0_countOnesLogic_11_14 = (_zz_s0_countOnesLogic_11_15 + _zz_s0_countOnesLogic_11_17);
  assign _zz_s0_countOnesLogic_12_9 = (_zz_s0_countOnesLogic_12_10 + _zz_s0_countOnesLogic_12_15);
  assign _zz_s0_countOnesLogic_12_10 = (_zz_s0_countOnesLogic_12_11 + _zz_s0_countOnesLogic_12_13);
  assign _zz_s0_countOnesLogic_12_15 = (_zz_s0_countOnesLogic_12_16 + _zz_s0_countOnesLogic_12_18);
  assign _zz_s0_countOnesLogic_12_22 = _zz_s0_countOnesLogic_12;
  assign _zz_s0_countOnesLogic_12_21 = {2'd0, _zz_s0_countOnesLogic_12_22};
  assign _zz_s0_countOnesLogic_13_9 = (_zz_s0_countOnesLogic_13_10 + _zz_s0_countOnesLogic_13_15);
  assign _zz_s0_countOnesLogic_13_10 = (_zz_s0_countOnesLogic_13_11 + _zz_s0_countOnesLogic_13_13);
  assign _zz_s0_countOnesLogic_13_15 = (_zz_s0_countOnesLogic_13_16 + _zz_s0_countOnesLogic_13_18);
  assign _zz_s0_countOnesLogic_13_22 = {_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12};
  assign _zz_s0_countOnesLogic_13_21 = {1'd0, _zz_s0_countOnesLogic_13_22};
  assign _zz_s0_countOnesLogic_14_9 = (_zz_s0_countOnesLogic_14_10 + _zz_s0_countOnesLogic_14_15);
  assign _zz_s0_countOnesLogic_14_10 = (_zz_s0_countOnesLogic_14_11 + _zz_s0_countOnesLogic_14_13);
  assign _zz_s0_countOnesLogic_14_15 = (_zz_s0_countOnesLogic_14_16 + _zz_s0_countOnesLogic_14_18);
  assign _zz_s0_countOnesLogic_15_9 = (_zz_s0_countOnesLogic_15_10 + _zz_s0_countOnesLogic_15_15);
  assign _zz_s0_countOnesLogic_15_10 = (_zz_s0_countOnesLogic_15_11 + _zz_s0_countOnesLogic_15_13);
  assign _zz_s0_countOnesLogic_15_15 = (_zz_s0_countOnesLogic_15_16 + _zz_s0_countOnesLogic_15_18);
  assign _zz_s0_countOnesLogic_15_20 = (_zz_s0_countOnesLogic_15_21 + _zz_s0_countOnesLogic_15_23);
  assign _zz_s0_countOnesLogic_15_25 = _zz_s0_countOnesLogic_15;
  assign _zz_s0_countOnesLogic_15_24 = {2'd0, _zz_s0_countOnesLogic_15_25};
  assign _zz_s0_countOnesLogic_16_9 = (_zz_s0_countOnesLogic_16_10 + _zz_s0_countOnesLogic_16_15);
  assign _zz_s0_countOnesLogic_16_10 = (_zz_s0_countOnesLogic_16_11 + _zz_s0_countOnesLogic_16_13);
  assign _zz_s0_countOnesLogic_16_15 = (_zz_s0_countOnesLogic_16_16 + _zz_s0_countOnesLogic_16_18);
  assign _zz_s0_countOnesLogic_16_20 = (_zz_s0_countOnesLogic_16_21 + _zz_s0_countOnesLogic_16_23);
  assign _zz_s0_countOnesLogic_16_25 = {_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15};
  assign _zz_s0_countOnesLogic_16_24 = {1'd0, _zz_s0_countOnesLogic_16_25};
  assign _zz_s0_countOnesLogic_17_9 = (_zz_s0_countOnesLogic_17_10 + _zz_s0_countOnesLogic_17_15);
  assign _zz_s0_countOnesLogic_17_10 = (_zz_s0_countOnesLogic_17_11 + _zz_s0_countOnesLogic_17_13);
  assign _zz_s0_countOnesLogic_17_15 = (_zz_s0_countOnesLogic_17_16 + _zz_s0_countOnesLogic_17_18);
  assign _zz_s0_countOnesLogic_17_20 = (_zz_s0_countOnesLogic_17_21 + _zz_s0_countOnesLogic_17_23);
  assign _zz_s0_countOnesLogic_18_9 = (_zz_s0_countOnesLogic_18_10 + _zz_s0_countOnesLogic_18_15);
  assign _zz_s0_countOnesLogic_18_10 = (_zz_s0_countOnesLogic_18_11 + _zz_s0_countOnesLogic_18_13);
  assign _zz_s0_countOnesLogic_18_15 = (_zz_s0_countOnesLogic_18_16 + _zz_s0_countOnesLogic_18_18);
  assign _zz_s0_countOnesLogic_18_20 = (_zz_s0_countOnesLogic_18_21 + _zz_s0_countOnesLogic_18_26);
  assign _zz_s0_countOnesLogic_18_21 = (_zz_s0_countOnesLogic_18_22 + _zz_s0_countOnesLogic_18_24);
  assign _zz_s0_countOnesLogic_18_28 = _zz_s0_countOnesLogic_18;
  assign _zz_s0_countOnesLogic_18_27 = {2'd0, _zz_s0_countOnesLogic_18_28};
  assign _zz_s0_countOnesLogic_19_9 = (_zz_s0_countOnesLogic_19_10 + _zz_s0_countOnesLogic_19_15);
  assign _zz_s0_countOnesLogic_19_10 = (_zz_s0_countOnesLogic_19_11 + _zz_s0_countOnesLogic_19_13);
  assign _zz_s0_countOnesLogic_19_15 = (_zz_s0_countOnesLogic_19_16 + _zz_s0_countOnesLogic_19_18);
  assign _zz_s0_countOnesLogic_19_20 = (_zz_s0_countOnesLogic_19_21 + _zz_s0_countOnesLogic_19_26);
  assign _zz_s0_countOnesLogic_19_21 = (_zz_s0_countOnesLogic_19_22 + _zz_s0_countOnesLogic_19_24);
  assign _zz_s0_countOnesLogic_19_28 = {_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18};
  assign _zz_s0_countOnesLogic_19_27 = {1'd0, _zz_s0_countOnesLogic_19_28};
  assign _zz_s0_countOnesLogic_20_9 = (_zz_s0_countOnesLogic_20_10 + _zz_s0_countOnesLogic_20_15);
  assign _zz_s0_countOnesLogic_20_10 = (_zz_s0_countOnesLogic_20_11 + _zz_s0_countOnesLogic_20_13);
  assign _zz_s0_countOnesLogic_20_15 = (_zz_s0_countOnesLogic_20_16 + _zz_s0_countOnesLogic_20_18);
  assign _zz_s0_countOnesLogic_20_20 = (_zz_s0_countOnesLogic_20_21 + _zz_s0_countOnesLogic_20_26);
  assign _zz_s0_countOnesLogic_20_21 = (_zz_s0_countOnesLogic_20_22 + _zz_s0_countOnesLogic_20_24);
  assign _zz_s0_countOnesLogic_21_9 = (_zz_s0_countOnesLogic_21_10 + _zz_s0_countOnesLogic_21_15);
  assign _zz_s0_countOnesLogic_21_10 = (_zz_s0_countOnesLogic_21_11 + _zz_s0_countOnesLogic_21_13);
  assign _zz_s0_countOnesLogic_21_15 = (_zz_s0_countOnesLogic_21_16 + _zz_s0_countOnesLogic_21_18);
  assign _zz_s0_countOnesLogic_21_20 = (_zz_s0_countOnesLogic_21_21 + _zz_s0_countOnesLogic_21_26);
  assign _zz_s0_countOnesLogic_21_21 = (_zz_s0_countOnesLogic_21_22 + _zz_s0_countOnesLogic_21_24);
  assign _zz_s0_countOnesLogic_21_26 = (_zz_s0_countOnesLogic_21_27 + _zz_s0_countOnesLogic_21_29);
  assign _zz_s0_countOnesLogic_21_31 = _zz_s0_countOnesLogic_21;
  assign _zz_s0_countOnesLogic_21_30 = {2'd0, _zz_s0_countOnesLogic_21_31};
  assign _zz_s0_countOnesLogic_22_9 = (_zz_s0_countOnesLogic_22_10 + _zz_s0_countOnesLogic_22_15);
  assign _zz_s0_countOnesLogic_22_10 = (_zz_s0_countOnesLogic_22_11 + _zz_s0_countOnesLogic_22_13);
  assign _zz_s0_countOnesLogic_22_15 = (_zz_s0_countOnesLogic_22_16 + _zz_s0_countOnesLogic_22_18);
  assign _zz_s0_countOnesLogic_22_20 = (_zz_s0_countOnesLogic_22_21 + _zz_s0_countOnesLogic_22_26);
  assign _zz_s0_countOnesLogic_22_21 = (_zz_s0_countOnesLogic_22_22 + _zz_s0_countOnesLogic_22_24);
  assign _zz_s0_countOnesLogic_22_26 = (_zz_s0_countOnesLogic_22_27 + _zz_s0_countOnesLogic_22_29);
  assign _zz_s0_countOnesLogic_22_31 = {_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21};
  assign _zz_s0_countOnesLogic_22_30 = {1'd0, _zz_s0_countOnesLogic_22_31};
  assign _zz_s0_countOnesLogic_23_9 = (_zz_s0_countOnesLogic_23_10 + _zz_s0_countOnesLogic_23_15);
  assign _zz_s0_countOnesLogic_23_10 = (_zz_s0_countOnesLogic_23_11 + _zz_s0_countOnesLogic_23_13);
  assign _zz_s0_countOnesLogic_23_15 = (_zz_s0_countOnesLogic_23_16 + _zz_s0_countOnesLogic_23_18);
  assign _zz_s0_countOnesLogic_23_20 = (_zz_s0_countOnesLogic_23_21 + _zz_s0_countOnesLogic_23_26);
  assign _zz_s0_countOnesLogic_23_21 = (_zz_s0_countOnesLogic_23_22 + _zz_s0_countOnesLogic_23_24);
  assign _zz_s0_countOnesLogic_23_26 = (_zz_s0_countOnesLogic_23_27 + _zz_s0_countOnesLogic_23_29);
  assign _zz_s0_countOnesLogic_24_9 = (_zz_s0_countOnesLogic_24_10 + _zz_s0_countOnesLogic_24_21);
  assign _zz_s0_countOnesLogic_24_10 = (_zz_s0_countOnesLogic_24_11 + _zz_s0_countOnesLogic_24_16);
  assign _zz_s0_countOnesLogic_24_11 = (_zz_s0_countOnesLogic_24_12 + _zz_s0_countOnesLogic_24_14);
  assign _zz_s0_countOnesLogic_24_16 = (_zz_s0_countOnesLogic_24_17 + _zz_s0_countOnesLogic_24_19);
  assign _zz_s0_countOnesLogic_24_21 = (_zz_s0_countOnesLogic_24_22 + _zz_s0_countOnesLogic_24_27);
  assign _zz_s0_countOnesLogic_24_22 = (_zz_s0_countOnesLogic_24_23 + _zz_s0_countOnesLogic_24_25);
  assign _zz_s0_countOnesLogic_24_27 = (_zz_s0_countOnesLogic_24_28 + _zz_s0_countOnesLogic_24_30);
  assign _zz_s0_countOnesLogic_24_34 = _zz_s0_countOnesLogic_24;
  assign _zz_s0_countOnesLogic_24_33 = {2'd0, _zz_s0_countOnesLogic_24_34};
  assign _zz_s0_countOnesLogic_25_9 = (_zz_s0_countOnesLogic_25_10 + _zz_s0_countOnesLogic_25_21);
  assign _zz_s0_countOnesLogic_25_10 = (_zz_s0_countOnesLogic_25_11 + _zz_s0_countOnesLogic_25_16);
  assign _zz_s0_countOnesLogic_25_11 = (_zz_s0_countOnesLogic_25_12 + _zz_s0_countOnesLogic_25_14);
  assign _zz_s0_countOnesLogic_25_16 = (_zz_s0_countOnesLogic_25_17 + _zz_s0_countOnesLogic_25_19);
  assign _zz_s0_countOnesLogic_25_21 = (_zz_s0_countOnesLogic_25_22 + _zz_s0_countOnesLogic_25_27);
  assign _zz_s0_countOnesLogic_25_22 = (_zz_s0_countOnesLogic_25_23 + _zz_s0_countOnesLogic_25_25);
  assign _zz_s0_countOnesLogic_25_27 = (_zz_s0_countOnesLogic_25_28 + _zz_s0_countOnesLogic_25_30);
  assign _zz_s0_countOnesLogic_25_34 = {_zz_s0_countOnesLogic_25,_zz_s0_countOnesLogic_24};
  assign _zz_s0_countOnesLogic_25_33 = {1'd0, _zz_s0_countOnesLogic_25_34};
  assign _zz_s0_countOnesLogic_26_9 = (_zz_s0_countOnesLogic_26_10 + _zz_s0_countOnesLogic_26_21);
  assign _zz_s0_countOnesLogic_26_10 = (_zz_s0_countOnesLogic_26_11 + _zz_s0_countOnesLogic_26_16);
  assign _zz_s0_countOnesLogic_26_11 = (_zz_s0_countOnesLogic_26_12 + _zz_s0_countOnesLogic_26_14);
  assign _zz_s0_countOnesLogic_26_16 = (_zz_s0_countOnesLogic_26_17 + _zz_s0_countOnesLogic_26_19);
  assign _zz_s0_countOnesLogic_26_21 = (_zz_s0_countOnesLogic_26_22 + _zz_s0_countOnesLogic_26_27);
  assign _zz_s0_countOnesLogic_26_22 = (_zz_s0_countOnesLogic_26_23 + _zz_s0_countOnesLogic_26_25);
  assign _zz_s0_countOnesLogic_26_27 = (_zz_s0_countOnesLogic_26_28 + _zz_s0_countOnesLogic_26_30);
  assign _zz_s0_countOnesLogic_27_9 = (_zz_s0_countOnesLogic_27_10 + _zz_s0_countOnesLogic_27_21);
  assign _zz_s0_countOnesLogic_27_10 = (_zz_s0_countOnesLogic_27_11 + _zz_s0_countOnesLogic_27_16);
  assign _zz_s0_countOnesLogic_27_11 = (_zz_s0_countOnesLogic_27_12 + _zz_s0_countOnesLogic_27_14);
  assign _zz_s0_countOnesLogic_27_16 = (_zz_s0_countOnesLogic_27_17 + _zz_s0_countOnesLogic_27_19);
  assign _zz_s0_countOnesLogic_27_21 = (_zz_s0_countOnesLogic_27_22 + _zz_s0_countOnesLogic_27_27);
  assign _zz_s0_countOnesLogic_27_22 = (_zz_s0_countOnesLogic_27_23 + _zz_s0_countOnesLogic_27_25);
  assign _zz_s0_countOnesLogic_27_27 = (_zz_s0_countOnesLogic_27_28 + _zz_s0_countOnesLogic_27_30);
  assign _zz_s0_countOnesLogic_27_32 = (_zz_s0_countOnesLogic_27_33 + _zz_s0_countOnesLogic_27_35);
  assign _zz_s0_countOnesLogic_27_37 = _zz_s0_countOnesLogic_27;
  assign _zz_s0_countOnesLogic_27_36 = {2'd0, _zz_s0_countOnesLogic_27_37};
  assign _zz_s0_countOnesLogic_28_9 = (_zz_s0_countOnesLogic_28_10 + _zz_s0_countOnesLogic_28_21);
  assign _zz_s0_countOnesLogic_28_10 = (_zz_s0_countOnesLogic_28_11 + _zz_s0_countOnesLogic_28_16);
  assign _zz_s0_countOnesLogic_28_11 = (_zz_s0_countOnesLogic_28_12 + _zz_s0_countOnesLogic_28_14);
  assign _zz_s0_countOnesLogic_28_16 = (_zz_s0_countOnesLogic_28_17 + _zz_s0_countOnesLogic_28_19);
  assign _zz_s0_countOnesLogic_28_21 = (_zz_s0_countOnesLogic_28_22 + _zz_s0_countOnesLogic_28_27);
  assign _zz_s0_countOnesLogic_28_22 = (_zz_s0_countOnesLogic_28_23 + _zz_s0_countOnesLogic_28_25);
  assign _zz_s0_countOnesLogic_28_27 = (_zz_s0_countOnesLogic_28_28 + _zz_s0_countOnesLogic_28_30);
  assign _zz_s0_countOnesLogic_28_32 = (_zz_s0_countOnesLogic_28_33 + _zz_s0_countOnesLogic_28_35);
  assign _zz_s0_countOnesLogic_28_37 = {_zz_s0_countOnesLogic_28,_zz_s0_countOnesLogic_27};
  assign _zz_s0_countOnesLogic_28_36 = {1'd0, _zz_s0_countOnesLogic_28_37};
  assign _zz_s0_countOnesLogic_29_9 = (_zz_s0_countOnesLogic_29_10 + _zz_s0_countOnesLogic_29_21);
  assign _zz_s0_countOnesLogic_29_10 = (_zz_s0_countOnesLogic_29_11 + _zz_s0_countOnesLogic_29_16);
  assign _zz_s0_countOnesLogic_29_11 = (_zz_s0_countOnesLogic_29_12 + _zz_s0_countOnesLogic_29_14);
  assign _zz_s0_countOnesLogic_29_16 = (_zz_s0_countOnesLogic_29_17 + _zz_s0_countOnesLogic_29_19);
  assign _zz_s0_countOnesLogic_29_21 = (_zz_s0_countOnesLogic_29_22 + _zz_s0_countOnesLogic_29_27);
  assign _zz_s0_countOnesLogic_29_22 = (_zz_s0_countOnesLogic_29_23 + _zz_s0_countOnesLogic_29_25);
  assign _zz_s0_countOnesLogic_29_27 = (_zz_s0_countOnesLogic_29_28 + _zz_s0_countOnesLogic_29_30);
  assign _zz_s0_countOnesLogic_29_32 = (_zz_s0_countOnesLogic_29_33 + _zz_s0_countOnesLogic_29_35);
  assign _zz_s0_countOnesLogic_30_9 = (_zz_s0_countOnesLogic_30_10 + _zz_s0_countOnesLogic_30_21);
  assign _zz_s0_countOnesLogic_30_10 = (_zz_s0_countOnesLogic_30_11 + _zz_s0_countOnesLogic_30_16);
  assign _zz_s0_countOnesLogic_30_11 = (_zz_s0_countOnesLogic_30_12 + _zz_s0_countOnesLogic_30_14);
  assign _zz_s0_countOnesLogic_30_16 = (_zz_s0_countOnesLogic_30_17 + _zz_s0_countOnesLogic_30_19);
  assign _zz_s0_countOnesLogic_30_21 = (_zz_s0_countOnesLogic_30_22 + _zz_s0_countOnesLogic_30_27);
  assign _zz_s0_countOnesLogic_30_22 = (_zz_s0_countOnesLogic_30_23 + _zz_s0_countOnesLogic_30_25);
  assign _zz_s0_countOnesLogic_30_27 = (_zz_s0_countOnesLogic_30_28 + _zz_s0_countOnesLogic_30_30);
  assign _zz_s0_countOnesLogic_30_32 = (_zz_s0_countOnesLogic_30_33 + _zz_s0_countOnesLogic_30_38);
  assign _zz_s0_countOnesLogic_30_33 = (_zz_s0_countOnesLogic_30_34 + _zz_s0_countOnesLogic_30_36);
  assign _zz_s0_countOnesLogic_30_40 = _zz_s0_countOnesLogic_30;
  assign _zz_s0_countOnesLogic_30_39 = {2'd0, _zz_s0_countOnesLogic_30_40};
  assign _zz_s0_countOnesLogic_31_8 = (_zz_s0_countOnesLogic_31_9 + _zz_s0_countOnesLogic_31_20);
  assign _zz_s0_countOnesLogic_31_9 = (_zz_s0_countOnesLogic_31_10 + _zz_s0_countOnesLogic_31_15);
  assign _zz_s0_countOnesLogic_31_10 = (_zz_s0_countOnesLogic_31_11 + _zz_s0_countOnesLogic_31_13);
  assign _zz_s0_countOnesLogic_31_15 = (_zz_s0_countOnesLogic_31_16 + _zz_s0_countOnesLogic_31_18);
  assign _zz_s0_countOnesLogic_31_20 = (_zz_s0_countOnesLogic_31_21 + _zz_s0_countOnesLogic_31_26);
  assign _zz_s0_countOnesLogic_31_21 = (_zz_s0_countOnesLogic_31_22 + _zz_s0_countOnesLogic_31_24);
  assign _zz_s0_countOnesLogic_31_26 = (_zz_s0_countOnesLogic_31_27 + _zz_s0_countOnesLogic_31_29);
  assign _zz_s0_countOnesLogic_31_31 = (_zz_s0_countOnesLogic_31_32 + _zz_s0_countOnesLogic_31_37);
  assign _zz_s0_countOnesLogic_31_32 = (_zz_s0_countOnesLogic_31_33 + _zz_s0_countOnesLogic_31_35);
  assign _zz_s0_countOnesLogic_31_39 = {s0_input_payload_mask[31],_zz_s0_countOnesLogic_30};
  assign _zz_s0_countOnesLogic_31_38 = {1'd0, _zz_s0_countOnesLogic_31_39};
  assign _zz_s1_offsetNext = {1'd0, s1_offset};
  assign _zz_s1_byteCounter = {8'd0, s1_input_payload_countOnes_31};
  assign _zz_s1_inputIndexes_1 = {4'd0, s1_input_payload_countOnes_0};
  assign _zz_s1_inputIndexes_2 = {3'd0, s1_input_payload_countOnes_1};
  assign _zz_s1_inputIndexes_3 = {3'd0, s1_input_payload_countOnes_2};
  assign _zz_s1_inputIndexes_4 = {2'd0, s1_input_payload_countOnes_3};
  assign _zz_s1_inputIndexes_5 = {2'd0, s1_input_payload_countOnes_4};
  assign _zz_s1_inputIndexes_6 = {2'd0, s1_input_payload_countOnes_5};
  assign _zz_s1_inputIndexes_7 = {2'd0, s1_input_payload_countOnes_6};
  assign _zz_s1_inputIndexes_8 = {1'd0, s1_input_payload_countOnes_7};
  assign _zz_s1_inputIndexes_9 = {1'd0, s1_input_payload_countOnes_8};
  assign _zz_s1_inputIndexes_10 = {1'd0, s1_input_payload_countOnes_9};
  assign _zz_s1_inputIndexes_11 = {1'd0, s1_input_payload_countOnes_10};
  assign _zz_s1_inputIndexes_12 = {1'd0, s1_input_payload_countOnes_11};
  assign _zz_s1_inputIndexes_13 = {1'd0, s1_input_payload_countOnes_12};
  assign _zz_s1_inputIndexes_14 = {1'd0, s1_input_payload_countOnes_13};
  assign _zz_s1_inputIndexes_15 = {1'd0, s1_input_payload_countOnes_14};
  assign _zz_when_DmaSg_l1464 = {1'd0, io_burstLength};
  assign _zz_s0_countOnesLogic_0_2 = _zz_s0_countOnesLogic_0;
  assign _zz_s0_countOnesLogic_1_2 = {_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0};
  assign _zz_s0_countOnesLogic_2_2 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_3_10 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_4_10 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_5_10 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_5_12 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_6_11 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_6_13 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_7_11 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_7_13 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_8_11 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_8_13 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_8_15 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_9_11 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_9_13 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_9_16 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_10_11 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_10_13 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_10_16 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_11_11 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_11_13 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_11_16 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_11_18 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_12_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_12_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_12_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_12_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_13_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_13_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_13_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_13_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_14_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_14_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_14_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_14_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_14_21 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_15_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_15_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_15_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_15_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_15_22 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_16_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_16_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_16_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_16_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_16_22 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_17_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_17_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_17_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_17_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_17_22 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_17_24 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_18_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_18_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_18_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_18_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_18_23 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_18_25 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_19_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_19_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_19_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_19_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_19_23 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_19_25 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_20_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_20_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_20_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_20_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_20_23 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_20_25 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_20_27 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_21_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_21_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_21_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_21_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_21_23 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_21_25 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_21_28 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_22_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_22_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_22_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_22_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_22_23 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_22_25 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_22_28 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_23_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_23_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_23_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_23_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_23_23 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_23_25 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_23_28 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_23_30 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_24_13 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_24_15 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_24_18 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_24_20 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_24_24 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_24_26 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_24_29 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_24_31 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_25_13 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_25_15 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_25_18 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_25_20 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_25_24 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_25_26 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_25_29 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_25_31 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_26_13 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_26_15 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_26_18 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_26_20 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_26_24 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_26_26 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_26_29 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_26_31 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_26_33 = {_zz_s0_countOnesLogic_26,{_zz_s0_countOnesLogic_25,_zz_s0_countOnesLogic_24}};
  assign _zz_s0_countOnesLogic_27_13 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_27_15 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_27_18 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_27_20 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_27_24 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_27_26 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_27_29 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_27_31 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_27_34 = {_zz_s0_countOnesLogic_26,{_zz_s0_countOnesLogic_25,_zz_s0_countOnesLogic_24}};
  assign _zz_s0_countOnesLogic_28_13 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_28_15 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_28_18 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_28_20 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_28_24 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_28_26 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_28_29 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_28_31 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_28_34 = {_zz_s0_countOnesLogic_26,{_zz_s0_countOnesLogic_25,_zz_s0_countOnesLogic_24}};
  assign _zz_s0_countOnesLogic_29_13 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_29_15 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_29_18 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_29_20 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_29_24 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_29_26 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_29_29 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_29_31 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_29_34 = {_zz_s0_countOnesLogic_26,{_zz_s0_countOnesLogic_25,_zz_s0_countOnesLogic_24}};
  assign _zz_s0_countOnesLogic_29_36 = {_zz_s0_countOnesLogic_29,{_zz_s0_countOnesLogic_28,_zz_s0_countOnesLogic_27}};
  assign _zz_s0_countOnesLogic_30_13 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_30_15 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_30_18 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_30_20 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_30_24 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_30_26 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_30_29 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_30_31 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_30_35 = {_zz_s0_countOnesLogic_26,{_zz_s0_countOnesLogic_25,_zz_s0_countOnesLogic_24}};
  assign _zz_s0_countOnesLogic_30_37 = {_zz_s0_countOnesLogic_29,{_zz_s0_countOnesLogic_28,_zz_s0_countOnesLogic_27}};
  assign _zz_s0_countOnesLogic_31_12 = {_zz_s0_countOnesLogic_2,{_zz_s0_countOnesLogic_1,_zz_s0_countOnesLogic_0}};
  assign _zz_s0_countOnesLogic_31_14 = {_zz_s0_countOnesLogic_5,{_zz_s0_countOnesLogic_4,_zz_s0_countOnesLogic_3}};
  assign _zz_s0_countOnesLogic_31_17 = {_zz_s0_countOnesLogic_8,{_zz_s0_countOnesLogic_7,_zz_s0_countOnesLogic_6}};
  assign _zz_s0_countOnesLogic_31_19 = {_zz_s0_countOnesLogic_11,{_zz_s0_countOnesLogic_10,_zz_s0_countOnesLogic_9}};
  assign _zz_s0_countOnesLogic_31_23 = {_zz_s0_countOnesLogic_14,{_zz_s0_countOnesLogic_13,_zz_s0_countOnesLogic_12}};
  assign _zz_s0_countOnesLogic_31_25 = {_zz_s0_countOnesLogic_17,{_zz_s0_countOnesLogic_16,_zz_s0_countOnesLogic_15}};
  assign _zz_s0_countOnesLogic_31_28 = {_zz_s0_countOnesLogic_20,{_zz_s0_countOnesLogic_19,_zz_s0_countOnesLogic_18}};
  assign _zz_s0_countOnesLogic_31_30 = {_zz_s0_countOnesLogic_23,{_zz_s0_countOnesLogic_22,_zz_s0_countOnesLogic_21}};
  assign _zz_s0_countOnesLogic_31_34 = {_zz_s0_countOnesLogic_26,{_zz_s0_countOnesLogic_25,_zz_s0_countOnesLogic_24}};
  assign _zz_s0_countOnesLogic_31_36 = {_zz_s0_countOnesLogic_29,{_zz_s0_countOnesLogic_28,_zz_s0_countOnesLogic_27}};
  assign _zz_io_output_usedUntil_6 = {_zz_io_output_usedUntil_4,{_zz_io_output_usedUntil_3,{_zz_io_output_usedUntil_2,{_zz_io_output_usedUntil_1,_zz_io_output_usedUntil}}}};
  assign _zz_s1_outputPayload_selValid_992 = _zz_s1_outputPayload_selValid_22;
  assign _zz_s1_outputPayload_selValid_993 = {_zz_s1_outputPayload_selValid_21,{_zz_s1_outputPayload_selValid_20,{_zz_s1_outputPayload_selValid_19,{_zz_s1_outputPayload_selValid_18,{_zz_s1_outputPayload_selValid_17,{_zz_s1_outputPayload_selValid_16,{_zz_s1_outputPayload_selValid_15,{_zz_s1_outputPayload_selValid_14,{_zz_s1_outputPayload_selValid_13,{_zz_s1_outputPayload_selValid_12,{_zz_s1_outputPayload_selValid_994,_zz_s1_outputPayload_selValid_995}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_994 = _zz_s1_outputPayload_selValid_11;
  assign _zz_s1_outputPayload_selValid_995 = {_zz_s1_outputPayload_selValid_10,{_zz_s1_outputPayload_selValid_9,{_zz_s1_outputPayload_selValid_8,{_zz_s1_outputPayload_selValid_7,{_zz_s1_outputPayload_selValid_6,{_zz_s1_outputPayload_selValid_5,{_zz_s1_outputPayload_selValid_4,{_zz_s1_outputPayload_selValid_3,{_zz_s1_outputPayload_selValid_2,{_zz_s1_outputPayload_selValid_1,{_zz_s1_outputPayload_selValid_996,_zz_s1_outputPayload_selValid_997}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_996 = _zz_s1_outputPayload_selValid;
  assign _zz_s1_outputPayload_selValid_997 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h0));
  assign _zz_s1_outputPayload_selValid_998 = _zz_s1_outputPayload_selValid_53;
  assign _zz_s1_outputPayload_selValid_999 = {_zz_s1_outputPayload_selValid_52,{_zz_s1_outputPayload_selValid_51,{_zz_s1_outputPayload_selValid_50,{_zz_s1_outputPayload_selValid_49,{_zz_s1_outputPayload_selValid_48,{_zz_s1_outputPayload_selValid_47,{_zz_s1_outputPayload_selValid_46,{_zz_s1_outputPayload_selValid_45,{_zz_s1_outputPayload_selValid_44,{_zz_s1_outputPayload_selValid_43,{_zz_s1_outputPayload_selValid_1000,_zz_s1_outputPayload_selValid_1001}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1000 = _zz_s1_outputPayload_selValid_42;
  assign _zz_s1_outputPayload_selValid_1001 = {_zz_s1_outputPayload_selValid_41,{_zz_s1_outputPayload_selValid_40,{_zz_s1_outputPayload_selValid_39,{_zz_s1_outputPayload_selValid_38,{_zz_s1_outputPayload_selValid_37,{_zz_s1_outputPayload_selValid_36,{_zz_s1_outputPayload_selValid_35,{_zz_s1_outputPayload_selValid_34,{_zz_s1_outputPayload_selValid_33,{_zz_s1_outputPayload_selValid_32,{_zz_s1_outputPayload_selValid_1002,_zz_s1_outputPayload_selValid_1003}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1002 = _zz_s1_outputPayload_selValid_31;
  assign _zz_s1_outputPayload_selValid_1003 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h01));
  assign _zz_s1_outputPayload_selValid_1004 = _zz_s1_outputPayload_selValid_84;
  assign _zz_s1_outputPayload_selValid_1005 = {_zz_s1_outputPayload_selValid_83,{_zz_s1_outputPayload_selValid_82,{_zz_s1_outputPayload_selValid_81,{_zz_s1_outputPayload_selValid_80,{_zz_s1_outputPayload_selValid_79,{_zz_s1_outputPayload_selValid_78,{_zz_s1_outputPayload_selValid_77,{_zz_s1_outputPayload_selValid_76,{_zz_s1_outputPayload_selValid_75,{_zz_s1_outputPayload_selValid_74,{_zz_s1_outputPayload_selValid_1006,_zz_s1_outputPayload_selValid_1007}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1006 = _zz_s1_outputPayload_selValid_73;
  assign _zz_s1_outputPayload_selValid_1007 = {_zz_s1_outputPayload_selValid_72,{_zz_s1_outputPayload_selValid_71,{_zz_s1_outputPayload_selValid_70,{_zz_s1_outputPayload_selValid_69,{_zz_s1_outputPayload_selValid_68,{_zz_s1_outputPayload_selValid_67,{_zz_s1_outputPayload_selValid_66,{_zz_s1_outputPayload_selValid_65,{_zz_s1_outputPayload_selValid_64,{_zz_s1_outputPayload_selValid_63,{_zz_s1_outputPayload_selValid_1008,_zz_s1_outputPayload_selValid_1009}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1008 = _zz_s1_outputPayload_selValid_62;
  assign _zz_s1_outputPayload_selValid_1009 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h02));
  assign _zz_s1_outputPayload_selValid_1010 = _zz_s1_outputPayload_selValid_115;
  assign _zz_s1_outputPayload_selValid_1011 = {_zz_s1_outputPayload_selValid_114,{_zz_s1_outputPayload_selValid_113,{_zz_s1_outputPayload_selValid_112,{_zz_s1_outputPayload_selValid_111,{_zz_s1_outputPayload_selValid_110,{_zz_s1_outputPayload_selValid_109,{_zz_s1_outputPayload_selValid_108,{_zz_s1_outputPayload_selValid_107,{_zz_s1_outputPayload_selValid_106,{_zz_s1_outputPayload_selValid_105,{_zz_s1_outputPayload_selValid_1012,_zz_s1_outputPayload_selValid_1013}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1012 = _zz_s1_outputPayload_selValid_104;
  assign _zz_s1_outputPayload_selValid_1013 = {_zz_s1_outputPayload_selValid_103,{_zz_s1_outputPayload_selValid_102,{_zz_s1_outputPayload_selValid_101,{_zz_s1_outputPayload_selValid_100,{_zz_s1_outputPayload_selValid_99,{_zz_s1_outputPayload_selValid_98,{_zz_s1_outputPayload_selValid_97,{_zz_s1_outputPayload_selValid_96,{_zz_s1_outputPayload_selValid_95,{_zz_s1_outputPayload_selValid_94,{_zz_s1_outputPayload_selValid_1014,_zz_s1_outputPayload_selValid_1015}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1014 = _zz_s1_outputPayload_selValid_93;
  assign _zz_s1_outputPayload_selValid_1015 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h03));
  assign _zz_s1_outputPayload_selValid_1016 = _zz_s1_outputPayload_selValid_146;
  assign _zz_s1_outputPayload_selValid_1017 = {_zz_s1_outputPayload_selValid_145,{_zz_s1_outputPayload_selValid_144,{_zz_s1_outputPayload_selValid_143,{_zz_s1_outputPayload_selValid_142,{_zz_s1_outputPayload_selValid_141,{_zz_s1_outputPayload_selValid_140,{_zz_s1_outputPayload_selValid_139,{_zz_s1_outputPayload_selValid_138,{_zz_s1_outputPayload_selValid_137,{_zz_s1_outputPayload_selValid_136,{_zz_s1_outputPayload_selValid_1018,_zz_s1_outputPayload_selValid_1019}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1018 = _zz_s1_outputPayload_selValid_135;
  assign _zz_s1_outputPayload_selValid_1019 = {_zz_s1_outputPayload_selValid_134,{_zz_s1_outputPayload_selValid_133,{_zz_s1_outputPayload_selValid_132,{_zz_s1_outputPayload_selValid_131,{_zz_s1_outputPayload_selValid_130,{_zz_s1_outputPayload_selValid_129,{_zz_s1_outputPayload_selValid_128,{_zz_s1_outputPayload_selValid_127,{_zz_s1_outputPayload_selValid_126,{_zz_s1_outputPayload_selValid_125,{_zz_s1_outputPayload_selValid_1020,_zz_s1_outputPayload_selValid_1021}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1020 = _zz_s1_outputPayload_selValid_124;
  assign _zz_s1_outputPayload_selValid_1021 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h04));
  assign _zz_s1_outputPayload_selValid_1022 = _zz_s1_outputPayload_selValid_177;
  assign _zz_s1_outputPayload_selValid_1023 = {_zz_s1_outputPayload_selValid_176,{_zz_s1_outputPayload_selValid_175,{_zz_s1_outputPayload_selValid_174,{_zz_s1_outputPayload_selValid_173,{_zz_s1_outputPayload_selValid_172,{_zz_s1_outputPayload_selValid_171,{_zz_s1_outputPayload_selValid_170,{_zz_s1_outputPayload_selValid_169,{_zz_s1_outputPayload_selValid_168,{_zz_s1_outputPayload_selValid_167,{_zz_s1_outputPayload_selValid_1024,_zz_s1_outputPayload_selValid_1025}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1024 = _zz_s1_outputPayload_selValid_166;
  assign _zz_s1_outputPayload_selValid_1025 = {_zz_s1_outputPayload_selValid_165,{_zz_s1_outputPayload_selValid_164,{_zz_s1_outputPayload_selValid_163,{_zz_s1_outputPayload_selValid_162,{_zz_s1_outputPayload_selValid_161,{_zz_s1_outputPayload_selValid_160,{_zz_s1_outputPayload_selValid_159,{_zz_s1_outputPayload_selValid_158,{_zz_s1_outputPayload_selValid_157,{_zz_s1_outputPayload_selValid_156,{_zz_s1_outputPayload_selValid_1026,_zz_s1_outputPayload_selValid_1027}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1026 = _zz_s1_outputPayload_selValid_155;
  assign _zz_s1_outputPayload_selValid_1027 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h05));
  assign _zz_s1_outputPayload_selValid_1028 = _zz_s1_outputPayload_selValid_208;
  assign _zz_s1_outputPayload_selValid_1029 = {_zz_s1_outputPayload_selValid_207,{_zz_s1_outputPayload_selValid_206,{_zz_s1_outputPayload_selValid_205,{_zz_s1_outputPayload_selValid_204,{_zz_s1_outputPayload_selValid_203,{_zz_s1_outputPayload_selValid_202,{_zz_s1_outputPayload_selValid_201,{_zz_s1_outputPayload_selValid_200,{_zz_s1_outputPayload_selValid_199,{_zz_s1_outputPayload_selValid_198,{_zz_s1_outputPayload_selValid_1030,_zz_s1_outputPayload_selValid_1031}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1030 = _zz_s1_outputPayload_selValid_197;
  assign _zz_s1_outputPayload_selValid_1031 = {_zz_s1_outputPayload_selValid_196,{_zz_s1_outputPayload_selValid_195,{_zz_s1_outputPayload_selValid_194,{_zz_s1_outputPayload_selValid_193,{_zz_s1_outputPayload_selValid_192,{_zz_s1_outputPayload_selValid_191,{_zz_s1_outputPayload_selValid_190,{_zz_s1_outputPayload_selValid_189,{_zz_s1_outputPayload_selValid_188,{_zz_s1_outputPayload_selValid_187,{_zz_s1_outputPayload_selValid_1032,_zz_s1_outputPayload_selValid_1033}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1032 = _zz_s1_outputPayload_selValid_186;
  assign _zz_s1_outputPayload_selValid_1033 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h06));
  assign _zz_s1_outputPayload_selValid_1034 = _zz_s1_outputPayload_selValid_239;
  assign _zz_s1_outputPayload_selValid_1035 = {_zz_s1_outputPayload_selValid_238,{_zz_s1_outputPayload_selValid_237,{_zz_s1_outputPayload_selValid_236,{_zz_s1_outputPayload_selValid_235,{_zz_s1_outputPayload_selValid_234,{_zz_s1_outputPayload_selValid_233,{_zz_s1_outputPayload_selValid_232,{_zz_s1_outputPayload_selValid_231,{_zz_s1_outputPayload_selValid_230,{_zz_s1_outputPayload_selValid_229,{_zz_s1_outputPayload_selValid_1036,_zz_s1_outputPayload_selValid_1037}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1036 = _zz_s1_outputPayload_selValid_228;
  assign _zz_s1_outputPayload_selValid_1037 = {_zz_s1_outputPayload_selValid_227,{_zz_s1_outputPayload_selValid_226,{_zz_s1_outputPayload_selValid_225,{_zz_s1_outputPayload_selValid_224,{_zz_s1_outputPayload_selValid_223,{_zz_s1_outputPayload_selValid_222,{_zz_s1_outputPayload_selValid_221,{_zz_s1_outputPayload_selValid_220,{_zz_s1_outputPayload_selValid_219,{_zz_s1_outputPayload_selValid_218,{_zz_s1_outputPayload_selValid_1038,_zz_s1_outputPayload_selValid_1039}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1038 = _zz_s1_outputPayload_selValid_217;
  assign _zz_s1_outputPayload_selValid_1039 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h07));
  assign _zz_s1_outputPayload_selValid_1040 = _zz_s1_outputPayload_selValid_270;
  assign _zz_s1_outputPayload_selValid_1041 = {_zz_s1_outputPayload_selValid_269,{_zz_s1_outputPayload_selValid_268,{_zz_s1_outputPayload_selValid_267,{_zz_s1_outputPayload_selValid_266,{_zz_s1_outputPayload_selValid_265,{_zz_s1_outputPayload_selValid_264,{_zz_s1_outputPayload_selValid_263,{_zz_s1_outputPayload_selValid_262,{_zz_s1_outputPayload_selValid_261,{_zz_s1_outputPayload_selValid_260,{_zz_s1_outputPayload_selValid_1042,_zz_s1_outputPayload_selValid_1043}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1042 = _zz_s1_outputPayload_selValid_259;
  assign _zz_s1_outputPayload_selValid_1043 = {_zz_s1_outputPayload_selValid_258,{_zz_s1_outputPayload_selValid_257,{_zz_s1_outputPayload_selValid_256,{_zz_s1_outputPayload_selValid_255,{_zz_s1_outputPayload_selValid_254,{_zz_s1_outputPayload_selValid_253,{_zz_s1_outputPayload_selValid_252,{_zz_s1_outputPayload_selValid_251,{_zz_s1_outputPayload_selValid_250,{_zz_s1_outputPayload_selValid_249,{_zz_s1_outputPayload_selValid_1044,_zz_s1_outputPayload_selValid_1045}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1044 = _zz_s1_outputPayload_selValid_248;
  assign _zz_s1_outputPayload_selValid_1045 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h08));
  assign _zz_s1_outputPayload_selValid_1046 = _zz_s1_outputPayload_selValid_301;
  assign _zz_s1_outputPayload_selValid_1047 = {_zz_s1_outputPayload_selValid_300,{_zz_s1_outputPayload_selValid_299,{_zz_s1_outputPayload_selValid_298,{_zz_s1_outputPayload_selValid_297,{_zz_s1_outputPayload_selValid_296,{_zz_s1_outputPayload_selValid_295,{_zz_s1_outputPayload_selValid_294,{_zz_s1_outputPayload_selValid_293,{_zz_s1_outputPayload_selValid_292,{_zz_s1_outputPayload_selValid_291,{_zz_s1_outputPayload_selValid_1048,_zz_s1_outputPayload_selValid_1049}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1048 = _zz_s1_outputPayload_selValid_290;
  assign _zz_s1_outputPayload_selValid_1049 = {_zz_s1_outputPayload_selValid_289,{_zz_s1_outputPayload_selValid_288,{_zz_s1_outputPayload_selValid_287,{_zz_s1_outputPayload_selValid_286,{_zz_s1_outputPayload_selValid_285,{_zz_s1_outputPayload_selValid_284,{_zz_s1_outputPayload_selValid_283,{_zz_s1_outputPayload_selValid_282,{_zz_s1_outputPayload_selValid_281,{_zz_s1_outputPayload_selValid_280,{_zz_s1_outputPayload_selValid_1050,_zz_s1_outputPayload_selValid_1051}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1050 = _zz_s1_outputPayload_selValid_279;
  assign _zz_s1_outputPayload_selValid_1051 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h09));
  assign _zz_s1_outputPayload_selValid_1052 = _zz_s1_outputPayload_selValid_332;
  assign _zz_s1_outputPayload_selValid_1053 = {_zz_s1_outputPayload_selValid_331,{_zz_s1_outputPayload_selValid_330,{_zz_s1_outputPayload_selValid_329,{_zz_s1_outputPayload_selValid_328,{_zz_s1_outputPayload_selValid_327,{_zz_s1_outputPayload_selValid_326,{_zz_s1_outputPayload_selValid_325,{_zz_s1_outputPayload_selValid_324,{_zz_s1_outputPayload_selValid_323,{_zz_s1_outputPayload_selValid_322,{_zz_s1_outputPayload_selValid_1054,_zz_s1_outputPayload_selValid_1055}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1054 = _zz_s1_outputPayload_selValid_321;
  assign _zz_s1_outputPayload_selValid_1055 = {_zz_s1_outputPayload_selValid_320,{_zz_s1_outputPayload_selValid_319,{_zz_s1_outputPayload_selValid_318,{_zz_s1_outputPayload_selValid_317,{_zz_s1_outputPayload_selValid_316,{_zz_s1_outputPayload_selValid_315,{_zz_s1_outputPayload_selValid_314,{_zz_s1_outputPayload_selValid_313,{_zz_s1_outputPayload_selValid_312,{_zz_s1_outputPayload_selValid_311,{_zz_s1_outputPayload_selValid_1056,_zz_s1_outputPayload_selValid_1057}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1056 = _zz_s1_outputPayload_selValid_310;
  assign _zz_s1_outputPayload_selValid_1057 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_1058 = _zz_s1_outputPayload_selValid_363;
  assign _zz_s1_outputPayload_selValid_1059 = {_zz_s1_outputPayload_selValid_362,{_zz_s1_outputPayload_selValid_361,{_zz_s1_outputPayload_selValid_360,{_zz_s1_outputPayload_selValid_359,{_zz_s1_outputPayload_selValid_358,{_zz_s1_outputPayload_selValid_357,{_zz_s1_outputPayload_selValid_356,{_zz_s1_outputPayload_selValid_355,{_zz_s1_outputPayload_selValid_354,{_zz_s1_outputPayload_selValid_353,{_zz_s1_outputPayload_selValid_1060,_zz_s1_outputPayload_selValid_1061}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1060 = _zz_s1_outputPayload_selValid_352;
  assign _zz_s1_outputPayload_selValid_1061 = {_zz_s1_outputPayload_selValid_351,{_zz_s1_outputPayload_selValid_350,{_zz_s1_outputPayload_selValid_349,{_zz_s1_outputPayload_selValid_348,{_zz_s1_outputPayload_selValid_347,{_zz_s1_outputPayload_selValid_346,{_zz_s1_outputPayload_selValid_345,{_zz_s1_outputPayload_selValid_344,{_zz_s1_outputPayload_selValid_343,{_zz_s1_outputPayload_selValid_342,{_zz_s1_outputPayload_selValid_1062,_zz_s1_outputPayload_selValid_1063}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1062 = _zz_s1_outputPayload_selValid_341;
  assign _zz_s1_outputPayload_selValid_1063 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_1064 = _zz_s1_outputPayload_selValid_394;
  assign _zz_s1_outputPayload_selValid_1065 = {_zz_s1_outputPayload_selValid_393,{_zz_s1_outputPayload_selValid_392,{_zz_s1_outputPayload_selValid_391,{_zz_s1_outputPayload_selValid_390,{_zz_s1_outputPayload_selValid_389,{_zz_s1_outputPayload_selValid_388,{_zz_s1_outputPayload_selValid_387,{_zz_s1_outputPayload_selValid_386,{_zz_s1_outputPayload_selValid_385,{_zz_s1_outputPayload_selValid_384,{_zz_s1_outputPayload_selValid_1066,_zz_s1_outputPayload_selValid_1067}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1066 = _zz_s1_outputPayload_selValid_383;
  assign _zz_s1_outputPayload_selValid_1067 = {_zz_s1_outputPayload_selValid_382,{_zz_s1_outputPayload_selValid_381,{_zz_s1_outputPayload_selValid_380,{_zz_s1_outputPayload_selValid_379,{_zz_s1_outputPayload_selValid_378,{_zz_s1_outputPayload_selValid_377,{_zz_s1_outputPayload_selValid_376,{_zz_s1_outputPayload_selValid_375,{_zz_s1_outputPayload_selValid_374,{_zz_s1_outputPayload_selValid_373,{_zz_s1_outputPayload_selValid_1068,_zz_s1_outputPayload_selValid_1069}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1068 = _zz_s1_outputPayload_selValid_372;
  assign _zz_s1_outputPayload_selValid_1069 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_1070 = _zz_s1_outputPayload_selValid_425;
  assign _zz_s1_outputPayload_selValid_1071 = {_zz_s1_outputPayload_selValid_424,{_zz_s1_outputPayload_selValid_423,{_zz_s1_outputPayload_selValid_422,{_zz_s1_outputPayload_selValid_421,{_zz_s1_outputPayload_selValid_420,{_zz_s1_outputPayload_selValid_419,{_zz_s1_outputPayload_selValid_418,{_zz_s1_outputPayload_selValid_417,{_zz_s1_outputPayload_selValid_416,{_zz_s1_outputPayload_selValid_415,{_zz_s1_outputPayload_selValid_1072,_zz_s1_outputPayload_selValid_1073}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1072 = _zz_s1_outputPayload_selValid_414;
  assign _zz_s1_outputPayload_selValid_1073 = {_zz_s1_outputPayload_selValid_413,{_zz_s1_outputPayload_selValid_412,{_zz_s1_outputPayload_selValid_411,{_zz_s1_outputPayload_selValid_410,{_zz_s1_outputPayload_selValid_409,{_zz_s1_outputPayload_selValid_408,{_zz_s1_outputPayload_selValid_407,{_zz_s1_outputPayload_selValid_406,{_zz_s1_outputPayload_selValid_405,{_zz_s1_outputPayload_selValid_404,{_zz_s1_outputPayload_selValid_1074,_zz_s1_outputPayload_selValid_1075}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1074 = _zz_s1_outputPayload_selValid_403;
  assign _zz_s1_outputPayload_selValid_1075 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_1076 = _zz_s1_outputPayload_selValid_456;
  assign _zz_s1_outputPayload_selValid_1077 = {_zz_s1_outputPayload_selValid_455,{_zz_s1_outputPayload_selValid_454,{_zz_s1_outputPayload_selValid_453,{_zz_s1_outputPayload_selValid_452,{_zz_s1_outputPayload_selValid_451,{_zz_s1_outputPayload_selValid_450,{_zz_s1_outputPayload_selValid_449,{_zz_s1_outputPayload_selValid_448,{_zz_s1_outputPayload_selValid_447,{_zz_s1_outputPayload_selValid_446,{_zz_s1_outputPayload_selValid_1078,_zz_s1_outputPayload_selValid_1079}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1078 = _zz_s1_outputPayload_selValid_445;
  assign _zz_s1_outputPayload_selValid_1079 = {_zz_s1_outputPayload_selValid_444,{_zz_s1_outputPayload_selValid_443,{_zz_s1_outputPayload_selValid_442,{_zz_s1_outputPayload_selValid_441,{_zz_s1_outputPayload_selValid_440,{_zz_s1_outputPayload_selValid_439,{_zz_s1_outputPayload_selValid_438,{_zz_s1_outputPayload_selValid_437,{_zz_s1_outputPayload_selValid_436,{_zz_s1_outputPayload_selValid_435,{_zz_s1_outputPayload_selValid_1080,_zz_s1_outputPayload_selValid_1081}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1080 = _zz_s1_outputPayload_selValid_434;
  assign _zz_s1_outputPayload_selValid_1081 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_1082 = _zz_s1_outputPayload_selValid_487;
  assign _zz_s1_outputPayload_selValid_1083 = {_zz_s1_outputPayload_selValid_486,{_zz_s1_outputPayload_selValid_485,{_zz_s1_outputPayload_selValid_484,{_zz_s1_outputPayload_selValid_483,{_zz_s1_outputPayload_selValid_482,{_zz_s1_outputPayload_selValid_481,{_zz_s1_outputPayload_selValid_480,{_zz_s1_outputPayload_selValid_479,{_zz_s1_outputPayload_selValid_478,{_zz_s1_outputPayload_selValid_477,{_zz_s1_outputPayload_selValid_1084,_zz_s1_outputPayload_selValid_1085}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1084 = _zz_s1_outputPayload_selValid_476;
  assign _zz_s1_outputPayload_selValid_1085 = {_zz_s1_outputPayload_selValid_475,{_zz_s1_outputPayload_selValid_474,{_zz_s1_outputPayload_selValid_473,{_zz_s1_outputPayload_selValid_472,{_zz_s1_outputPayload_selValid_471,{_zz_s1_outputPayload_selValid_470,{_zz_s1_outputPayload_selValid_469,{_zz_s1_outputPayload_selValid_468,{_zz_s1_outputPayload_selValid_467,{_zz_s1_outputPayload_selValid_466,{_zz_s1_outputPayload_selValid_1086,_zz_s1_outputPayload_selValid_1087}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1086 = _zz_s1_outputPayload_selValid_465;
  assign _zz_s1_outputPayload_selValid_1087 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_1088 = _zz_s1_outputPayload_selValid_518;
  assign _zz_s1_outputPayload_selValid_1089 = {_zz_s1_outputPayload_selValid_517,{_zz_s1_outputPayload_selValid_516,{_zz_s1_outputPayload_selValid_515,{_zz_s1_outputPayload_selValid_514,{_zz_s1_outputPayload_selValid_513,{_zz_s1_outputPayload_selValid_512,{_zz_s1_outputPayload_selValid_511,{_zz_s1_outputPayload_selValid_510,{_zz_s1_outputPayload_selValid_509,{_zz_s1_outputPayload_selValid_508,{_zz_s1_outputPayload_selValid_1090,_zz_s1_outputPayload_selValid_1091}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1090 = _zz_s1_outputPayload_selValid_507;
  assign _zz_s1_outputPayload_selValid_1091 = {_zz_s1_outputPayload_selValid_506,{_zz_s1_outputPayload_selValid_505,{_zz_s1_outputPayload_selValid_504,{_zz_s1_outputPayload_selValid_503,{_zz_s1_outputPayload_selValid_502,{_zz_s1_outputPayload_selValid_501,{_zz_s1_outputPayload_selValid_500,{_zz_s1_outputPayload_selValid_499,{_zz_s1_outputPayload_selValid_498,{_zz_s1_outputPayload_selValid_497,{_zz_s1_outputPayload_selValid_1092,_zz_s1_outputPayload_selValid_1093}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1092 = _zz_s1_outputPayload_selValid_496;
  assign _zz_s1_outputPayload_selValid_1093 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h10));
  assign _zz_s1_outputPayload_selValid_1094 = _zz_s1_outputPayload_selValid_549;
  assign _zz_s1_outputPayload_selValid_1095 = {_zz_s1_outputPayload_selValid_548,{_zz_s1_outputPayload_selValid_547,{_zz_s1_outputPayload_selValid_546,{_zz_s1_outputPayload_selValid_545,{_zz_s1_outputPayload_selValid_544,{_zz_s1_outputPayload_selValid_543,{_zz_s1_outputPayload_selValid_542,{_zz_s1_outputPayload_selValid_541,{_zz_s1_outputPayload_selValid_540,{_zz_s1_outputPayload_selValid_539,{_zz_s1_outputPayload_selValid_1096,_zz_s1_outputPayload_selValid_1097}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1096 = _zz_s1_outputPayload_selValid_538;
  assign _zz_s1_outputPayload_selValid_1097 = {_zz_s1_outputPayload_selValid_537,{_zz_s1_outputPayload_selValid_536,{_zz_s1_outputPayload_selValid_535,{_zz_s1_outputPayload_selValid_534,{_zz_s1_outputPayload_selValid_533,{_zz_s1_outputPayload_selValid_532,{_zz_s1_outputPayload_selValid_531,{_zz_s1_outputPayload_selValid_530,{_zz_s1_outputPayload_selValid_529,{_zz_s1_outputPayload_selValid_528,{_zz_s1_outputPayload_selValid_1098,_zz_s1_outputPayload_selValid_1099}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1098 = _zz_s1_outputPayload_selValid_527;
  assign _zz_s1_outputPayload_selValid_1099 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h11));
  assign _zz_s1_outputPayload_selValid_1100 = _zz_s1_outputPayload_selValid_580;
  assign _zz_s1_outputPayload_selValid_1101 = {_zz_s1_outputPayload_selValid_579,{_zz_s1_outputPayload_selValid_578,{_zz_s1_outputPayload_selValid_577,{_zz_s1_outputPayload_selValid_576,{_zz_s1_outputPayload_selValid_575,{_zz_s1_outputPayload_selValid_574,{_zz_s1_outputPayload_selValid_573,{_zz_s1_outputPayload_selValid_572,{_zz_s1_outputPayload_selValid_571,{_zz_s1_outputPayload_selValid_570,{_zz_s1_outputPayload_selValid_1102,_zz_s1_outputPayload_selValid_1103}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1102 = _zz_s1_outputPayload_selValid_569;
  assign _zz_s1_outputPayload_selValid_1103 = {_zz_s1_outputPayload_selValid_568,{_zz_s1_outputPayload_selValid_567,{_zz_s1_outputPayload_selValid_566,{_zz_s1_outputPayload_selValid_565,{_zz_s1_outputPayload_selValid_564,{_zz_s1_outputPayload_selValid_563,{_zz_s1_outputPayload_selValid_562,{_zz_s1_outputPayload_selValid_561,{_zz_s1_outputPayload_selValid_560,{_zz_s1_outputPayload_selValid_559,{_zz_s1_outputPayload_selValid_1104,_zz_s1_outputPayload_selValid_1105}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1104 = _zz_s1_outputPayload_selValid_558;
  assign _zz_s1_outputPayload_selValid_1105 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h12));
  assign _zz_s1_outputPayload_selValid_1106 = _zz_s1_outputPayload_selValid_611;
  assign _zz_s1_outputPayload_selValid_1107 = {_zz_s1_outputPayload_selValid_610,{_zz_s1_outputPayload_selValid_609,{_zz_s1_outputPayload_selValid_608,{_zz_s1_outputPayload_selValid_607,{_zz_s1_outputPayload_selValid_606,{_zz_s1_outputPayload_selValid_605,{_zz_s1_outputPayload_selValid_604,{_zz_s1_outputPayload_selValid_603,{_zz_s1_outputPayload_selValid_602,{_zz_s1_outputPayload_selValid_601,{_zz_s1_outputPayload_selValid_1108,_zz_s1_outputPayload_selValid_1109}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1108 = _zz_s1_outputPayload_selValid_600;
  assign _zz_s1_outputPayload_selValid_1109 = {_zz_s1_outputPayload_selValid_599,{_zz_s1_outputPayload_selValid_598,{_zz_s1_outputPayload_selValid_597,{_zz_s1_outputPayload_selValid_596,{_zz_s1_outputPayload_selValid_595,{_zz_s1_outputPayload_selValid_594,{_zz_s1_outputPayload_selValid_593,{_zz_s1_outputPayload_selValid_592,{_zz_s1_outputPayload_selValid_591,{_zz_s1_outputPayload_selValid_590,{_zz_s1_outputPayload_selValid_1110,_zz_s1_outputPayload_selValid_1111}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1110 = _zz_s1_outputPayload_selValid_589;
  assign _zz_s1_outputPayload_selValid_1111 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h13));
  assign _zz_s1_outputPayload_selValid_1112 = _zz_s1_outputPayload_selValid_642;
  assign _zz_s1_outputPayload_selValid_1113 = {_zz_s1_outputPayload_selValid_641,{_zz_s1_outputPayload_selValid_640,{_zz_s1_outputPayload_selValid_639,{_zz_s1_outputPayload_selValid_638,{_zz_s1_outputPayload_selValid_637,{_zz_s1_outputPayload_selValid_636,{_zz_s1_outputPayload_selValid_635,{_zz_s1_outputPayload_selValid_634,{_zz_s1_outputPayload_selValid_633,{_zz_s1_outputPayload_selValid_632,{_zz_s1_outputPayload_selValid_1114,_zz_s1_outputPayload_selValid_1115}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1114 = _zz_s1_outputPayload_selValid_631;
  assign _zz_s1_outputPayload_selValid_1115 = {_zz_s1_outputPayload_selValid_630,{_zz_s1_outputPayload_selValid_629,{_zz_s1_outputPayload_selValid_628,{_zz_s1_outputPayload_selValid_627,{_zz_s1_outputPayload_selValid_626,{_zz_s1_outputPayload_selValid_625,{_zz_s1_outputPayload_selValid_624,{_zz_s1_outputPayload_selValid_623,{_zz_s1_outputPayload_selValid_622,{_zz_s1_outputPayload_selValid_621,{_zz_s1_outputPayload_selValid_1116,_zz_s1_outputPayload_selValid_1117}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1116 = _zz_s1_outputPayload_selValid_620;
  assign _zz_s1_outputPayload_selValid_1117 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h14));
  assign _zz_s1_outputPayload_selValid_1118 = _zz_s1_outputPayload_selValid_673;
  assign _zz_s1_outputPayload_selValid_1119 = {_zz_s1_outputPayload_selValid_672,{_zz_s1_outputPayload_selValid_671,{_zz_s1_outputPayload_selValid_670,{_zz_s1_outputPayload_selValid_669,{_zz_s1_outputPayload_selValid_668,{_zz_s1_outputPayload_selValid_667,{_zz_s1_outputPayload_selValid_666,{_zz_s1_outputPayload_selValid_665,{_zz_s1_outputPayload_selValid_664,{_zz_s1_outputPayload_selValid_663,{_zz_s1_outputPayload_selValid_1120,_zz_s1_outputPayload_selValid_1121}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1120 = _zz_s1_outputPayload_selValid_662;
  assign _zz_s1_outputPayload_selValid_1121 = {_zz_s1_outputPayload_selValid_661,{_zz_s1_outputPayload_selValid_660,{_zz_s1_outputPayload_selValid_659,{_zz_s1_outputPayload_selValid_658,{_zz_s1_outputPayload_selValid_657,{_zz_s1_outputPayload_selValid_656,{_zz_s1_outputPayload_selValid_655,{_zz_s1_outputPayload_selValid_654,{_zz_s1_outputPayload_selValid_653,{_zz_s1_outputPayload_selValid_652,{_zz_s1_outputPayload_selValid_1122,_zz_s1_outputPayload_selValid_1123}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1122 = _zz_s1_outputPayload_selValid_651;
  assign _zz_s1_outputPayload_selValid_1123 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h15));
  assign _zz_s1_outputPayload_selValid_1124 = _zz_s1_outputPayload_selValid_704;
  assign _zz_s1_outputPayload_selValid_1125 = {_zz_s1_outputPayload_selValid_703,{_zz_s1_outputPayload_selValid_702,{_zz_s1_outputPayload_selValid_701,{_zz_s1_outputPayload_selValid_700,{_zz_s1_outputPayload_selValid_699,{_zz_s1_outputPayload_selValid_698,{_zz_s1_outputPayload_selValid_697,{_zz_s1_outputPayload_selValid_696,{_zz_s1_outputPayload_selValid_695,{_zz_s1_outputPayload_selValid_694,{_zz_s1_outputPayload_selValid_1126,_zz_s1_outputPayload_selValid_1127}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1126 = _zz_s1_outputPayload_selValid_693;
  assign _zz_s1_outputPayload_selValid_1127 = {_zz_s1_outputPayload_selValid_692,{_zz_s1_outputPayload_selValid_691,{_zz_s1_outputPayload_selValid_690,{_zz_s1_outputPayload_selValid_689,{_zz_s1_outputPayload_selValid_688,{_zz_s1_outputPayload_selValid_687,{_zz_s1_outputPayload_selValid_686,{_zz_s1_outputPayload_selValid_685,{_zz_s1_outputPayload_selValid_684,{_zz_s1_outputPayload_selValid_683,{_zz_s1_outputPayload_selValid_1128,_zz_s1_outputPayload_selValid_1129}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1128 = _zz_s1_outputPayload_selValid_682;
  assign _zz_s1_outputPayload_selValid_1129 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h16));
  assign _zz_s1_outputPayload_selValid_1130 = _zz_s1_outputPayload_selValid_735;
  assign _zz_s1_outputPayload_selValid_1131 = {_zz_s1_outputPayload_selValid_734,{_zz_s1_outputPayload_selValid_733,{_zz_s1_outputPayload_selValid_732,{_zz_s1_outputPayload_selValid_731,{_zz_s1_outputPayload_selValid_730,{_zz_s1_outputPayload_selValid_729,{_zz_s1_outputPayload_selValid_728,{_zz_s1_outputPayload_selValid_727,{_zz_s1_outputPayload_selValid_726,{_zz_s1_outputPayload_selValid_725,{_zz_s1_outputPayload_selValid_1132,_zz_s1_outputPayload_selValid_1133}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1132 = _zz_s1_outputPayload_selValid_724;
  assign _zz_s1_outputPayload_selValid_1133 = {_zz_s1_outputPayload_selValid_723,{_zz_s1_outputPayload_selValid_722,{_zz_s1_outputPayload_selValid_721,{_zz_s1_outputPayload_selValid_720,{_zz_s1_outputPayload_selValid_719,{_zz_s1_outputPayload_selValid_718,{_zz_s1_outputPayload_selValid_717,{_zz_s1_outputPayload_selValid_716,{_zz_s1_outputPayload_selValid_715,{_zz_s1_outputPayload_selValid_714,{_zz_s1_outputPayload_selValid_1134,_zz_s1_outputPayload_selValid_1135}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1134 = _zz_s1_outputPayload_selValid_713;
  assign _zz_s1_outputPayload_selValid_1135 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h17));
  assign _zz_s1_outputPayload_selValid_1136 = _zz_s1_outputPayload_selValid_766;
  assign _zz_s1_outputPayload_selValid_1137 = {_zz_s1_outputPayload_selValid_765,{_zz_s1_outputPayload_selValid_764,{_zz_s1_outputPayload_selValid_763,{_zz_s1_outputPayload_selValid_762,{_zz_s1_outputPayload_selValid_761,{_zz_s1_outputPayload_selValid_760,{_zz_s1_outputPayload_selValid_759,{_zz_s1_outputPayload_selValid_758,{_zz_s1_outputPayload_selValid_757,{_zz_s1_outputPayload_selValid_756,{_zz_s1_outputPayload_selValid_1138,_zz_s1_outputPayload_selValid_1139}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1138 = _zz_s1_outputPayload_selValid_755;
  assign _zz_s1_outputPayload_selValid_1139 = {_zz_s1_outputPayload_selValid_754,{_zz_s1_outputPayload_selValid_753,{_zz_s1_outputPayload_selValid_752,{_zz_s1_outputPayload_selValid_751,{_zz_s1_outputPayload_selValid_750,{_zz_s1_outputPayload_selValid_749,{_zz_s1_outputPayload_selValid_748,{_zz_s1_outputPayload_selValid_747,{_zz_s1_outputPayload_selValid_746,{_zz_s1_outputPayload_selValid_745,{_zz_s1_outputPayload_selValid_1140,_zz_s1_outputPayload_selValid_1141}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1140 = _zz_s1_outputPayload_selValid_744;
  assign _zz_s1_outputPayload_selValid_1141 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h18));
  assign _zz_s1_outputPayload_selValid_1142 = _zz_s1_outputPayload_selValid_797;
  assign _zz_s1_outputPayload_selValid_1143 = {_zz_s1_outputPayload_selValid_796,{_zz_s1_outputPayload_selValid_795,{_zz_s1_outputPayload_selValid_794,{_zz_s1_outputPayload_selValid_793,{_zz_s1_outputPayload_selValid_792,{_zz_s1_outputPayload_selValid_791,{_zz_s1_outputPayload_selValid_790,{_zz_s1_outputPayload_selValid_789,{_zz_s1_outputPayload_selValid_788,{_zz_s1_outputPayload_selValid_787,{_zz_s1_outputPayload_selValid_1144,_zz_s1_outputPayload_selValid_1145}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1144 = _zz_s1_outputPayload_selValid_786;
  assign _zz_s1_outputPayload_selValid_1145 = {_zz_s1_outputPayload_selValid_785,{_zz_s1_outputPayload_selValid_784,{_zz_s1_outputPayload_selValid_783,{_zz_s1_outputPayload_selValid_782,{_zz_s1_outputPayload_selValid_781,{_zz_s1_outputPayload_selValid_780,{_zz_s1_outputPayload_selValid_779,{_zz_s1_outputPayload_selValid_778,{_zz_s1_outputPayload_selValid_777,{_zz_s1_outputPayload_selValid_776,{_zz_s1_outputPayload_selValid_1146,_zz_s1_outputPayload_selValid_1147}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1146 = _zz_s1_outputPayload_selValid_775;
  assign _zz_s1_outputPayload_selValid_1147 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h19));
  assign _zz_s1_outputPayload_selValid_1148 = _zz_s1_outputPayload_selValid_828;
  assign _zz_s1_outputPayload_selValid_1149 = {_zz_s1_outputPayload_selValid_827,{_zz_s1_outputPayload_selValid_826,{_zz_s1_outputPayload_selValid_825,{_zz_s1_outputPayload_selValid_824,{_zz_s1_outputPayload_selValid_823,{_zz_s1_outputPayload_selValid_822,{_zz_s1_outputPayload_selValid_821,{_zz_s1_outputPayload_selValid_820,{_zz_s1_outputPayload_selValid_819,{_zz_s1_outputPayload_selValid_818,{_zz_s1_outputPayload_selValid_1150,_zz_s1_outputPayload_selValid_1151}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1150 = _zz_s1_outputPayload_selValid_817;
  assign _zz_s1_outputPayload_selValid_1151 = {_zz_s1_outputPayload_selValid_816,{_zz_s1_outputPayload_selValid_815,{_zz_s1_outputPayload_selValid_814,{_zz_s1_outputPayload_selValid_813,{_zz_s1_outputPayload_selValid_812,{_zz_s1_outputPayload_selValid_811,{_zz_s1_outputPayload_selValid_810,{_zz_s1_outputPayload_selValid_809,{_zz_s1_outputPayload_selValid_808,{_zz_s1_outputPayload_selValid_807,{_zz_s1_outputPayload_selValid_1152,_zz_s1_outputPayload_selValid_1153}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1152 = _zz_s1_outputPayload_selValid_806;
  assign _zz_s1_outputPayload_selValid_1153 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_1154 = _zz_s1_outputPayload_selValid_859;
  assign _zz_s1_outputPayload_selValid_1155 = {_zz_s1_outputPayload_selValid_858,{_zz_s1_outputPayload_selValid_857,{_zz_s1_outputPayload_selValid_856,{_zz_s1_outputPayload_selValid_855,{_zz_s1_outputPayload_selValid_854,{_zz_s1_outputPayload_selValid_853,{_zz_s1_outputPayload_selValid_852,{_zz_s1_outputPayload_selValid_851,{_zz_s1_outputPayload_selValid_850,{_zz_s1_outputPayload_selValid_849,{_zz_s1_outputPayload_selValid_1156,_zz_s1_outputPayload_selValid_1157}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1156 = _zz_s1_outputPayload_selValid_848;
  assign _zz_s1_outputPayload_selValid_1157 = {_zz_s1_outputPayload_selValid_847,{_zz_s1_outputPayload_selValid_846,{_zz_s1_outputPayload_selValid_845,{_zz_s1_outputPayload_selValid_844,{_zz_s1_outputPayload_selValid_843,{_zz_s1_outputPayload_selValid_842,{_zz_s1_outputPayload_selValid_841,{_zz_s1_outputPayload_selValid_840,{_zz_s1_outputPayload_selValid_839,{_zz_s1_outputPayload_selValid_838,{_zz_s1_outputPayload_selValid_1158,_zz_s1_outputPayload_selValid_1159}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1158 = _zz_s1_outputPayload_selValid_837;
  assign _zz_s1_outputPayload_selValid_1159 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_1160 = _zz_s1_outputPayload_selValid_890;
  assign _zz_s1_outputPayload_selValid_1161 = {_zz_s1_outputPayload_selValid_889,{_zz_s1_outputPayload_selValid_888,{_zz_s1_outputPayload_selValid_887,{_zz_s1_outputPayload_selValid_886,{_zz_s1_outputPayload_selValid_885,{_zz_s1_outputPayload_selValid_884,{_zz_s1_outputPayload_selValid_883,{_zz_s1_outputPayload_selValid_882,{_zz_s1_outputPayload_selValid_881,{_zz_s1_outputPayload_selValid_880,{_zz_s1_outputPayload_selValid_1162,_zz_s1_outputPayload_selValid_1163}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1162 = _zz_s1_outputPayload_selValid_879;
  assign _zz_s1_outputPayload_selValid_1163 = {_zz_s1_outputPayload_selValid_878,{_zz_s1_outputPayload_selValid_877,{_zz_s1_outputPayload_selValid_876,{_zz_s1_outputPayload_selValid_875,{_zz_s1_outputPayload_selValid_874,{_zz_s1_outputPayload_selValid_873,{_zz_s1_outputPayload_selValid_872,{_zz_s1_outputPayload_selValid_871,{_zz_s1_outputPayload_selValid_870,{_zz_s1_outputPayload_selValid_869,{_zz_s1_outputPayload_selValid_1164,_zz_s1_outputPayload_selValid_1165}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1164 = _zz_s1_outputPayload_selValid_868;
  assign _zz_s1_outputPayload_selValid_1165 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_1166 = _zz_s1_outputPayload_selValid_921;
  assign _zz_s1_outputPayload_selValid_1167 = {_zz_s1_outputPayload_selValid_920,{_zz_s1_outputPayload_selValid_919,{_zz_s1_outputPayload_selValid_918,{_zz_s1_outputPayload_selValid_917,{_zz_s1_outputPayload_selValid_916,{_zz_s1_outputPayload_selValid_915,{_zz_s1_outputPayload_selValid_914,{_zz_s1_outputPayload_selValid_913,{_zz_s1_outputPayload_selValid_912,{_zz_s1_outputPayload_selValid_911,{_zz_s1_outputPayload_selValid_1168,_zz_s1_outputPayload_selValid_1169}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1168 = _zz_s1_outputPayload_selValid_910;
  assign _zz_s1_outputPayload_selValid_1169 = {_zz_s1_outputPayload_selValid_909,{_zz_s1_outputPayload_selValid_908,{_zz_s1_outputPayload_selValid_907,{_zz_s1_outputPayload_selValid_906,{_zz_s1_outputPayload_selValid_905,{_zz_s1_outputPayload_selValid_904,{_zz_s1_outputPayload_selValid_903,{_zz_s1_outputPayload_selValid_902,{_zz_s1_outputPayload_selValid_901,{_zz_s1_outputPayload_selValid_900,{_zz_s1_outputPayload_selValid_1170,_zz_s1_outputPayload_selValid_1171}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1170 = _zz_s1_outputPayload_selValid_899;
  assign _zz_s1_outputPayload_selValid_1171 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_1172 = _zz_s1_outputPayload_selValid_952;
  assign _zz_s1_outputPayload_selValid_1173 = {_zz_s1_outputPayload_selValid_951,{_zz_s1_outputPayload_selValid_950,{_zz_s1_outputPayload_selValid_949,{_zz_s1_outputPayload_selValid_948,{_zz_s1_outputPayload_selValid_947,{_zz_s1_outputPayload_selValid_946,{_zz_s1_outputPayload_selValid_945,{_zz_s1_outputPayload_selValid_944,{_zz_s1_outputPayload_selValid_943,{_zz_s1_outputPayload_selValid_942,{_zz_s1_outputPayload_selValid_1174,_zz_s1_outputPayload_selValid_1175}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1174 = _zz_s1_outputPayload_selValid_941;
  assign _zz_s1_outputPayload_selValid_1175 = {_zz_s1_outputPayload_selValid_940,{_zz_s1_outputPayload_selValid_939,{_zz_s1_outputPayload_selValid_938,{_zz_s1_outputPayload_selValid_937,{_zz_s1_outputPayload_selValid_936,{_zz_s1_outputPayload_selValid_935,{_zz_s1_outputPayload_selValid_934,{_zz_s1_outputPayload_selValid_933,{_zz_s1_outputPayload_selValid_932,{_zz_s1_outputPayload_selValid_931,{_zz_s1_outputPayload_selValid_1176,_zz_s1_outputPayload_selValid_1177}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1176 = _zz_s1_outputPayload_selValid_930;
  assign _zz_s1_outputPayload_selValid_1177 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_1178 = _zz_s1_outputPayload_selValid_983;
  assign _zz_s1_outputPayload_selValid_1179 = {_zz_s1_outputPayload_selValid_982,{_zz_s1_outputPayload_selValid_981,{_zz_s1_outputPayload_selValid_980,{_zz_s1_outputPayload_selValid_979,{_zz_s1_outputPayload_selValid_978,{_zz_s1_outputPayload_selValid_977,{_zz_s1_outputPayload_selValid_976,{_zz_s1_outputPayload_selValid_975,{_zz_s1_outputPayload_selValid_974,{_zz_s1_outputPayload_selValid_973,{_zz_s1_outputPayload_selValid_1180,_zz_s1_outputPayload_selValid_1181}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1180 = _zz_s1_outputPayload_selValid_972;
  assign _zz_s1_outputPayload_selValid_1181 = {_zz_s1_outputPayload_selValid_971,{_zz_s1_outputPayload_selValid_970,{_zz_s1_outputPayload_selValid_969,{_zz_s1_outputPayload_selValid_968,{_zz_s1_outputPayload_selValid_967,{_zz_s1_outputPayload_selValid_966,{_zz_s1_outputPayload_selValid_965,{_zz_s1_outputPayload_selValid_964,{_zz_s1_outputPayload_selValid_963,{_zz_s1_outputPayload_selValid_962,{_zz_s1_outputPayload_selValid_1182,_zz_s1_outputPayload_selValid_1183}}}}}}}}}}};
  assign _zz_s1_outputPayload_selValid_1182 = _zz_s1_outputPayload_selValid_961;
  assign _zz_s1_outputPayload_selValid_1183 = (s1_input_payload_cmd_mask[0] && (s1_inputIndexes_0 == 5'h1f));
  always @(*) begin
    case(_zz_s0_countOnesLogic_0_2)
      1'b0 : _zz_s0_countOnesLogic_0_1 = 1'b0;
      default : _zz_s0_countOnesLogic_0_1 = 1'b1;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_1_2)
      2'b00 : _zz_s0_countOnesLogic_1_1 = 2'b00;
      2'b01 : _zz_s0_countOnesLogic_1_1 = 2'b01;
      2'b10 : _zz_s0_countOnesLogic_1_1 = 2'b01;
      default : _zz_s0_countOnesLogic_1_1 = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_2_2)
      3'b000 : _zz_s0_countOnesLogic_2_1 = 2'b00;
      3'b001 : _zz_s0_countOnesLogic_2_1 = 2'b01;
      3'b010 : _zz_s0_countOnesLogic_2_1 = 2'b01;
      3'b011 : _zz_s0_countOnesLogic_2_1 = 2'b10;
      3'b100 : _zz_s0_countOnesLogic_2_1 = 2'b01;
      3'b101 : _zz_s0_countOnesLogic_2_1 = 2'b10;
      3'b110 : _zz_s0_countOnesLogic_2_1 = 2'b10;
      default : _zz_s0_countOnesLogic_2_1 = 2'b11;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_3_10)
      3'b000 : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_1;
      3'b001 : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_2;
      3'b010 : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_3;
      3'b011 : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_4;
      3'b100 : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_5;
      3'b101 : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_6;
      3'b110 : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_7;
      default : _zz_s0_countOnesLogic_3_9 = _zz_s0_countOnesLogic_3_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_3_12)
      3'b000 : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_1;
      3'b001 : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_2;
      3'b010 : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_3;
      3'b011 : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_4;
      3'b100 : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_5;
      3'b101 : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_6;
      3'b110 : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_7;
      default : _zz_s0_countOnesLogic_3_11 = _zz_s0_countOnesLogic_3_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_4_10)
      3'b000 : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_1;
      3'b001 : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_2;
      3'b010 : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_3;
      3'b011 : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_4;
      3'b100 : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_5;
      3'b101 : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_6;
      3'b110 : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_7;
      default : _zz_s0_countOnesLogic_4_9 = _zz_s0_countOnesLogic_4_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_4_12)
      3'b000 : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_1;
      3'b001 : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_2;
      3'b010 : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_3;
      3'b011 : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_4;
      3'b100 : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_5;
      3'b101 : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_6;
      3'b110 : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_7;
      default : _zz_s0_countOnesLogic_4_11 = _zz_s0_countOnesLogic_4_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_5_10)
      3'b000 : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_1;
      3'b001 : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_2;
      3'b010 : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_3;
      3'b011 : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_4;
      3'b100 : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_5;
      3'b101 : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_6;
      3'b110 : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_7;
      default : _zz_s0_countOnesLogic_5_9 = _zz_s0_countOnesLogic_5_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_5_12)
      3'b000 : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_1;
      3'b001 : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_2;
      3'b010 : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_3;
      3'b011 : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_4;
      3'b100 : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_5;
      3'b101 : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_6;
      3'b110 : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_7;
      default : _zz_s0_countOnesLogic_5_11 = _zz_s0_countOnesLogic_5_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_6_11)
      3'b000 : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_1;
      3'b001 : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_2;
      3'b010 : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_3;
      3'b011 : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_4;
      3'b100 : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_5;
      3'b101 : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_6;
      3'b110 : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_7;
      default : _zz_s0_countOnesLogic_6_10 = _zz_s0_countOnesLogic_6_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_6_13)
      3'b000 : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_1;
      3'b001 : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_2;
      3'b010 : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_3;
      3'b011 : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_4;
      3'b100 : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_5;
      3'b101 : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_6;
      3'b110 : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_7;
      default : _zz_s0_countOnesLogic_6_12 = _zz_s0_countOnesLogic_6_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_6_15)
      3'b000 : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_1;
      3'b001 : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_2;
      3'b010 : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_3;
      3'b011 : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_4;
      3'b100 : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_5;
      3'b101 : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_6;
      3'b110 : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_7;
      default : _zz_s0_countOnesLogic_6_14 = _zz_s0_countOnesLogic_6_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_7_11)
      3'b000 : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_1;
      3'b001 : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_2;
      3'b010 : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_3;
      3'b011 : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_4;
      3'b100 : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_5;
      3'b101 : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_6;
      3'b110 : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_7;
      default : _zz_s0_countOnesLogic_7_10 = _zz_s0_countOnesLogic_7_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_7_13)
      3'b000 : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_1;
      3'b001 : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_2;
      3'b010 : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_3;
      3'b011 : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_4;
      3'b100 : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_5;
      3'b101 : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_6;
      3'b110 : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_7;
      default : _zz_s0_countOnesLogic_7_12 = _zz_s0_countOnesLogic_7_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_7_15)
      3'b000 : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_1;
      3'b001 : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_2;
      3'b010 : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_3;
      3'b011 : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_4;
      3'b100 : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_5;
      3'b101 : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_6;
      3'b110 : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_7;
      default : _zz_s0_countOnesLogic_7_14 = _zz_s0_countOnesLogic_7_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_8_11)
      3'b000 : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_1;
      3'b001 : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_2;
      3'b010 : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_3;
      3'b011 : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_4;
      3'b100 : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_5;
      3'b101 : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_6;
      3'b110 : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_7;
      default : _zz_s0_countOnesLogic_8_10 = _zz_s0_countOnesLogic_8_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_8_13)
      3'b000 : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_1;
      3'b001 : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_2;
      3'b010 : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_3;
      3'b011 : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_4;
      3'b100 : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_5;
      3'b101 : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_6;
      3'b110 : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_7;
      default : _zz_s0_countOnesLogic_8_12 = _zz_s0_countOnesLogic_8_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_8_15)
      3'b000 : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_1;
      3'b001 : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_2;
      3'b010 : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_3;
      3'b011 : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_4;
      3'b100 : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_5;
      3'b101 : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_6;
      3'b110 : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_7;
      default : _zz_s0_countOnesLogic_8_14 = _zz_s0_countOnesLogic_8_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_9_11)
      3'b000 : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_1;
      3'b001 : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_2;
      3'b010 : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_3;
      3'b011 : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_4;
      3'b100 : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_5;
      3'b101 : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_6;
      3'b110 : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_7;
      default : _zz_s0_countOnesLogic_9_10 = _zz_s0_countOnesLogic_9_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_9_13)
      3'b000 : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_1;
      3'b001 : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_2;
      3'b010 : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_3;
      3'b011 : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_4;
      3'b100 : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_5;
      3'b101 : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_6;
      3'b110 : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_7;
      default : _zz_s0_countOnesLogic_9_12 = _zz_s0_countOnesLogic_9_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_9_16)
      3'b000 : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_1;
      3'b001 : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_2;
      3'b010 : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_3;
      3'b011 : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_4;
      3'b100 : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_5;
      3'b101 : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_6;
      3'b110 : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_7;
      default : _zz_s0_countOnesLogic_9_15 = _zz_s0_countOnesLogic_9_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_9_18)
      3'b000 : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_1;
      3'b001 : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_2;
      3'b010 : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_3;
      3'b011 : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_4;
      3'b100 : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_5;
      3'b101 : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_6;
      3'b110 : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_7;
      default : _zz_s0_countOnesLogic_9_17 = _zz_s0_countOnesLogic_9_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_10_11)
      3'b000 : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_1;
      3'b001 : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_2;
      3'b010 : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_3;
      3'b011 : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_4;
      3'b100 : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_5;
      3'b101 : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_6;
      3'b110 : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_7;
      default : _zz_s0_countOnesLogic_10_10 = _zz_s0_countOnesLogic_10_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_10_13)
      3'b000 : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_1;
      3'b001 : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_2;
      3'b010 : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_3;
      3'b011 : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_4;
      3'b100 : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_5;
      3'b101 : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_6;
      3'b110 : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_7;
      default : _zz_s0_countOnesLogic_10_12 = _zz_s0_countOnesLogic_10_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_10_16)
      3'b000 : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_1;
      3'b001 : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_2;
      3'b010 : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_3;
      3'b011 : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_4;
      3'b100 : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_5;
      3'b101 : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_6;
      3'b110 : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_7;
      default : _zz_s0_countOnesLogic_10_15 = _zz_s0_countOnesLogic_10_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_10_18)
      3'b000 : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_1;
      3'b001 : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_2;
      3'b010 : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_3;
      3'b011 : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_4;
      3'b100 : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_5;
      3'b101 : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_6;
      3'b110 : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_7;
      default : _zz_s0_countOnesLogic_10_17 = _zz_s0_countOnesLogic_10_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_11_11)
      3'b000 : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_1;
      3'b001 : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_2;
      3'b010 : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_3;
      3'b011 : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_4;
      3'b100 : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_5;
      3'b101 : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_6;
      3'b110 : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_7;
      default : _zz_s0_countOnesLogic_11_10 = _zz_s0_countOnesLogic_11_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_11_13)
      3'b000 : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_1;
      3'b001 : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_2;
      3'b010 : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_3;
      3'b011 : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_4;
      3'b100 : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_5;
      3'b101 : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_6;
      3'b110 : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_7;
      default : _zz_s0_countOnesLogic_11_12 = _zz_s0_countOnesLogic_11_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_11_16)
      3'b000 : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_1;
      3'b001 : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_2;
      3'b010 : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_3;
      3'b011 : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_4;
      3'b100 : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_5;
      3'b101 : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_6;
      3'b110 : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_7;
      default : _zz_s0_countOnesLogic_11_15 = _zz_s0_countOnesLogic_11_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_11_18)
      3'b000 : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_1;
      3'b001 : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_2;
      3'b010 : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_3;
      3'b011 : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_4;
      3'b100 : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_5;
      3'b101 : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_6;
      3'b110 : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_7;
      default : _zz_s0_countOnesLogic_11_17 = _zz_s0_countOnesLogic_11_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_12_12)
      3'b000 : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_1;
      3'b001 : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_2;
      3'b010 : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_3;
      3'b011 : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_4;
      3'b100 : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_5;
      3'b101 : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_6;
      3'b110 : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_7;
      default : _zz_s0_countOnesLogic_12_11 = _zz_s0_countOnesLogic_12_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_12_14)
      3'b000 : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_1;
      3'b001 : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_2;
      3'b010 : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_3;
      3'b011 : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_4;
      3'b100 : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_5;
      3'b101 : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_6;
      3'b110 : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_7;
      default : _zz_s0_countOnesLogic_12_13 = _zz_s0_countOnesLogic_12_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_12_17)
      3'b000 : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_1;
      3'b001 : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_2;
      3'b010 : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_3;
      3'b011 : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_4;
      3'b100 : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_5;
      3'b101 : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_6;
      3'b110 : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_7;
      default : _zz_s0_countOnesLogic_12_16 = _zz_s0_countOnesLogic_12_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_12_19)
      3'b000 : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_1;
      3'b001 : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_2;
      3'b010 : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_3;
      3'b011 : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_4;
      3'b100 : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_5;
      3'b101 : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_6;
      3'b110 : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_7;
      default : _zz_s0_countOnesLogic_12_18 = _zz_s0_countOnesLogic_12_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_12_21)
      3'b000 : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_1;
      3'b001 : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_2;
      3'b010 : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_3;
      3'b011 : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_4;
      3'b100 : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_5;
      3'b101 : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_6;
      3'b110 : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_7;
      default : _zz_s0_countOnesLogic_12_20 = _zz_s0_countOnesLogic_12_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_13_12)
      3'b000 : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_1;
      3'b001 : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_2;
      3'b010 : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_3;
      3'b011 : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_4;
      3'b100 : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_5;
      3'b101 : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_6;
      3'b110 : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_7;
      default : _zz_s0_countOnesLogic_13_11 = _zz_s0_countOnesLogic_13_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_13_14)
      3'b000 : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_1;
      3'b001 : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_2;
      3'b010 : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_3;
      3'b011 : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_4;
      3'b100 : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_5;
      3'b101 : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_6;
      3'b110 : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_7;
      default : _zz_s0_countOnesLogic_13_13 = _zz_s0_countOnesLogic_13_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_13_17)
      3'b000 : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_1;
      3'b001 : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_2;
      3'b010 : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_3;
      3'b011 : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_4;
      3'b100 : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_5;
      3'b101 : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_6;
      3'b110 : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_7;
      default : _zz_s0_countOnesLogic_13_16 = _zz_s0_countOnesLogic_13_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_13_19)
      3'b000 : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_1;
      3'b001 : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_2;
      3'b010 : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_3;
      3'b011 : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_4;
      3'b100 : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_5;
      3'b101 : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_6;
      3'b110 : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_7;
      default : _zz_s0_countOnesLogic_13_18 = _zz_s0_countOnesLogic_13_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_13_21)
      3'b000 : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_1;
      3'b001 : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_2;
      3'b010 : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_3;
      3'b011 : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_4;
      3'b100 : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_5;
      3'b101 : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_6;
      3'b110 : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_7;
      default : _zz_s0_countOnesLogic_13_20 = _zz_s0_countOnesLogic_13_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_14_12)
      3'b000 : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_1;
      3'b001 : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_2;
      3'b010 : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_3;
      3'b011 : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_4;
      3'b100 : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_5;
      3'b101 : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_6;
      3'b110 : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_7;
      default : _zz_s0_countOnesLogic_14_11 = _zz_s0_countOnesLogic_14_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_14_14)
      3'b000 : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_1;
      3'b001 : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_2;
      3'b010 : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_3;
      3'b011 : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_4;
      3'b100 : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_5;
      3'b101 : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_6;
      3'b110 : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_7;
      default : _zz_s0_countOnesLogic_14_13 = _zz_s0_countOnesLogic_14_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_14_17)
      3'b000 : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_1;
      3'b001 : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_2;
      3'b010 : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_3;
      3'b011 : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_4;
      3'b100 : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_5;
      3'b101 : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_6;
      3'b110 : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_7;
      default : _zz_s0_countOnesLogic_14_16 = _zz_s0_countOnesLogic_14_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_14_19)
      3'b000 : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_1;
      3'b001 : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_2;
      3'b010 : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_3;
      3'b011 : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_4;
      3'b100 : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_5;
      3'b101 : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_6;
      3'b110 : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_7;
      default : _zz_s0_countOnesLogic_14_18 = _zz_s0_countOnesLogic_14_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_14_21)
      3'b000 : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_1;
      3'b001 : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_2;
      3'b010 : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_3;
      3'b011 : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_4;
      3'b100 : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_5;
      3'b101 : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_6;
      3'b110 : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_7;
      default : _zz_s0_countOnesLogic_14_20 = _zz_s0_countOnesLogic_14_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_15_12)
      3'b000 : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_1;
      3'b001 : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_2;
      3'b010 : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_3;
      3'b011 : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_4;
      3'b100 : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_5;
      3'b101 : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_6;
      3'b110 : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_7;
      default : _zz_s0_countOnesLogic_15_11 = _zz_s0_countOnesLogic_15_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_15_14)
      3'b000 : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_1;
      3'b001 : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_2;
      3'b010 : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_3;
      3'b011 : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_4;
      3'b100 : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_5;
      3'b101 : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_6;
      3'b110 : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_7;
      default : _zz_s0_countOnesLogic_15_13 = _zz_s0_countOnesLogic_15_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_15_17)
      3'b000 : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_1;
      3'b001 : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_2;
      3'b010 : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_3;
      3'b011 : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_4;
      3'b100 : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_5;
      3'b101 : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_6;
      3'b110 : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_7;
      default : _zz_s0_countOnesLogic_15_16 = _zz_s0_countOnesLogic_15_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_15_19)
      3'b000 : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_1;
      3'b001 : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_2;
      3'b010 : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_3;
      3'b011 : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_4;
      3'b100 : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_5;
      3'b101 : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_6;
      3'b110 : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_7;
      default : _zz_s0_countOnesLogic_15_18 = _zz_s0_countOnesLogic_15_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_15_22)
      3'b000 : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_1;
      3'b001 : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_2;
      3'b010 : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_3;
      3'b011 : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_4;
      3'b100 : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_5;
      3'b101 : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_6;
      3'b110 : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_7;
      default : _zz_s0_countOnesLogic_15_21 = _zz_s0_countOnesLogic_15_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_15_24)
      3'b000 : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_1;
      3'b001 : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_2;
      3'b010 : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_3;
      3'b011 : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_4;
      3'b100 : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_5;
      3'b101 : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_6;
      3'b110 : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_7;
      default : _zz_s0_countOnesLogic_15_23 = _zz_s0_countOnesLogic_15_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_16_12)
      3'b000 : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_1;
      3'b001 : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_2;
      3'b010 : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_3;
      3'b011 : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_4;
      3'b100 : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_5;
      3'b101 : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_6;
      3'b110 : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_7;
      default : _zz_s0_countOnesLogic_16_11 = _zz_s0_countOnesLogic_16_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_16_14)
      3'b000 : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_1;
      3'b001 : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_2;
      3'b010 : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_3;
      3'b011 : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_4;
      3'b100 : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_5;
      3'b101 : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_6;
      3'b110 : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_7;
      default : _zz_s0_countOnesLogic_16_13 = _zz_s0_countOnesLogic_16_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_16_17)
      3'b000 : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_1;
      3'b001 : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_2;
      3'b010 : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_3;
      3'b011 : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_4;
      3'b100 : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_5;
      3'b101 : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_6;
      3'b110 : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_7;
      default : _zz_s0_countOnesLogic_16_16 = _zz_s0_countOnesLogic_16_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_16_19)
      3'b000 : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_1;
      3'b001 : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_2;
      3'b010 : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_3;
      3'b011 : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_4;
      3'b100 : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_5;
      3'b101 : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_6;
      3'b110 : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_7;
      default : _zz_s0_countOnesLogic_16_18 = _zz_s0_countOnesLogic_16_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_16_22)
      3'b000 : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_1;
      3'b001 : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_2;
      3'b010 : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_3;
      3'b011 : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_4;
      3'b100 : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_5;
      3'b101 : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_6;
      3'b110 : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_7;
      default : _zz_s0_countOnesLogic_16_21 = _zz_s0_countOnesLogic_16_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_16_24)
      3'b000 : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_1;
      3'b001 : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_2;
      3'b010 : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_3;
      3'b011 : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_4;
      3'b100 : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_5;
      3'b101 : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_6;
      3'b110 : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_7;
      default : _zz_s0_countOnesLogic_16_23 = _zz_s0_countOnesLogic_16_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_17_12)
      3'b000 : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_1;
      3'b001 : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_2;
      3'b010 : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_3;
      3'b011 : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_4;
      3'b100 : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_5;
      3'b101 : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_6;
      3'b110 : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_7;
      default : _zz_s0_countOnesLogic_17_11 = _zz_s0_countOnesLogic_17_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_17_14)
      3'b000 : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_1;
      3'b001 : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_2;
      3'b010 : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_3;
      3'b011 : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_4;
      3'b100 : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_5;
      3'b101 : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_6;
      3'b110 : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_7;
      default : _zz_s0_countOnesLogic_17_13 = _zz_s0_countOnesLogic_17_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_17_17)
      3'b000 : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_1;
      3'b001 : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_2;
      3'b010 : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_3;
      3'b011 : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_4;
      3'b100 : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_5;
      3'b101 : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_6;
      3'b110 : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_7;
      default : _zz_s0_countOnesLogic_17_16 = _zz_s0_countOnesLogic_17_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_17_19)
      3'b000 : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_1;
      3'b001 : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_2;
      3'b010 : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_3;
      3'b011 : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_4;
      3'b100 : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_5;
      3'b101 : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_6;
      3'b110 : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_7;
      default : _zz_s0_countOnesLogic_17_18 = _zz_s0_countOnesLogic_17_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_17_22)
      3'b000 : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_1;
      3'b001 : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_2;
      3'b010 : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_3;
      3'b011 : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_4;
      3'b100 : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_5;
      3'b101 : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_6;
      3'b110 : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_7;
      default : _zz_s0_countOnesLogic_17_21 = _zz_s0_countOnesLogic_17_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_17_24)
      3'b000 : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_1;
      3'b001 : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_2;
      3'b010 : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_3;
      3'b011 : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_4;
      3'b100 : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_5;
      3'b101 : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_6;
      3'b110 : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_7;
      default : _zz_s0_countOnesLogic_17_23 = _zz_s0_countOnesLogic_17_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_18_12)
      3'b000 : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_1;
      3'b001 : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_2;
      3'b010 : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_3;
      3'b011 : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_4;
      3'b100 : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_5;
      3'b101 : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_6;
      3'b110 : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_7;
      default : _zz_s0_countOnesLogic_18_11 = _zz_s0_countOnesLogic_18_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_18_14)
      3'b000 : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_1;
      3'b001 : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_2;
      3'b010 : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_3;
      3'b011 : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_4;
      3'b100 : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_5;
      3'b101 : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_6;
      3'b110 : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_7;
      default : _zz_s0_countOnesLogic_18_13 = _zz_s0_countOnesLogic_18_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_18_17)
      3'b000 : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_1;
      3'b001 : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_2;
      3'b010 : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_3;
      3'b011 : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_4;
      3'b100 : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_5;
      3'b101 : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_6;
      3'b110 : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_7;
      default : _zz_s0_countOnesLogic_18_16 = _zz_s0_countOnesLogic_18_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_18_19)
      3'b000 : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_1;
      3'b001 : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_2;
      3'b010 : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_3;
      3'b011 : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_4;
      3'b100 : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_5;
      3'b101 : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_6;
      3'b110 : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_7;
      default : _zz_s0_countOnesLogic_18_18 = _zz_s0_countOnesLogic_18_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_18_23)
      3'b000 : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_1;
      3'b001 : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_2;
      3'b010 : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_3;
      3'b011 : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_4;
      3'b100 : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_5;
      3'b101 : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_6;
      3'b110 : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_7;
      default : _zz_s0_countOnesLogic_18_22 = _zz_s0_countOnesLogic_18_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_18_25)
      3'b000 : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_1;
      3'b001 : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_2;
      3'b010 : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_3;
      3'b011 : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_4;
      3'b100 : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_5;
      3'b101 : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_6;
      3'b110 : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_7;
      default : _zz_s0_countOnesLogic_18_24 = _zz_s0_countOnesLogic_18_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_18_27)
      3'b000 : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_1;
      3'b001 : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_2;
      3'b010 : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_3;
      3'b011 : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_4;
      3'b100 : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_5;
      3'b101 : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_6;
      3'b110 : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_7;
      default : _zz_s0_countOnesLogic_18_26 = _zz_s0_countOnesLogic_18_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_19_12)
      3'b000 : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_1;
      3'b001 : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_2;
      3'b010 : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_3;
      3'b011 : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_4;
      3'b100 : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_5;
      3'b101 : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_6;
      3'b110 : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_7;
      default : _zz_s0_countOnesLogic_19_11 = _zz_s0_countOnesLogic_19_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_19_14)
      3'b000 : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_1;
      3'b001 : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_2;
      3'b010 : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_3;
      3'b011 : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_4;
      3'b100 : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_5;
      3'b101 : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_6;
      3'b110 : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_7;
      default : _zz_s0_countOnesLogic_19_13 = _zz_s0_countOnesLogic_19_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_19_17)
      3'b000 : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_1;
      3'b001 : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_2;
      3'b010 : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_3;
      3'b011 : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_4;
      3'b100 : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_5;
      3'b101 : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_6;
      3'b110 : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_7;
      default : _zz_s0_countOnesLogic_19_16 = _zz_s0_countOnesLogic_19_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_19_19)
      3'b000 : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_1;
      3'b001 : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_2;
      3'b010 : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_3;
      3'b011 : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_4;
      3'b100 : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_5;
      3'b101 : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_6;
      3'b110 : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_7;
      default : _zz_s0_countOnesLogic_19_18 = _zz_s0_countOnesLogic_19_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_19_23)
      3'b000 : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_1;
      3'b001 : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_2;
      3'b010 : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_3;
      3'b011 : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_4;
      3'b100 : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_5;
      3'b101 : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_6;
      3'b110 : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_7;
      default : _zz_s0_countOnesLogic_19_22 = _zz_s0_countOnesLogic_19_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_19_25)
      3'b000 : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_1;
      3'b001 : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_2;
      3'b010 : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_3;
      3'b011 : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_4;
      3'b100 : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_5;
      3'b101 : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_6;
      3'b110 : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_7;
      default : _zz_s0_countOnesLogic_19_24 = _zz_s0_countOnesLogic_19_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_19_27)
      3'b000 : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_1;
      3'b001 : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_2;
      3'b010 : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_3;
      3'b011 : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_4;
      3'b100 : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_5;
      3'b101 : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_6;
      3'b110 : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_7;
      default : _zz_s0_countOnesLogic_19_26 = _zz_s0_countOnesLogic_19_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_20_12)
      3'b000 : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_1;
      3'b001 : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_2;
      3'b010 : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_3;
      3'b011 : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_4;
      3'b100 : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_5;
      3'b101 : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_6;
      3'b110 : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_7;
      default : _zz_s0_countOnesLogic_20_11 = _zz_s0_countOnesLogic_20_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_20_14)
      3'b000 : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_1;
      3'b001 : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_2;
      3'b010 : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_3;
      3'b011 : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_4;
      3'b100 : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_5;
      3'b101 : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_6;
      3'b110 : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_7;
      default : _zz_s0_countOnesLogic_20_13 = _zz_s0_countOnesLogic_20_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_20_17)
      3'b000 : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_1;
      3'b001 : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_2;
      3'b010 : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_3;
      3'b011 : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_4;
      3'b100 : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_5;
      3'b101 : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_6;
      3'b110 : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_7;
      default : _zz_s0_countOnesLogic_20_16 = _zz_s0_countOnesLogic_20_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_20_19)
      3'b000 : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_1;
      3'b001 : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_2;
      3'b010 : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_3;
      3'b011 : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_4;
      3'b100 : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_5;
      3'b101 : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_6;
      3'b110 : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_7;
      default : _zz_s0_countOnesLogic_20_18 = _zz_s0_countOnesLogic_20_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_20_23)
      3'b000 : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_1;
      3'b001 : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_2;
      3'b010 : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_3;
      3'b011 : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_4;
      3'b100 : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_5;
      3'b101 : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_6;
      3'b110 : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_7;
      default : _zz_s0_countOnesLogic_20_22 = _zz_s0_countOnesLogic_20_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_20_25)
      3'b000 : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_1;
      3'b001 : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_2;
      3'b010 : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_3;
      3'b011 : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_4;
      3'b100 : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_5;
      3'b101 : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_6;
      3'b110 : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_7;
      default : _zz_s0_countOnesLogic_20_24 = _zz_s0_countOnesLogic_20_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_20_27)
      3'b000 : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_1;
      3'b001 : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_2;
      3'b010 : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_3;
      3'b011 : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_4;
      3'b100 : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_5;
      3'b101 : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_6;
      3'b110 : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_7;
      default : _zz_s0_countOnesLogic_20_26 = _zz_s0_countOnesLogic_20_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_12)
      3'b000 : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_11 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_14)
      3'b000 : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_13 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_17)
      3'b000 : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_16 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_19)
      3'b000 : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_18 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_23)
      3'b000 : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_22 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_25)
      3'b000 : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_24 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_28)
      3'b000 : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_27 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_21_30)
      3'b000 : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_1;
      3'b001 : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_2;
      3'b010 : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_3;
      3'b011 : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_4;
      3'b100 : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_5;
      3'b101 : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_6;
      3'b110 : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_7;
      default : _zz_s0_countOnesLogic_21_29 = _zz_s0_countOnesLogic_21_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_12)
      3'b000 : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_11 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_14)
      3'b000 : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_13 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_17)
      3'b000 : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_16 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_19)
      3'b000 : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_18 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_23)
      3'b000 : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_22 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_25)
      3'b000 : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_24 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_28)
      3'b000 : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_27 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_22_30)
      3'b000 : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_1;
      3'b001 : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_2;
      3'b010 : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_3;
      3'b011 : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_4;
      3'b100 : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_5;
      3'b101 : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_6;
      3'b110 : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_7;
      default : _zz_s0_countOnesLogic_22_29 = _zz_s0_countOnesLogic_22_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_12)
      3'b000 : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_11 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_14)
      3'b000 : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_13 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_17)
      3'b000 : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_16 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_19)
      3'b000 : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_18 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_23)
      3'b000 : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_22 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_25)
      3'b000 : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_24 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_28)
      3'b000 : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_27 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_23_30)
      3'b000 : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_1;
      3'b001 : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_2;
      3'b010 : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_3;
      3'b011 : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_4;
      3'b100 : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_5;
      3'b101 : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_6;
      3'b110 : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_7;
      default : _zz_s0_countOnesLogic_23_29 = _zz_s0_countOnesLogic_23_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_13)
      3'b000 : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_12 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_15)
      3'b000 : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_14 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_18)
      3'b000 : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_17 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_20)
      3'b000 : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_19 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_24)
      3'b000 : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_23 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_26)
      3'b000 : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_25 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_29)
      3'b000 : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_28 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_31)
      3'b000 : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_30 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_24_33)
      3'b000 : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_1;
      3'b001 : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_2;
      3'b010 : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_3;
      3'b011 : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_4;
      3'b100 : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_5;
      3'b101 : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_6;
      3'b110 : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_7;
      default : _zz_s0_countOnesLogic_24_32 = _zz_s0_countOnesLogic_24_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_13)
      3'b000 : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_12 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_15)
      3'b000 : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_14 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_18)
      3'b000 : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_17 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_20)
      3'b000 : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_19 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_24)
      3'b000 : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_23 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_26)
      3'b000 : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_25 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_29)
      3'b000 : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_28 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_31)
      3'b000 : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_30 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_25_33)
      3'b000 : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_1;
      3'b001 : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_2;
      3'b010 : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_3;
      3'b011 : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_4;
      3'b100 : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_5;
      3'b101 : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_6;
      3'b110 : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_7;
      default : _zz_s0_countOnesLogic_25_32 = _zz_s0_countOnesLogic_25_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_13)
      3'b000 : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_12 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_15)
      3'b000 : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_14 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_18)
      3'b000 : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_17 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_20)
      3'b000 : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_19 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_24)
      3'b000 : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_23 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_26)
      3'b000 : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_25 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_29)
      3'b000 : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_28 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_31)
      3'b000 : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_30 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_26_33)
      3'b000 : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_1;
      3'b001 : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_2;
      3'b010 : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_3;
      3'b011 : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_4;
      3'b100 : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_5;
      3'b101 : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_6;
      3'b110 : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_7;
      default : _zz_s0_countOnesLogic_26_32 = _zz_s0_countOnesLogic_26_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_13)
      3'b000 : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_12 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_15)
      3'b000 : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_14 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_18)
      3'b000 : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_17 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_20)
      3'b000 : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_19 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_24)
      3'b000 : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_23 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_26)
      3'b000 : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_25 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_29)
      3'b000 : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_28 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_31)
      3'b000 : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_30 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_34)
      3'b000 : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_33 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_27_36)
      3'b000 : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_1;
      3'b001 : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_2;
      3'b010 : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_3;
      3'b011 : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_4;
      3'b100 : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_5;
      3'b101 : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_6;
      3'b110 : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_7;
      default : _zz_s0_countOnesLogic_27_35 = _zz_s0_countOnesLogic_27_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_13)
      3'b000 : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_12 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_15)
      3'b000 : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_14 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_18)
      3'b000 : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_17 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_20)
      3'b000 : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_19 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_24)
      3'b000 : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_23 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_26)
      3'b000 : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_25 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_29)
      3'b000 : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_28 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_31)
      3'b000 : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_30 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_34)
      3'b000 : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_33 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_28_36)
      3'b000 : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_1;
      3'b001 : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_2;
      3'b010 : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_3;
      3'b011 : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_4;
      3'b100 : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_5;
      3'b101 : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_6;
      3'b110 : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_7;
      default : _zz_s0_countOnesLogic_28_35 = _zz_s0_countOnesLogic_28_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_13)
      3'b000 : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_12 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_15)
      3'b000 : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_14 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_18)
      3'b000 : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_17 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_20)
      3'b000 : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_19 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_24)
      3'b000 : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_23 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_26)
      3'b000 : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_25 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_29)
      3'b000 : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_28 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_31)
      3'b000 : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_30 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_34)
      3'b000 : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_33 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_29_36)
      3'b000 : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_1;
      3'b001 : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_2;
      3'b010 : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_3;
      3'b011 : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_4;
      3'b100 : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_5;
      3'b101 : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_6;
      3'b110 : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_7;
      default : _zz_s0_countOnesLogic_29_35 = _zz_s0_countOnesLogic_29_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_13)
      3'b000 : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_12 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_15)
      3'b000 : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_14 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_18)
      3'b000 : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_17 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_20)
      3'b000 : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_19 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_24)
      3'b000 : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_23 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_26)
      3'b000 : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_25 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_29)
      3'b000 : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_28 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_31)
      3'b000 : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_30 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_35)
      3'b000 : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_34 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_37)
      3'b000 : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_36 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_30_39)
      3'b000 : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_1;
      3'b001 : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_2;
      3'b010 : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_3;
      3'b011 : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_4;
      3'b100 : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_5;
      3'b101 : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_6;
      3'b110 : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_7;
      default : _zz_s0_countOnesLogic_30_38 = _zz_s0_countOnesLogic_30_8;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_12)
      3'b000 : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_11 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_14)
      3'b000 : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_13 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_17)
      3'b000 : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_16 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_19)
      3'b000 : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_18 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_23)
      3'b000 : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_22 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_25)
      3'b000 : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_24 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_28)
      3'b000 : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_27 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_30)
      3'b000 : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_29 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_34)
      3'b000 : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_33 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_36)
      3'b000 : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_35 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(_zz_s0_countOnesLogic_31_38)
      3'b000 : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31;
      3'b001 : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31_1;
      3'b010 : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31_2;
      3'b011 : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31_3;
      3'b100 : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31_4;
      3'b101 : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31_5;
      3'b110 : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31_6;
      default : _zz_s0_countOnesLogic_31_37 = _zz_s0_countOnesLogic_31_7;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_0)
      5'b00000 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_0_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_1)
      5'b00000 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_1_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_2)
      5'b00000 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_2_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_3)
      5'b00000 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_3_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_4)
      5'b00000 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_4_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_5)
      5'b00000 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_5_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_6)
      5'b00000 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_6_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_7)
      5'b00000 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_7_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_8)
      5'b00000 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_8_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_9)
      5'b00000 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_9_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_10)
      5'b00000 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_10_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_11)
      5'b00000 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_11_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_12)
      5'b00000 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_12_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_13)
      5'b00000 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_13_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_14)
      5'b00000 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_14_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_15)
      5'b00000 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_15_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_16)
      5'b00000 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_16_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_17)
      5'b00000 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_17_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_18)
      5'b00000 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_18_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_19)
      5'b00000 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_19_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_20)
      5'b00000 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_20_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_21)
      5'b00000 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_21_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_22)
      5'b00000 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_22_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_23)
      5'b00000 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_23_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_24)
      5'b00000 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_24_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_25)
      5'b00000 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_25_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_26)
      5'b00000 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_26_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_27)
      5'b00000 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_27_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_28)
      5'b00000 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_28_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_29)
      5'b00000 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_29_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_30)
      5'b00000 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_30_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(s2_input_payload_sel_31)
      5'b00000 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_0;
      5'b00001 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_1;
      5'b00010 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_2;
      5'b00011 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_3;
      5'b00100 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_4;
      5'b00101 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_5;
      5'b00110 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_6;
      5'b00111 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_7;
      5'b01000 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_8;
      5'b01001 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_9;
      5'b01010 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_10;
      5'b01011 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_11;
      5'b01100 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_12;
      5'b01101 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_13;
      5'b01110 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_14;
      5'b01111 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_15;
      5'b10000 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_16;
      5'b10001 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_17;
      5'b10010 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_18;
      5'b10011 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_19;
      5'b10100 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_20;
      5'b10101 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_21;
      5'b10110 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_22;
      5'b10111 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_23;
      5'b11000 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_24;
      5'b11001 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_25;
      5'b11010 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_26;
      5'b11011 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_27;
      5'b11100 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_28;
      5'b11101 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_29;
      5'b11110 : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_30;
      default : _zz_s2_byteLogic_31_inputData = s2_inputDataBytes_31;
    endcase
  end

  always @(*) begin
    case(_zz_io_output_usedUntil_6)
      5'b00000 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_0;
      5'b00001 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_1;
      5'b00010 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_2;
      5'b00011 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_3;
      5'b00100 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_4;
      5'b00101 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_5;
      5'b00110 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_6;
      5'b00111 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_7;
      5'b01000 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_8;
      5'b01001 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_9;
      5'b01010 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_10;
      5'b01011 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_11;
      5'b01100 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_12;
      5'b01101 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_13;
      5'b01110 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_14;
      5'b01111 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_15;
      5'b10000 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_16;
      5'b10001 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_17;
      5'b10010 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_18;
      5'b10011 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_19;
      5'b10100 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_20;
      5'b10101 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_21;
      5'b10110 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_22;
      5'b10111 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_23;
      5'b11000 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_24;
      5'b11001 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_25;
      5'b11010 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_26;
      5'b11011 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_27;
      5'b11100 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_28;
      5'b11101 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_29;
      5'b11110 : _zz_io_output_usedUntil_5 = s2_input_payload_sel_30;
      default : _zz_io_output_usedUntil_5 = s2_input_payload_sel_31;
    endcase
  end

  always @(*) begin
    io_input_ready = s0_input_ready;
    if(when_Stream_l375) begin
      io_input_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! s0_input_valid);
  assign s0_input_valid = io_input_rValid;
  assign s0_input_payload_data = io_input_rData_data;
  assign s0_input_payload_mask = io_input_rData_mask;
  assign _zz_s0_countOnesLogic_0 = s0_input_payload_mask[0];
  assign _zz_s0_countOnesLogic_1 = s0_input_payload_mask[1];
  assign _zz_s0_countOnesLogic_2 = s0_input_payload_mask[2];
  assign _zz_s0_countOnesLogic_3 = s0_input_payload_mask[3];
  assign _zz_s0_countOnesLogic_4 = s0_input_payload_mask[4];
  assign _zz_s0_countOnesLogic_5 = s0_input_payload_mask[5];
  assign _zz_s0_countOnesLogic_6 = s0_input_payload_mask[6];
  assign _zz_s0_countOnesLogic_7 = s0_input_payload_mask[7];
  assign _zz_s0_countOnesLogic_8 = s0_input_payload_mask[8];
  assign _zz_s0_countOnesLogic_9 = s0_input_payload_mask[9];
  assign _zz_s0_countOnesLogic_10 = s0_input_payload_mask[10];
  assign _zz_s0_countOnesLogic_11 = s0_input_payload_mask[11];
  assign _zz_s0_countOnesLogic_12 = s0_input_payload_mask[12];
  assign _zz_s0_countOnesLogic_13 = s0_input_payload_mask[13];
  assign _zz_s0_countOnesLogic_14 = s0_input_payload_mask[14];
  assign _zz_s0_countOnesLogic_15 = s0_input_payload_mask[15];
  assign _zz_s0_countOnesLogic_16 = s0_input_payload_mask[16];
  assign _zz_s0_countOnesLogic_17 = s0_input_payload_mask[17];
  assign _zz_s0_countOnesLogic_18 = s0_input_payload_mask[18];
  assign _zz_s0_countOnesLogic_19 = s0_input_payload_mask[19];
  assign _zz_s0_countOnesLogic_20 = s0_input_payload_mask[20];
  assign _zz_s0_countOnesLogic_21 = s0_input_payload_mask[21];
  assign _zz_s0_countOnesLogic_22 = s0_input_payload_mask[22];
  assign _zz_s0_countOnesLogic_23 = s0_input_payload_mask[23];
  assign _zz_s0_countOnesLogic_24 = s0_input_payload_mask[24];
  assign _zz_s0_countOnesLogic_25 = s0_input_payload_mask[25];
  assign _zz_s0_countOnesLogic_26 = s0_input_payload_mask[26];
  assign _zz_s0_countOnesLogic_27 = s0_input_payload_mask[27];
  assign _zz_s0_countOnesLogic_28 = s0_input_payload_mask[28];
  assign _zz_s0_countOnesLogic_29 = s0_input_payload_mask[29];
  assign _zz_s0_countOnesLogic_30 = s0_input_payload_mask[30];
  assign s0_countOnesLogic_0 = _zz_s0_countOnesLogic_0_1;
  assign s0_countOnesLogic_1 = _zz_s0_countOnesLogic_1_1;
  assign s0_countOnesLogic_2 = _zz_s0_countOnesLogic_2_1;
  assign _zz_s0_countOnesLogic_3_1 = 3'b000;
  assign _zz_s0_countOnesLogic_3_2 = 3'b001;
  assign _zz_s0_countOnesLogic_3_3 = 3'b001;
  assign _zz_s0_countOnesLogic_3_4 = 3'b010;
  assign _zz_s0_countOnesLogic_3_5 = 3'b001;
  assign _zz_s0_countOnesLogic_3_6 = 3'b010;
  assign _zz_s0_countOnesLogic_3_7 = 3'b010;
  assign _zz_s0_countOnesLogic_3_8 = 3'b011;
  assign s0_countOnesLogic_3 = (_zz_s0_countOnesLogic_3_9 + _zz_s0_countOnesLogic_3_11);
  assign _zz_s0_countOnesLogic_4_1 = 3'b000;
  assign _zz_s0_countOnesLogic_4_2 = 3'b001;
  assign _zz_s0_countOnesLogic_4_3 = 3'b001;
  assign _zz_s0_countOnesLogic_4_4 = 3'b010;
  assign _zz_s0_countOnesLogic_4_5 = 3'b001;
  assign _zz_s0_countOnesLogic_4_6 = 3'b010;
  assign _zz_s0_countOnesLogic_4_7 = 3'b010;
  assign _zz_s0_countOnesLogic_4_8 = 3'b011;
  assign s0_countOnesLogic_4 = (_zz_s0_countOnesLogic_4_9 + _zz_s0_countOnesLogic_4_11);
  assign _zz_s0_countOnesLogic_5_1 = 3'b000;
  assign _zz_s0_countOnesLogic_5_2 = 3'b001;
  assign _zz_s0_countOnesLogic_5_3 = 3'b001;
  assign _zz_s0_countOnesLogic_5_4 = 3'b010;
  assign _zz_s0_countOnesLogic_5_5 = 3'b001;
  assign _zz_s0_countOnesLogic_5_6 = 3'b010;
  assign _zz_s0_countOnesLogic_5_7 = 3'b010;
  assign _zz_s0_countOnesLogic_5_8 = 3'b011;
  assign s0_countOnesLogic_5 = (_zz_s0_countOnesLogic_5_9 + _zz_s0_countOnesLogic_5_11);
  assign _zz_s0_countOnesLogic_6_1 = 3'b000;
  assign _zz_s0_countOnesLogic_6_2 = 3'b001;
  assign _zz_s0_countOnesLogic_6_3 = 3'b001;
  assign _zz_s0_countOnesLogic_6_4 = 3'b010;
  assign _zz_s0_countOnesLogic_6_5 = 3'b001;
  assign _zz_s0_countOnesLogic_6_6 = 3'b010;
  assign _zz_s0_countOnesLogic_6_7 = 3'b010;
  assign _zz_s0_countOnesLogic_6_8 = 3'b011;
  assign s0_countOnesLogic_6 = (_zz_s0_countOnesLogic_6_9 + _zz_s0_countOnesLogic_6_14);
  assign _zz_s0_countOnesLogic_7_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_7_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_7_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_7_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_7_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_7_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_7_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_7_8 = 4'b0011;
  assign s0_countOnesLogic_7 = (_zz_s0_countOnesLogic_7_9 + _zz_s0_countOnesLogic_7_14);
  assign _zz_s0_countOnesLogic_8_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_8_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_8_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_8_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_8_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_8_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_8_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_8_8 = 4'b0011;
  assign s0_countOnesLogic_8 = (_zz_s0_countOnesLogic_8_9 + _zz_s0_countOnesLogic_8_14);
  assign _zz_s0_countOnesLogic_9_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_9_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_9_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_9_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_9_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_9_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_9_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_9_8 = 4'b0011;
  assign s0_countOnesLogic_9 = (_zz_s0_countOnesLogic_9_9 + _zz_s0_countOnesLogic_9_14);
  assign _zz_s0_countOnesLogic_10_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_10_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_10_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_10_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_10_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_10_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_10_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_10_8 = 4'b0011;
  assign s0_countOnesLogic_10 = (_zz_s0_countOnesLogic_10_9 + _zz_s0_countOnesLogic_10_14);
  assign _zz_s0_countOnesLogic_11_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_11_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_11_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_11_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_11_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_11_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_11_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_11_8 = 4'b0011;
  assign s0_countOnesLogic_11 = (_zz_s0_countOnesLogic_11_9 + _zz_s0_countOnesLogic_11_14);
  assign _zz_s0_countOnesLogic_12_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_12_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_12_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_12_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_12_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_12_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_12_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_12_8 = 4'b0011;
  assign s0_countOnesLogic_12 = (_zz_s0_countOnesLogic_12_9 + _zz_s0_countOnesLogic_12_20);
  assign _zz_s0_countOnesLogic_13_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_13_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_13_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_13_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_13_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_13_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_13_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_13_8 = 4'b0011;
  assign s0_countOnesLogic_13 = (_zz_s0_countOnesLogic_13_9 + _zz_s0_countOnesLogic_13_20);
  assign _zz_s0_countOnesLogic_14_1 = 4'b0000;
  assign _zz_s0_countOnesLogic_14_2 = 4'b0001;
  assign _zz_s0_countOnesLogic_14_3 = 4'b0001;
  assign _zz_s0_countOnesLogic_14_4 = 4'b0010;
  assign _zz_s0_countOnesLogic_14_5 = 4'b0001;
  assign _zz_s0_countOnesLogic_14_6 = 4'b0010;
  assign _zz_s0_countOnesLogic_14_7 = 4'b0010;
  assign _zz_s0_countOnesLogic_14_8 = 4'b0011;
  assign s0_countOnesLogic_14 = (_zz_s0_countOnesLogic_14_9 + _zz_s0_countOnesLogic_14_20);
  assign _zz_s0_countOnesLogic_15_1 = 5'h0;
  assign _zz_s0_countOnesLogic_15_2 = 5'h01;
  assign _zz_s0_countOnesLogic_15_3 = 5'h01;
  assign _zz_s0_countOnesLogic_15_4 = 5'h02;
  assign _zz_s0_countOnesLogic_15_5 = 5'h01;
  assign _zz_s0_countOnesLogic_15_6 = 5'h02;
  assign _zz_s0_countOnesLogic_15_7 = 5'h02;
  assign _zz_s0_countOnesLogic_15_8 = 5'h03;
  assign s0_countOnesLogic_15 = (_zz_s0_countOnesLogic_15_9 + _zz_s0_countOnesLogic_15_20);
  assign _zz_s0_countOnesLogic_16_1 = 5'h0;
  assign _zz_s0_countOnesLogic_16_2 = 5'h01;
  assign _zz_s0_countOnesLogic_16_3 = 5'h01;
  assign _zz_s0_countOnesLogic_16_4 = 5'h02;
  assign _zz_s0_countOnesLogic_16_5 = 5'h01;
  assign _zz_s0_countOnesLogic_16_6 = 5'h02;
  assign _zz_s0_countOnesLogic_16_7 = 5'h02;
  assign _zz_s0_countOnesLogic_16_8 = 5'h03;
  assign s0_countOnesLogic_16 = (_zz_s0_countOnesLogic_16_9 + _zz_s0_countOnesLogic_16_20);
  assign _zz_s0_countOnesLogic_17_1 = 5'h0;
  assign _zz_s0_countOnesLogic_17_2 = 5'h01;
  assign _zz_s0_countOnesLogic_17_3 = 5'h01;
  assign _zz_s0_countOnesLogic_17_4 = 5'h02;
  assign _zz_s0_countOnesLogic_17_5 = 5'h01;
  assign _zz_s0_countOnesLogic_17_6 = 5'h02;
  assign _zz_s0_countOnesLogic_17_7 = 5'h02;
  assign _zz_s0_countOnesLogic_17_8 = 5'h03;
  assign s0_countOnesLogic_17 = (_zz_s0_countOnesLogic_17_9 + _zz_s0_countOnesLogic_17_20);
  assign _zz_s0_countOnesLogic_18_1 = 5'h0;
  assign _zz_s0_countOnesLogic_18_2 = 5'h01;
  assign _zz_s0_countOnesLogic_18_3 = 5'h01;
  assign _zz_s0_countOnesLogic_18_4 = 5'h02;
  assign _zz_s0_countOnesLogic_18_5 = 5'h01;
  assign _zz_s0_countOnesLogic_18_6 = 5'h02;
  assign _zz_s0_countOnesLogic_18_7 = 5'h02;
  assign _zz_s0_countOnesLogic_18_8 = 5'h03;
  assign s0_countOnesLogic_18 = (_zz_s0_countOnesLogic_18_9 + _zz_s0_countOnesLogic_18_20);
  assign _zz_s0_countOnesLogic_19_1 = 5'h0;
  assign _zz_s0_countOnesLogic_19_2 = 5'h01;
  assign _zz_s0_countOnesLogic_19_3 = 5'h01;
  assign _zz_s0_countOnesLogic_19_4 = 5'h02;
  assign _zz_s0_countOnesLogic_19_5 = 5'h01;
  assign _zz_s0_countOnesLogic_19_6 = 5'h02;
  assign _zz_s0_countOnesLogic_19_7 = 5'h02;
  assign _zz_s0_countOnesLogic_19_8 = 5'h03;
  assign s0_countOnesLogic_19 = (_zz_s0_countOnesLogic_19_9 + _zz_s0_countOnesLogic_19_20);
  assign _zz_s0_countOnesLogic_20_1 = 5'h0;
  assign _zz_s0_countOnesLogic_20_2 = 5'h01;
  assign _zz_s0_countOnesLogic_20_3 = 5'h01;
  assign _zz_s0_countOnesLogic_20_4 = 5'h02;
  assign _zz_s0_countOnesLogic_20_5 = 5'h01;
  assign _zz_s0_countOnesLogic_20_6 = 5'h02;
  assign _zz_s0_countOnesLogic_20_7 = 5'h02;
  assign _zz_s0_countOnesLogic_20_8 = 5'h03;
  assign s0_countOnesLogic_20 = (_zz_s0_countOnesLogic_20_9 + _zz_s0_countOnesLogic_20_20);
  assign _zz_s0_countOnesLogic_21_1 = 5'h0;
  assign _zz_s0_countOnesLogic_21_2 = 5'h01;
  assign _zz_s0_countOnesLogic_21_3 = 5'h01;
  assign _zz_s0_countOnesLogic_21_4 = 5'h02;
  assign _zz_s0_countOnesLogic_21_5 = 5'h01;
  assign _zz_s0_countOnesLogic_21_6 = 5'h02;
  assign _zz_s0_countOnesLogic_21_7 = 5'h02;
  assign _zz_s0_countOnesLogic_21_8 = 5'h03;
  assign s0_countOnesLogic_21 = (_zz_s0_countOnesLogic_21_9 + _zz_s0_countOnesLogic_21_20);
  assign _zz_s0_countOnesLogic_22_1 = 5'h0;
  assign _zz_s0_countOnesLogic_22_2 = 5'h01;
  assign _zz_s0_countOnesLogic_22_3 = 5'h01;
  assign _zz_s0_countOnesLogic_22_4 = 5'h02;
  assign _zz_s0_countOnesLogic_22_5 = 5'h01;
  assign _zz_s0_countOnesLogic_22_6 = 5'h02;
  assign _zz_s0_countOnesLogic_22_7 = 5'h02;
  assign _zz_s0_countOnesLogic_22_8 = 5'h03;
  assign s0_countOnesLogic_22 = (_zz_s0_countOnesLogic_22_9 + _zz_s0_countOnesLogic_22_20);
  assign _zz_s0_countOnesLogic_23_1 = 5'h0;
  assign _zz_s0_countOnesLogic_23_2 = 5'h01;
  assign _zz_s0_countOnesLogic_23_3 = 5'h01;
  assign _zz_s0_countOnesLogic_23_4 = 5'h02;
  assign _zz_s0_countOnesLogic_23_5 = 5'h01;
  assign _zz_s0_countOnesLogic_23_6 = 5'h02;
  assign _zz_s0_countOnesLogic_23_7 = 5'h02;
  assign _zz_s0_countOnesLogic_23_8 = 5'h03;
  assign s0_countOnesLogic_23 = (_zz_s0_countOnesLogic_23_9 + _zz_s0_countOnesLogic_23_20);
  assign _zz_s0_countOnesLogic_24_1 = 5'h0;
  assign _zz_s0_countOnesLogic_24_2 = 5'h01;
  assign _zz_s0_countOnesLogic_24_3 = 5'h01;
  assign _zz_s0_countOnesLogic_24_4 = 5'h02;
  assign _zz_s0_countOnesLogic_24_5 = 5'h01;
  assign _zz_s0_countOnesLogic_24_6 = 5'h02;
  assign _zz_s0_countOnesLogic_24_7 = 5'h02;
  assign _zz_s0_countOnesLogic_24_8 = 5'h03;
  assign s0_countOnesLogic_24 = (_zz_s0_countOnesLogic_24_9 + _zz_s0_countOnesLogic_24_32);
  assign _zz_s0_countOnesLogic_25_1 = 5'h0;
  assign _zz_s0_countOnesLogic_25_2 = 5'h01;
  assign _zz_s0_countOnesLogic_25_3 = 5'h01;
  assign _zz_s0_countOnesLogic_25_4 = 5'h02;
  assign _zz_s0_countOnesLogic_25_5 = 5'h01;
  assign _zz_s0_countOnesLogic_25_6 = 5'h02;
  assign _zz_s0_countOnesLogic_25_7 = 5'h02;
  assign _zz_s0_countOnesLogic_25_8 = 5'h03;
  assign s0_countOnesLogic_25 = (_zz_s0_countOnesLogic_25_9 + _zz_s0_countOnesLogic_25_32);
  assign _zz_s0_countOnesLogic_26_1 = 5'h0;
  assign _zz_s0_countOnesLogic_26_2 = 5'h01;
  assign _zz_s0_countOnesLogic_26_3 = 5'h01;
  assign _zz_s0_countOnesLogic_26_4 = 5'h02;
  assign _zz_s0_countOnesLogic_26_5 = 5'h01;
  assign _zz_s0_countOnesLogic_26_6 = 5'h02;
  assign _zz_s0_countOnesLogic_26_7 = 5'h02;
  assign _zz_s0_countOnesLogic_26_8 = 5'h03;
  assign s0_countOnesLogic_26 = (_zz_s0_countOnesLogic_26_9 + _zz_s0_countOnesLogic_26_32);
  assign _zz_s0_countOnesLogic_27_1 = 5'h0;
  assign _zz_s0_countOnesLogic_27_2 = 5'h01;
  assign _zz_s0_countOnesLogic_27_3 = 5'h01;
  assign _zz_s0_countOnesLogic_27_4 = 5'h02;
  assign _zz_s0_countOnesLogic_27_5 = 5'h01;
  assign _zz_s0_countOnesLogic_27_6 = 5'h02;
  assign _zz_s0_countOnesLogic_27_7 = 5'h02;
  assign _zz_s0_countOnesLogic_27_8 = 5'h03;
  assign s0_countOnesLogic_27 = (_zz_s0_countOnesLogic_27_9 + _zz_s0_countOnesLogic_27_32);
  assign _zz_s0_countOnesLogic_28_1 = 5'h0;
  assign _zz_s0_countOnesLogic_28_2 = 5'h01;
  assign _zz_s0_countOnesLogic_28_3 = 5'h01;
  assign _zz_s0_countOnesLogic_28_4 = 5'h02;
  assign _zz_s0_countOnesLogic_28_5 = 5'h01;
  assign _zz_s0_countOnesLogic_28_6 = 5'h02;
  assign _zz_s0_countOnesLogic_28_7 = 5'h02;
  assign _zz_s0_countOnesLogic_28_8 = 5'h03;
  assign s0_countOnesLogic_28 = (_zz_s0_countOnesLogic_28_9 + _zz_s0_countOnesLogic_28_32);
  assign _zz_s0_countOnesLogic_29_1 = 5'h0;
  assign _zz_s0_countOnesLogic_29_2 = 5'h01;
  assign _zz_s0_countOnesLogic_29_3 = 5'h01;
  assign _zz_s0_countOnesLogic_29_4 = 5'h02;
  assign _zz_s0_countOnesLogic_29_5 = 5'h01;
  assign _zz_s0_countOnesLogic_29_6 = 5'h02;
  assign _zz_s0_countOnesLogic_29_7 = 5'h02;
  assign _zz_s0_countOnesLogic_29_8 = 5'h03;
  assign s0_countOnesLogic_29 = (_zz_s0_countOnesLogic_29_9 + _zz_s0_countOnesLogic_29_32);
  assign _zz_s0_countOnesLogic_30_1 = 5'h0;
  assign _zz_s0_countOnesLogic_30_2 = 5'h01;
  assign _zz_s0_countOnesLogic_30_3 = 5'h01;
  assign _zz_s0_countOnesLogic_30_4 = 5'h02;
  assign _zz_s0_countOnesLogic_30_5 = 5'h01;
  assign _zz_s0_countOnesLogic_30_6 = 5'h02;
  assign _zz_s0_countOnesLogic_30_7 = 5'h02;
  assign _zz_s0_countOnesLogic_30_8 = 5'h03;
  assign s0_countOnesLogic_30 = (_zz_s0_countOnesLogic_30_9 + _zz_s0_countOnesLogic_30_32);
  assign _zz_s0_countOnesLogic_31 = 6'h0;
  assign _zz_s0_countOnesLogic_31_1 = 6'h01;
  assign _zz_s0_countOnesLogic_31_2 = 6'h01;
  assign _zz_s0_countOnesLogic_31_3 = 6'h02;
  assign _zz_s0_countOnesLogic_31_4 = 6'h01;
  assign _zz_s0_countOnesLogic_31_5 = 6'h02;
  assign _zz_s0_countOnesLogic_31_6 = 6'h02;
  assign _zz_s0_countOnesLogic_31_7 = 6'h03;
  assign s0_countOnesLogic_31 = (_zz_s0_countOnesLogic_31_8 + _zz_s0_countOnesLogic_31_31);
  assign s0_outputPayload_cmd_data = s0_input_payload_data;
  assign s0_outputPayload_cmd_mask = s0_input_payload_mask;
  assign s0_outputPayload_countOnes_0 = s0_countOnesLogic_0;
  assign s0_outputPayload_countOnes_1 = s0_countOnesLogic_1;
  assign s0_outputPayload_countOnes_2 = s0_countOnesLogic_2;
  assign s0_outputPayload_countOnes_3 = s0_countOnesLogic_3;
  assign s0_outputPayload_countOnes_4 = s0_countOnesLogic_4;
  assign s0_outputPayload_countOnes_5 = s0_countOnesLogic_5;
  assign s0_outputPayload_countOnes_6 = s0_countOnesLogic_6;
  assign s0_outputPayload_countOnes_7 = s0_countOnesLogic_7;
  assign s0_outputPayload_countOnes_8 = s0_countOnesLogic_8;
  assign s0_outputPayload_countOnes_9 = s0_countOnesLogic_9;
  assign s0_outputPayload_countOnes_10 = s0_countOnesLogic_10;
  assign s0_outputPayload_countOnes_11 = s0_countOnesLogic_11;
  assign s0_outputPayload_countOnes_12 = s0_countOnesLogic_12;
  assign s0_outputPayload_countOnes_13 = s0_countOnesLogic_13;
  assign s0_outputPayload_countOnes_14 = s0_countOnesLogic_14;
  assign s0_outputPayload_countOnes_15 = s0_countOnesLogic_15;
  assign s0_outputPayload_countOnes_16 = s0_countOnesLogic_16;
  assign s0_outputPayload_countOnes_17 = s0_countOnesLogic_17;
  assign s0_outputPayload_countOnes_18 = s0_countOnesLogic_18;
  assign s0_outputPayload_countOnes_19 = s0_countOnesLogic_19;
  assign s0_outputPayload_countOnes_20 = s0_countOnesLogic_20;
  assign s0_outputPayload_countOnes_21 = s0_countOnesLogic_21;
  assign s0_outputPayload_countOnes_22 = s0_countOnesLogic_22;
  assign s0_outputPayload_countOnes_23 = s0_countOnesLogic_23;
  assign s0_outputPayload_countOnes_24 = s0_countOnesLogic_24;
  assign s0_outputPayload_countOnes_25 = s0_countOnesLogic_25;
  assign s0_outputPayload_countOnes_26 = s0_countOnesLogic_26;
  assign s0_outputPayload_countOnes_27 = s0_countOnesLogic_27;
  assign s0_outputPayload_countOnes_28 = s0_countOnesLogic_28;
  assign s0_outputPayload_countOnes_29 = s0_countOnesLogic_29;
  assign s0_outputPayload_countOnes_30 = s0_countOnesLogic_30;
  assign s0_outputPayload_countOnes_31 = s0_countOnesLogic_31;
  assign s0_output_valid = s0_input_valid;
  assign s0_input_ready = s0_output_ready;
  assign s0_output_payload_cmd_data = s0_outputPayload_cmd_data;
  assign s0_output_payload_cmd_mask = s0_outputPayload_cmd_mask;
  assign s0_output_payload_countOnes_0 = s0_outputPayload_countOnes_0;
  assign s0_output_payload_countOnes_1 = s0_outputPayload_countOnes_1;
  assign s0_output_payload_countOnes_2 = s0_outputPayload_countOnes_2;
  assign s0_output_payload_countOnes_3 = s0_outputPayload_countOnes_3;
  assign s0_output_payload_countOnes_4 = s0_outputPayload_countOnes_4;
  assign s0_output_payload_countOnes_5 = s0_outputPayload_countOnes_5;
  assign s0_output_payload_countOnes_6 = s0_outputPayload_countOnes_6;
  assign s0_output_payload_countOnes_7 = s0_outputPayload_countOnes_7;
  assign s0_output_payload_countOnes_8 = s0_outputPayload_countOnes_8;
  assign s0_output_payload_countOnes_9 = s0_outputPayload_countOnes_9;
  assign s0_output_payload_countOnes_10 = s0_outputPayload_countOnes_10;
  assign s0_output_payload_countOnes_11 = s0_outputPayload_countOnes_11;
  assign s0_output_payload_countOnes_12 = s0_outputPayload_countOnes_12;
  assign s0_output_payload_countOnes_13 = s0_outputPayload_countOnes_13;
  assign s0_output_payload_countOnes_14 = s0_outputPayload_countOnes_14;
  assign s0_output_payload_countOnes_15 = s0_outputPayload_countOnes_15;
  assign s0_output_payload_countOnes_16 = s0_outputPayload_countOnes_16;
  assign s0_output_payload_countOnes_17 = s0_outputPayload_countOnes_17;
  assign s0_output_payload_countOnes_18 = s0_outputPayload_countOnes_18;
  assign s0_output_payload_countOnes_19 = s0_outputPayload_countOnes_19;
  assign s0_output_payload_countOnes_20 = s0_outputPayload_countOnes_20;
  assign s0_output_payload_countOnes_21 = s0_outputPayload_countOnes_21;
  assign s0_output_payload_countOnes_22 = s0_outputPayload_countOnes_22;
  assign s0_output_payload_countOnes_23 = s0_outputPayload_countOnes_23;
  assign s0_output_payload_countOnes_24 = s0_outputPayload_countOnes_24;
  assign s0_output_payload_countOnes_25 = s0_outputPayload_countOnes_25;
  assign s0_output_payload_countOnes_26 = s0_outputPayload_countOnes_26;
  assign s0_output_payload_countOnes_27 = s0_outputPayload_countOnes_27;
  assign s0_output_payload_countOnes_28 = s0_outputPayload_countOnes_28;
  assign s0_output_payload_countOnes_29 = s0_outputPayload_countOnes_29;
  assign s0_output_payload_countOnes_30 = s0_outputPayload_countOnes_30;
  assign s0_output_payload_countOnes_31 = s0_outputPayload_countOnes_31;
  always @(*) begin
    s0_output_ready = s1_input_ready;
    if(when_Stream_l375_1) begin
      s0_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! s1_input_valid);
  assign s1_input_valid = s0_output_rValid;
  assign s1_input_payload_cmd_data = s0_output_rData_cmd_data;
  assign s1_input_payload_cmd_mask = s0_output_rData_cmd_mask;
  assign s1_input_payload_countOnes_0 = s0_output_rData_countOnes_0;
  assign s1_input_payload_countOnes_1 = s0_output_rData_countOnes_1;
  assign s1_input_payload_countOnes_2 = s0_output_rData_countOnes_2;
  assign s1_input_payload_countOnes_3 = s0_output_rData_countOnes_3;
  assign s1_input_payload_countOnes_4 = s0_output_rData_countOnes_4;
  assign s1_input_payload_countOnes_5 = s0_output_rData_countOnes_5;
  assign s1_input_payload_countOnes_6 = s0_output_rData_countOnes_6;
  assign s1_input_payload_countOnes_7 = s0_output_rData_countOnes_7;
  assign s1_input_payload_countOnes_8 = s0_output_rData_countOnes_8;
  assign s1_input_payload_countOnes_9 = s0_output_rData_countOnes_9;
  assign s1_input_payload_countOnes_10 = s0_output_rData_countOnes_10;
  assign s1_input_payload_countOnes_11 = s0_output_rData_countOnes_11;
  assign s1_input_payload_countOnes_12 = s0_output_rData_countOnes_12;
  assign s1_input_payload_countOnes_13 = s0_output_rData_countOnes_13;
  assign s1_input_payload_countOnes_14 = s0_output_rData_countOnes_14;
  assign s1_input_payload_countOnes_15 = s0_output_rData_countOnes_15;
  assign s1_input_payload_countOnes_16 = s0_output_rData_countOnes_16;
  assign s1_input_payload_countOnes_17 = s0_output_rData_countOnes_17;
  assign s1_input_payload_countOnes_18 = s0_output_rData_countOnes_18;
  assign s1_input_payload_countOnes_19 = s0_output_rData_countOnes_19;
  assign s1_input_payload_countOnes_20 = s0_output_rData_countOnes_20;
  assign s1_input_payload_countOnes_21 = s0_output_rData_countOnes_21;
  assign s1_input_payload_countOnes_22 = s0_output_rData_countOnes_22;
  assign s1_input_payload_countOnes_23 = s0_output_rData_countOnes_23;
  assign s1_input_payload_countOnes_24 = s0_output_rData_countOnes_24;
  assign s1_input_payload_countOnes_25 = s0_output_rData_countOnes_25;
  assign s1_input_payload_countOnes_26 = s0_output_rData_countOnes_26;
  assign s1_input_payload_countOnes_27 = s0_output_rData_countOnes_27;
  assign s1_input_payload_countOnes_28 = s0_output_rData_countOnes_28;
  assign s1_input_payload_countOnes_29 = s0_output_rData_countOnes_29;
  assign s1_input_payload_countOnes_30 = s0_output_rData_countOnes_30;
  assign s1_input_payload_countOnes_31 = s0_output_rData_countOnes_31;
  assign s1_offsetNext = (_zz_s1_offsetNext + s1_input_payload_countOnes_31);
  assign s1_input_fire = (s1_input_valid && s1_input_ready);
  assign s1_inputIndexes_0 = (5'h0 + s1_offset);
  assign s1_inputIndexes_1 = (_zz_s1_inputIndexes_1 + s1_offset);
  assign s1_inputIndexes_2 = (_zz_s1_inputIndexes_2 + s1_offset);
  assign s1_inputIndexes_3 = (_zz_s1_inputIndexes_3 + s1_offset);
  assign s1_inputIndexes_4 = (_zz_s1_inputIndexes_4 + s1_offset);
  assign s1_inputIndexes_5 = (_zz_s1_inputIndexes_5 + s1_offset);
  assign s1_inputIndexes_6 = (_zz_s1_inputIndexes_6 + s1_offset);
  assign s1_inputIndexes_7 = (_zz_s1_inputIndexes_7 + s1_offset);
  assign s1_inputIndexes_8 = (_zz_s1_inputIndexes_8 + s1_offset);
  assign s1_inputIndexes_9 = (_zz_s1_inputIndexes_9 + s1_offset);
  assign s1_inputIndexes_10 = (_zz_s1_inputIndexes_10 + s1_offset);
  assign s1_inputIndexes_11 = (_zz_s1_inputIndexes_11 + s1_offset);
  assign s1_inputIndexes_12 = (_zz_s1_inputIndexes_12 + s1_offset);
  assign s1_inputIndexes_13 = (_zz_s1_inputIndexes_13 + s1_offset);
  assign s1_inputIndexes_14 = (_zz_s1_inputIndexes_14 + s1_offset);
  assign s1_inputIndexes_15 = (_zz_s1_inputIndexes_15 + s1_offset);
  assign s1_inputIndexes_16 = (s1_input_payload_countOnes_15 + s1_offset);
  assign s1_inputIndexes_17 = (s1_input_payload_countOnes_16 + s1_offset);
  assign s1_inputIndexes_18 = (s1_input_payload_countOnes_17 + s1_offset);
  assign s1_inputIndexes_19 = (s1_input_payload_countOnes_18 + s1_offset);
  assign s1_inputIndexes_20 = (s1_input_payload_countOnes_19 + s1_offset);
  assign s1_inputIndexes_21 = (s1_input_payload_countOnes_20 + s1_offset);
  assign s1_inputIndexes_22 = (s1_input_payload_countOnes_21 + s1_offset);
  assign s1_inputIndexes_23 = (s1_input_payload_countOnes_22 + s1_offset);
  assign s1_inputIndexes_24 = (s1_input_payload_countOnes_23 + s1_offset);
  assign s1_inputIndexes_25 = (s1_input_payload_countOnes_24 + s1_offset);
  assign s1_inputIndexes_26 = (s1_input_payload_countOnes_25 + s1_offset);
  assign s1_inputIndexes_27 = (s1_input_payload_countOnes_26 + s1_offset);
  assign s1_inputIndexes_28 = (s1_input_payload_countOnes_27 + s1_offset);
  assign s1_inputIndexes_29 = (s1_input_payload_countOnes_28 + s1_offset);
  assign s1_inputIndexes_30 = (s1_input_payload_countOnes_29 + s1_offset);
  assign s1_inputIndexes_31 = (s1_input_payload_countOnes_30 + s1_offset);
  assign s1_outputPayload_cmd_data = s1_input_payload_cmd_data;
  assign s1_outputPayload_cmd_mask = s1_input_payload_cmd_mask;
  assign s1_outputPayload_index_0 = s1_inputIndexes_0;
  assign s1_outputPayload_index_1 = s1_inputIndexes_1;
  assign s1_outputPayload_index_2 = s1_inputIndexes_2;
  assign s1_outputPayload_index_3 = s1_inputIndexes_3;
  assign s1_outputPayload_index_4 = s1_inputIndexes_4;
  assign s1_outputPayload_index_5 = s1_inputIndexes_5;
  assign s1_outputPayload_index_6 = s1_inputIndexes_6;
  assign s1_outputPayload_index_7 = s1_inputIndexes_7;
  assign s1_outputPayload_index_8 = s1_inputIndexes_8;
  assign s1_outputPayload_index_9 = s1_inputIndexes_9;
  assign s1_outputPayload_index_10 = s1_inputIndexes_10;
  assign s1_outputPayload_index_11 = s1_inputIndexes_11;
  assign s1_outputPayload_index_12 = s1_inputIndexes_12;
  assign s1_outputPayload_index_13 = s1_inputIndexes_13;
  assign s1_outputPayload_index_14 = s1_inputIndexes_14;
  assign s1_outputPayload_index_15 = s1_inputIndexes_15;
  assign s1_outputPayload_index_16 = s1_inputIndexes_16;
  assign s1_outputPayload_index_17 = s1_inputIndexes_17;
  assign s1_outputPayload_index_18 = s1_inputIndexes_18;
  assign s1_outputPayload_index_19 = s1_inputIndexes_19;
  assign s1_outputPayload_index_20 = s1_inputIndexes_20;
  assign s1_outputPayload_index_21 = s1_inputIndexes_21;
  assign s1_outputPayload_index_22 = s1_inputIndexes_22;
  assign s1_outputPayload_index_23 = s1_inputIndexes_23;
  assign s1_outputPayload_index_24 = s1_inputIndexes_24;
  assign s1_outputPayload_index_25 = s1_inputIndexes_25;
  assign s1_outputPayload_index_26 = s1_inputIndexes_26;
  assign s1_outputPayload_index_27 = s1_inputIndexes_27;
  assign s1_outputPayload_index_28 = s1_inputIndexes_28;
  assign s1_outputPayload_index_29 = s1_inputIndexes_29;
  assign s1_outputPayload_index_30 = s1_inputIndexes_30;
  assign s1_outputPayload_index_31 = s1_inputIndexes_31;
  assign s1_outputPayload_last = s1_offsetNext[5];
  assign _zz_s1_outputPayload_selValid = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h0));
  assign _zz_s1_outputPayload_selValid_1 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h0));
  assign _zz_s1_outputPayload_selValid_2 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h0));
  assign _zz_s1_outputPayload_selValid_3 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h0));
  assign _zz_s1_outputPayload_selValid_4 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h0));
  assign _zz_s1_outputPayload_selValid_5 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h0));
  assign _zz_s1_outputPayload_selValid_6 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h0));
  assign _zz_s1_outputPayload_selValid_7 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h0));
  assign _zz_s1_outputPayload_selValid_8 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h0));
  assign _zz_s1_outputPayload_selValid_9 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h0));
  assign _zz_s1_outputPayload_selValid_10 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h0));
  assign _zz_s1_outputPayload_selValid_11 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h0));
  assign _zz_s1_outputPayload_selValid_12 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h0));
  assign _zz_s1_outputPayload_selValid_13 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h0));
  assign _zz_s1_outputPayload_selValid_14 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h0));
  assign _zz_s1_outputPayload_selValid_15 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h0));
  assign _zz_s1_outputPayload_selValid_16 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h0));
  assign _zz_s1_outputPayload_selValid_17 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h0));
  assign _zz_s1_outputPayload_selValid_18 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h0));
  assign _zz_s1_outputPayload_selValid_19 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h0));
  assign _zz_s1_outputPayload_selValid_20 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h0));
  assign _zz_s1_outputPayload_selValid_21 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h0));
  assign _zz_s1_outputPayload_selValid_22 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h0));
  assign _zz_s1_outputPayload_selValid_23 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h0));
  assign _zz_s1_outputPayload_selValid_24 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h0));
  assign _zz_s1_outputPayload_selValid_25 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h0));
  assign _zz_s1_outputPayload_selValid_26 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h0));
  assign _zz_s1_outputPayload_selValid_27 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h0));
  assign _zz_s1_outputPayload_selValid_28 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h0));
  assign _zz_s1_outputPayload_selValid_29 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h0));
  assign _zz_s1_outputPayload_selValid_30 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h0));
  assign _zz_s1_outputPayload_sel_0 = (((((((((((((((_zz_s1_outputPayload_selValid || _zz_s1_outputPayload_selValid_2) || _zz_s1_outputPayload_selValid_4) || _zz_s1_outputPayload_selValid_6) || _zz_s1_outputPayload_selValid_8) || _zz_s1_outputPayload_selValid_10) || _zz_s1_outputPayload_selValid_12) || _zz_s1_outputPayload_selValid_14) || _zz_s1_outputPayload_selValid_16) || _zz_s1_outputPayload_selValid_18) || _zz_s1_outputPayload_selValid_20) || _zz_s1_outputPayload_selValid_22) || _zz_s1_outputPayload_selValid_24) || _zz_s1_outputPayload_selValid_26) || _zz_s1_outputPayload_selValid_28) || _zz_s1_outputPayload_selValid_30);
  assign _zz_s1_outputPayload_sel_0_1 = (((((((((((((((_zz_s1_outputPayload_selValid_1 || _zz_s1_outputPayload_selValid_2) || _zz_s1_outputPayload_selValid_5) || _zz_s1_outputPayload_selValid_6) || _zz_s1_outputPayload_selValid_9) || _zz_s1_outputPayload_selValid_10) || _zz_s1_outputPayload_selValid_13) || _zz_s1_outputPayload_selValid_14) || _zz_s1_outputPayload_selValid_17) || _zz_s1_outputPayload_selValid_18) || _zz_s1_outputPayload_selValid_21) || _zz_s1_outputPayload_selValid_22) || _zz_s1_outputPayload_selValid_25) || _zz_s1_outputPayload_selValid_26) || _zz_s1_outputPayload_selValid_29) || _zz_s1_outputPayload_selValid_30);
  assign _zz_s1_outputPayload_sel_0_2 = (((((((((((((((_zz_s1_outputPayload_selValid_3 || _zz_s1_outputPayload_selValid_4) || _zz_s1_outputPayload_selValid_5) || _zz_s1_outputPayload_selValid_6) || _zz_s1_outputPayload_selValid_11) || _zz_s1_outputPayload_selValid_12) || _zz_s1_outputPayload_selValid_13) || _zz_s1_outputPayload_selValid_14) || _zz_s1_outputPayload_selValid_19) || _zz_s1_outputPayload_selValid_20) || _zz_s1_outputPayload_selValid_21) || _zz_s1_outputPayload_selValid_22) || _zz_s1_outputPayload_selValid_27) || _zz_s1_outputPayload_selValid_28) || _zz_s1_outputPayload_selValid_29) || _zz_s1_outputPayload_selValid_30);
  assign _zz_s1_outputPayload_sel_0_3 = (((((((((((((((_zz_s1_outputPayload_selValid_7 || _zz_s1_outputPayload_selValid_8) || _zz_s1_outputPayload_selValid_9) || _zz_s1_outputPayload_selValid_10) || _zz_s1_outputPayload_selValid_11) || _zz_s1_outputPayload_selValid_12) || _zz_s1_outputPayload_selValid_13) || _zz_s1_outputPayload_selValid_14) || _zz_s1_outputPayload_selValid_23) || _zz_s1_outputPayload_selValid_24) || _zz_s1_outputPayload_selValid_25) || _zz_s1_outputPayload_selValid_26) || _zz_s1_outputPayload_selValid_27) || _zz_s1_outputPayload_selValid_28) || _zz_s1_outputPayload_selValid_29) || _zz_s1_outputPayload_selValid_30);
  assign _zz_s1_outputPayload_sel_0_4 = (((((((((((((((_zz_s1_outputPayload_selValid_15 || _zz_s1_outputPayload_selValid_16) || _zz_s1_outputPayload_selValid_17) || _zz_s1_outputPayload_selValid_18) || _zz_s1_outputPayload_selValid_19) || _zz_s1_outputPayload_selValid_20) || _zz_s1_outputPayload_selValid_21) || _zz_s1_outputPayload_selValid_22) || _zz_s1_outputPayload_selValid_23) || _zz_s1_outputPayload_selValid_24) || _zz_s1_outputPayload_selValid_25) || _zz_s1_outputPayload_selValid_26) || _zz_s1_outputPayload_selValid_27) || _zz_s1_outputPayload_selValid_28) || _zz_s1_outputPayload_selValid_29) || _zz_s1_outputPayload_selValid_30);
  assign s1_outputPayload_sel_0 = {_zz_s1_outputPayload_sel_0_4,{_zz_s1_outputPayload_sel_0_3,{_zz_s1_outputPayload_sel_0_2,{_zz_s1_outputPayload_sel_0_1,_zz_s1_outputPayload_sel_0}}}};
  always @(*) begin
    s1_outputPayload_selValid[0] = ((|{_zz_s1_outputPayload_selValid_30,{_zz_s1_outputPayload_selValid_29,{_zz_s1_outputPayload_selValid_28,{_zz_s1_outputPayload_selValid_27,{_zz_s1_outputPayload_selValid_26,{_zz_s1_outputPayload_selValid_25,{_zz_s1_outputPayload_selValid_24,{_zz_s1_outputPayload_selValid_23,{_zz_s1_outputPayload_selValid_992,_zz_s1_outputPayload_selValid_993}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_0]);
    s1_outputPayload_selValid[1] = ((|{_zz_s1_outputPayload_selValid_61,{_zz_s1_outputPayload_selValid_60,{_zz_s1_outputPayload_selValid_59,{_zz_s1_outputPayload_selValid_58,{_zz_s1_outputPayload_selValid_57,{_zz_s1_outputPayload_selValid_56,{_zz_s1_outputPayload_selValid_55,{_zz_s1_outputPayload_selValid_54,{_zz_s1_outputPayload_selValid_998,_zz_s1_outputPayload_selValid_999}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_1]);
    s1_outputPayload_selValid[2] = ((|{_zz_s1_outputPayload_selValid_92,{_zz_s1_outputPayload_selValid_91,{_zz_s1_outputPayload_selValid_90,{_zz_s1_outputPayload_selValid_89,{_zz_s1_outputPayload_selValid_88,{_zz_s1_outputPayload_selValid_87,{_zz_s1_outputPayload_selValid_86,{_zz_s1_outputPayload_selValid_85,{_zz_s1_outputPayload_selValid_1004,_zz_s1_outputPayload_selValid_1005}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_2]);
    s1_outputPayload_selValid[3] = ((|{_zz_s1_outputPayload_selValid_123,{_zz_s1_outputPayload_selValid_122,{_zz_s1_outputPayload_selValid_121,{_zz_s1_outputPayload_selValid_120,{_zz_s1_outputPayload_selValid_119,{_zz_s1_outputPayload_selValid_118,{_zz_s1_outputPayload_selValid_117,{_zz_s1_outputPayload_selValid_116,{_zz_s1_outputPayload_selValid_1010,_zz_s1_outputPayload_selValid_1011}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_3]);
    s1_outputPayload_selValid[4] = ((|{_zz_s1_outputPayload_selValid_154,{_zz_s1_outputPayload_selValid_153,{_zz_s1_outputPayload_selValid_152,{_zz_s1_outputPayload_selValid_151,{_zz_s1_outputPayload_selValid_150,{_zz_s1_outputPayload_selValid_149,{_zz_s1_outputPayload_selValid_148,{_zz_s1_outputPayload_selValid_147,{_zz_s1_outputPayload_selValid_1016,_zz_s1_outputPayload_selValid_1017}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_4]);
    s1_outputPayload_selValid[5] = ((|{_zz_s1_outputPayload_selValid_185,{_zz_s1_outputPayload_selValid_184,{_zz_s1_outputPayload_selValid_183,{_zz_s1_outputPayload_selValid_182,{_zz_s1_outputPayload_selValid_181,{_zz_s1_outputPayload_selValid_180,{_zz_s1_outputPayload_selValid_179,{_zz_s1_outputPayload_selValid_178,{_zz_s1_outputPayload_selValid_1022,_zz_s1_outputPayload_selValid_1023}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_5]);
    s1_outputPayload_selValid[6] = ((|{_zz_s1_outputPayload_selValid_216,{_zz_s1_outputPayload_selValid_215,{_zz_s1_outputPayload_selValid_214,{_zz_s1_outputPayload_selValid_213,{_zz_s1_outputPayload_selValid_212,{_zz_s1_outputPayload_selValid_211,{_zz_s1_outputPayload_selValid_210,{_zz_s1_outputPayload_selValid_209,{_zz_s1_outputPayload_selValid_1028,_zz_s1_outputPayload_selValid_1029}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_6]);
    s1_outputPayload_selValid[7] = ((|{_zz_s1_outputPayload_selValid_247,{_zz_s1_outputPayload_selValid_246,{_zz_s1_outputPayload_selValid_245,{_zz_s1_outputPayload_selValid_244,{_zz_s1_outputPayload_selValid_243,{_zz_s1_outputPayload_selValid_242,{_zz_s1_outputPayload_selValid_241,{_zz_s1_outputPayload_selValid_240,{_zz_s1_outputPayload_selValid_1034,_zz_s1_outputPayload_selValid_1035}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_7]);
    s1_outputPayload_selValid[8] = ((|{_zz_s1_outputPayload_selValid_278,{_zz_s1_outputPayload_selValid_277,{_zz_s1_outputPayload_selValid_276,{_zz_s1_outputPayload_selValid_275,{_zz_s1_outputPayload_selValid_274,{_zz_s1_outputPayload_selValid_273,{_zz_s1_outputPayload_selValid_272,{_zz_s1_outputPayload_selValid_271,{_zz_s1_outputPayload_selValid_1040,_zz_s1_outputPayload_selValid_1041}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_8]);
    s1_outputPayload_selValid[9] = ((|{_zz_s1_outputPayload_selValid_309,{_zz_s1_outputPayload_selValid_308,{_zz_s1_outputPayload_selValid_307,{_zz_s1_outputPayload_selValid_306,{_zz_s1_outputPayload_selValid_305,{_zz_s1_outputPayload_selValid_304,{_zz_s1_outputPayload_selValid_303,{_zz_s1_outputPayload_selValid_302,{_zz_s1_outputPayload_selValid_1046,_zz_s1_outputPayload_selValid_1047}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_9]);
    s1_outputPayload_selValid[10] = ((|{_zz_s1_outputPayload_selValid_340,{_zz_s1_outputPayload_selValid_339,{_zz_s1_outputPayload_selValid_338,{_zz_s1_outputPayload_selValid_337,{_zz_s1_outputPayload_selValid_336,{_zz_s1_outputPayload_selValid_335,{_zz_s1_outputPayload_selValid_334,{_zz_s1_outputPayload_selValid_333,{_zz_s1_outputPayload_selValid_1052,_zz_s1_outputPayload_selValid_1053}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_10]);
    s1_outputPayload_selValid[11] = ((|{_zz_s1_outputPayload_selValid_371,{_zz_s1_outputPayload_selValid_370,{_zz_s1_outputPayload_selValid_369,{_zz_s1_outputPayload_selValid_368,{_zz_s1_outputPayload_selValid_367,{_zz_s1_outputPayload_selValid_366,{_zz_s1_outputPayload_selValid_365,{_zz_s1_outputPayload_selValid_364,{_zz_s1_outputPayload_selValid_1058,_zz_s1_outputPayload_selValid_1059}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_11]);
    s1_outputPayload_selValid[12] = ((|{_zz_s1_outputPayload_selValid_402,{_zz_s1_outputPayload_selValid_401,{_zz_s1_outputPayload_selValid_400,{_zz_s1_outputPayload_selValid_399,{_zz_s1_outputPayload_selValid_398,{_zz_s1_outputPayload_selValid_397,{_zz_s1_outputPayload_selValid_396,{_zz_s1_outputPayload_selValid_395,{_zz_s1_outputPayload_selValid_1064,_zz_s1_outputPayload_selValid_1065}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_12]);
    s1_outputPayload_selValid[13] = ((|{_zz_s1_outputPayload_selValid_433,{_zz_s1_outputPayload_selValid_432,{_zz_s1_outputPayload_selValid_431,{_zz_s1_outputPayload_selValid_430,{_zz_s1_outputPayload_selValid_429,{_zz_s1_outputPayload_selValid_428,{_zz_s1_outputPayload_selValid_427,{_zz_s1_outputPayload_selValid_426,{_zz_s1_outputPayload_selValid_1070,_zz_s1_outputPayload_selValid_1071}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_13]);
    s1_outputPayload_selValid[14] = ((|{_zz_s1_outputPayload_selValid_464,{_zz_s1_outputPayload_selValid_463,{_zz_s1_outputPayload_selValid_462,{_zz_s1_outputPayload_selValid_461,{_zz_s1_outputPayload_selValid_460,{_zz_s1_outputPayload_selValid_459,{_zz_s1_outputPayload_selValid_458,{_zz_s1_outputPayload_selValid_457,{_zz_s1_outputPayload_selValid_1076,_zz_s1_outputPayload_selValid_1077}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_14]);
    s1_outputPayload_selValid[15] = ((|{_zz_s1_outputPayload_selValid_495,{_zz_s1_outputPayload_selValid_494,{_zz_s1_outputPayload_selValid_493,{_zz_s1_outputPayload_selValid_492,{_zz_s1_outputPayload_selValid_491,{_zz_s1_outputPayload_selValid_490,{_zz_s1_outputPayload_selValid_489,{_zz_s1_outputPayload_selValid_488,{_zz_s1_outputPayload_selValid_1082,_zz_s1_outputPayload_selValid_1083}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_15]);
    s1_outputPayload_selValid[16] = ((|{_zz_s1_outputPayload_selValid_526,{_zz_s1_outputPayload_selValid_525,{_zz_s1_outputPayload_selValid_524,{_zz_s1_outputPayload_selValid_523,{_zz_s1_outputPayload_selValid_522,{_zz_s1_outputPayload_selValid_521,{_zz_s1_outputPayload_selValid_520,{_zz_s1_outputPayload_selValid_519,{_zz_s1_outputPayload_selValid_1088,_zz_s1_outputPayload_selValid_1089}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_16]);
    s1_outputPayload_selValid[17] = ((|{_zz_s1_outputPayload_selValid_557,{_zz_s1_outputPayload_selValid_556,{_zz_s1_outputPayload_selValid_555,{_zz_s1_outputPayload_selValid_554,{_zz_s1_outputPayload_selValid_553,{_zz_s1_outputPayload_selValid_552,{_zz_s1_outputPayload_selValid_551,{_zz_s1_outputPayload_selValid_550,{_zz_s1_outputPayload_selValid_1094,_zz_s1_outputPayload_selValid_1095}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_17]);
    s1_outputPayload_selValid[18] = ((|{_zz_s1_outputPayload_selValid_588,{_zz_s1_outputPayload_selValid_587,{_zz_s1_outputPayload_selValid_586,{_zz_s1_outputPayload_selValid_585,{_zz_s1_outputPayload_selValid_584,{_zz_s1_outputPayload_selValid_583,{_zz_s1_outputPayload_selValid_582,{_zz_s1_outputPayload_selValid_581,{_zz_s1_outputPayload_selValid_1100,_zz_s1_outputPayload_selValid_1101}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_18]);
    s1_outputPayload_selValid[19] = ((|{_zz_s1_outputPayload_selValid_619,{_zz_s1_outputPayload_selValid_618,{_zz_s1_outputPayload_selValid_617,{_zz_s1_outputPayload_selValid_616,{_zz_s1_outputPayload_selValid_615,{_zz_s1_outputPayload_selValid_614,{_zz_s1_outputPayload_selValid_613,{_zz_s1_outputPayload_selValid_612,{_zz_s1_outputPayload_selValid_1106,_zz_s1_outputPayload_selValid_1107}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_19]);
    s1_outputPayload_selValid[20] = ((|{_zz_s1_outputPayload_selValid_650,{_zz_s1_outputPayload_selValid_649,{_zz_s1_outputPayload_selValid_648,{_zz_s1_outputPayload_selValid_647,{_zz_s1_outputPayload_selValid_646,{_zz_s1_outputPayload_selValid_645,{_zz_s1_outputPayload_selValid_644,{_zz_s1_outputPayload_selValid_643,{_zz_s1_outputPayload_selValid_1112,_zz_s1_outputPayload_selValid_1113}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_20]);
    s1_outputPayload_selValid[21] = ((|{_zz_s1_outputPayload_selValid_681,{_zz_s1_outputPayload_selValid_680,{_zz_s1_outputPayload_selValid_679,{_zz_s1_outputPayload_selValid_678,{_zz_s1_outputPayload_selValid_677,{_zz_s1_outputPayload_selValid_676,{_zz_s1_outputPayload_selValid_675,{_zz_s1_outputPayload_selValid_674,{_zz_s1_outputPayload_selValid_1118,_zz_s1_outputPayload_selValid_1119}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_21]);
    s1_outputPayload_selValid[22] = ((|{_zz_s1_outputPayload_selValid_712,{_zz_s1_outputPayload_selValid_711,{_zz_s1_outputPayload_selValid_710,{_zz_s1_outputPayload_selValid_709,{_zz_s1_outputPayload_selValid_708,{_zz_s1_outputPayload_selValid_707,{_zz_s1_outputPayload_selValid_706,{_zz_s1_outputPayload_selValid_705,{_zz_s1_outputPayload_selValid_1124,_zz_s1_outputPayload_selValid_1125}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_22]);
    s1_outputPayload_selValid[23] = ((|{_zz_s1_outputPayload_selValid_743,{_zz_s1_outputPayload_selValid_742,{_zz_s1_outputPayload_selValid_741,{_zz_s1_outputPayload_selValid_740,{_zz_s1_outputPayload_selValid_739,{_zz_s1_outputPayload_selValid_738,{_zz_s1_outputPayload_selValid_737,{_zz_s1_outputPayload_selValid_736,{_zz_s1_outputPayload_selValid_1130,_zz_s1_outputPayload_selValid_1131}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_23]);
    s1_outputPayload_selValid[24] = ((|{_zz_s1_outputPayload_selValid_774,{_zz_s1_outputPayload_selValid_773,{_zz_s1_outputPayload_selValid_772,{_zz_s1_outputPayload_selValid_771,{_zz_s1_outputPayload_selValid_770,{_zz_s1_outputPayload_selValid_769,{_zz_s1_outputPayload_selValid_768,{_zz_s1_outputPayload_selValid_767,{_zz_s1_outputPayload_selValid_1136,_zz_s1_outputPayload_selValid_1137}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_24]);
    s1_outputPayload_selValid[25] = ((|{_zz_s1_outputPayload_selValid_805,{_zz_s1_outputPayload_selValid_804,{_zz_s1_outputPayload_selValid_803,{_zz_s1_outputPayload_selValid_802,{_zz_s1_outputPayload_selValid_801,{_zz_s1_outputPayload_selValid_800,{_zz_s1_outputPayload_selValid_799,{_zz_s1_outputPayload_selValid_798,{_zz_s1_outputPayload_selValid_1142,_zz_s1_outputPayload_selValid_1143}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_25]);
    s1_outputPayload_selValid[26] = ((|{_zz_s1_outputPayload_selValid_836,{_zz_s1_outputPayload_selValid_835,{_zz_s1_outputPayload_selValid_834,{_zz_s1_outputPayload_selValid_833,{_zz_s1_outputPayload_selValid_832,{_zz_s1_outputPayload_selValid_831,{_zz_s1_outputPayload_selValid_830,{_zz_s1_outputPayload_selValid_829,{_zz_s1_outputPayload_selValid_1148,_zz_s1_outputPayload_selValid_1149}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_26]);
    s1_outputPayload_selValid[27] = ((|{_zz_s1_outputPayload_selValid_867,{_zz_s1_outputPayload_selValid_866,{_zz_s1_outputPayload_selValid_865,{_zz_s1_outputPayload_selValid_864,{_zz_s1_outputPayload_selValid_863,{_zz_s1_outputPayload_selValid_862,{_zz_s1_outputPayload_selValid_861,{_zz_s1_outputPayload_selValid_860,{_zz_s1_outputPayload_selValid_1154,_zz_s1_outputPayload_selValid_1155}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_27]);
    s1_outputPayload_selValid[28] = ((|{_zz_s1_outputPayload_selValid_898,{_zz_s1_outputPayload_selValid_897,{_zz_s1_outputPayload_selValid_896,{_zz_s1_outputPayload_selValid_895,{_zz_s1_outputPayload_selValid_894,{_zz_s1_outputPayload_selValid_893,{_zz_s1_outputPayload_selValid_892,{_zz_s1_outputPayload_selValid_891,{_zz_s1_outputPayload_selValid_1160,_zz_s1_outputPayload_selValid_1161}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_28]);
    s1_outputPayload_selValid[29] = ((|{_zz_s1_outputPayload_selValid_929,{_zz_s1_outputPayload_selValid_928,{_zz_s1_outputPayload_selValid_927,{_zz_s1_outputPayload_selValid_926,{_zz_s1_outputPayload_selValid_925,{_zz_s1_outputPayload_selValid_924,{_zz_s1_outputPayload_selValid_923,{_zz_s1_outputPayload_selValid_922,{_zz_s1_outputPayload_selValid_1166,_zz_s1_outputPayload_selValid_1167}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_29]);
    s1_outputPayload_selValid[30] = ((|{_zz_s1_outputPayload_selValid_960,{_zz_s1_outputPayload_selValid_959,{_zz_s1_outputPayload_selValid_958,{_zz_s1_outputPayload_selValid_957,{_zz_s1_outputPayload_selValid_956,{_zz_s1_outputPayload_selValid_955,{_zz_s1_outputPayload_selValid_954,{_zz_s1_outputPayload_selValid_953,{_zz_s1_outputPayload_selValid_1172,_zz_s1_outputPayload_selValid_1173}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_30]);
    s1_outputPayload_selValid[31] = ((|{_zz_s1_outputPayload_selValid_991,{_zz_s1_outputPayload_selValid_990,{_zz_s1_outputPayload_selValid_989,{_zz_s1_outputPayload_selValid_988,{_zz_s1_outputPayload_selValid_987,{_zz_s1_outputPayload_selValid_986,{_zz_s1_outputPayload_selValid_985,{_zz_s1_outputPayload_selValid_984,{_zz_s1_outputPayload_selValid_1178,_zz_s1_outputPayload_selValid_1179}}}}}}}}}) && s1_outputPayload_cmd_mask[s1_outputPayload_sel_31]);
  end

  assign _zz_s1_outputPayload_selValid_31 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h01));
  assign _zz_s1_outputPayload_selValid_32 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h01));
  assign _zz_s1_outputPayload_selValid_33 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h01));
  assign _zz_s1_outputPayload_selValid_34 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h01));
  assign _zz_s1_outputPayload_selValid_35 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h01));
  assign _zz_s1_outputPayload_selValid_36 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h01));
  assign _zz_s1_outputPayload_selValid_37 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h01));
  assign _zz_s1_outputPayload_selValid_38 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h01));
  assign _zz_s1_outputPayload_selValid_39 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h01));
  assign _zz_s1_outputPayload_selValid_40 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h01));
  assign _zz_s1_outputPayload_selValid_41 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h01));
  assign _zz_s1_outputPayload_selValid_42 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h01));
  assign _zz_s1_outputPayload_selValid_43 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h01));
  assign _zz_s1_outputPayload_selValid_44 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h01));
  assign _zz_s1_outputPayload_selValid_45 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h01));
  assign _zz_s1_outputPayload_selValid_46 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h01));
  assign _zz_s1_outputPayload_selValid_47 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h01));
  assign _zz_s1_outputPayload_selValid_48 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h01));
  assign _zz_s1_outputPayload_selValid_49 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h01));
  assign _zz_s1_outputPayload_selValid_50 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h01));
  assign _zz_s1_outputPayload_selValid_51 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h01));
  assign _zz_s1_outputPayload_selValid_52 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h01));
  assign _zz_s1_outputPayload_selValid_53 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h01));
  assign _zz_s1_outputPayload_selValid_54 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h01));
  assign _zz_s1_outputPayload_selValid_55 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h01));
  assign _zz_s1_outputPayload_selValid_56 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h01));
  assign _zz_s1_outputPayload_selValid_57 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h01));
  assign _zz_s1_outputPayload_selValid_58 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h01));
  assign _zz_s1_outputPayload_selValid_59 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h01));
  assign _zz_s1_outputPayload_selValid_60 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h01));
  assign _zz_s1_outputPayload_selValid_61 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h01));
  assign _zz_s1_outputPayload_sel_1 = (((((((((((((((_zz_s1_outputPayload_selValid_31 || _zz_s1_outputPayload_selValid_33) || _zz_s1_outputPayload_selValid_35) || _zz_s1_outputPayload_selValid_37) || _zz_s1_outputPayload_selValid_39) || _zz_s1_outputPayload_selValid_41) || _zz_s1_outputPayload_selValid_43) || _zz_s1_outputPayload_selValid_45) || _zz_s1_outputPayload_selValid_47) || _zz_s1_outputPayload_selValid_49) || _zz_s1_outputPayload_selValid_51) || _zz_s1_outputPayload_selValid_53) || _zz_s1_outputPayload_selValid_55) || _zz_s1_outputPayload_selValid_57) || _zz_s1_outputPayload_selValid_59) || _zz_s1_outputPayload_selValid_61);
  assign _zz_s1_outputPayload_sel_1_1 = (((((((((((((((_zz_s1_outputPayload_selValid_32 || _zz_s1_outputPayload_selValid_33) || _zz_s1_outputPayload_selValid_36) || _zz_s1_outputPayload_selValid_37) || _zz_s1_outputPayload_selValid_40) || _zz_s1_outputPayload_selValid_41) || _zz_s1_outputPayload_selValid_44) || _zz_s1_outputPayload_selValid_45) || _zz_s1_outputPayload_selValid_48) || _zz_s1_outputPayload_selValid_49) || _zz_s1_outputPayload_selValid_52) || _zz_s1_outputPayload_selValid_53) || _zz_s1_outputPayload_selValid_56) || _zz_s1_outputPayload_selValid_57) || _zz_s1_outputPayload_selValid_60) || _zz_s1_outputPayload_selValid_61);
  assign _zz_s1_outputPayload_sel_1_2 = (((((((((((((((_zz_s1_outputPayload_selValid_34 || _zz_s1_outputPayload_selValid_35) || _zz_s1_outputPayload_selValid_36) || _zz_s1_outputPayload_selValid_37) || _zz_s1_outputPayload_selValid_42) || _zz_s1_outputPayload_selValid_43) || _zz_s1_outputPayload_selValid_44) || _zz_s1_outputPayload_selValid_45) || _zz_s1_outputPayload_selValid_50) || _zz_s1_outputPayload_selValid_51) || _zz_s1_outputPayload_selValid_52) || _zz_s1_outputPayload_selValid_53) || _zz_s1_outputPayload_selValid_58) || _zz_s1_outputPayload_selValid_59) || _zz_s1_outputPayload_selValid_60) || _zz_s1_outputPayload_selValid_61);
  assign _zz_s1_outputPayload_sel_1_3 = (((((((((((((((_zz_s1_outputPayload_selValid_38 || _zz_s1_outputPayload_selValid_39) || _zz_s1_outputPayload_selValid_40) || _zz_s1_outputPayload_selValid_41) || _zz_s1_outputPayload_selValid_42) || _zz_s1_outputPayload_selValid_43) || _zz_s1_outputPayload_selValid_44) || _zz_s1_outputPayload_selValid_45) || _zz_s1_outputPayload_selValid_54) || _zz_s1_outputPayload_selValid_55) || _zz_s1_outputPayload_selValid_56) || _zz_s1_outputPayload_selValid_57) || _zz_s1_outputPayload_selValid_58) || _zz_s1_outputPayload_selValid_59) || _zz_s1_outputPayload_selValid_60) || _zz_s1_outputPayload_selValid_61);
  assign _zz_s1_outputPayload_sel_1_4 = (((((((((((((((_zz_s1_outputPayload_selValid_46 || _zz_s1_outputPayload_selValid_47) || _zz_s1_outputPayload_selValid_48) || _zz_s1_outputPayload_selValid_49) || _zz_s1_outputPayload_selValid_50) || _zz_s1_outputPayload_selValid_51) || _zz_s1_outputPayload_selValid_52) || _zz_s1_outputPayload_selValid_53) || _zz_s1_outputPayload_selValid_54) || _zz_s1_outputPayload_selValid_55) || _zz_s1_outputPayload_selValid_56) || _zz_s1_outputPayload_selValid_57) || _zz_s1_outputPayload_selValid_58) || _zz_s1_outputPayload_selValid_59) || _zz_s1_outputPayload_selValid_60) || _zz_s1_outputPayload_selValid_61);
  assign s1_outputPayload_sel_1 = {_zz_s1_outputPayload_sel_1_4,{_zz_s1_outputPayload_sel_1_3,{_zz_s1_outputPayload_sel_1_2,{_zz_s1_outputPayload_sel_1_1,_zz_s1_outputPayload_sel_1}}}};
  assign _zz_s1_outputPayload_selValid_62 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h02));
  assign _zz_s1_outputPayload_selValid_63 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h02));
  assign _zz_s1_outputPayload_selValid_64 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h02));
  assign _zz_s1_outputPayload_selValid_65 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h02));
  assign _zz_s1_outputPayload_selValid_66 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h02));
  assign _zz_s1_outputPayload_selValid_67 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h02));
  assign _zz_s1_outputPayload_selValid_68 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h02));
  assign _zz_s1_outputPayload_selValid_69 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h02));
  assign _zz_s1_outputPayload_selValid_70 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h02));
  assign _zz_s1_outputPayload_selValid_71 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h02));
  assign _zz_s1_outputPayload_selValid_72 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h02));
  assign _zz_s1_outputPayload_selValid_73 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h02));
  assign _zz_s1_outputPayload_selValid_74 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h02));
  assign _zz_s1_outputPayload_selValid_75 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h02));
  assign _zz_s1_outputPayload_selValid_76 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h02));
  assign _zz_s1_outputPayload_selValid_77 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h02));
  assign _zz_s1_outputPayload_selValid_78 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h02));
  assign _zz_s1_outputPayload_selValid_79 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h02));
  assign _zz_s1_outputPayload_selValid_80 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h02));
  assign _zz_s1_outputPayload_selValid_81 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h02));
  assign _zz_s1_outputPayload_selValid_82 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h02));
  assign _zz_s1_outputPayload_selValid_83 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h02));
  assign _zz_s1_outputPayload_selValid_84 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h02));
  assign _zz_s1_outputPayload_selValid_85 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h02));
  assign _zz_s1_outputPayload_selValid_86 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h02));
  assign _zz_s1_outputPayload_selValid_87 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h02));
  assign _zz_s1_outputPayload_selValid_88 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h02));
  assign _zz_s1_outputPayload_selValid_89 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h02));
  assign _zz_s1_outputPayload_selValid_90 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h02));
  assign _zz_s1_outputPayload_selValid_91 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h02));
  assign _zz_s1_outputPayload_selValid_92 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h02));
  assign _zz_s1_outputPayload_sel_2 = (((((((((((((((_zz_s1_outputPayload_selValid_62 || _zz_s1_outputPayload_selValid_64) || _zz_s1_outputPayload_selValid_66) || _zz_s1_outputPayload_selValid_68) || _zz_s1_outputPayload_selValid_70) || _zz_s1_outputPayload_selValid_72) || _zz_s1_outputPayload_selValid_74) || _zz_s1_outputPayload_selValid_76) || _zz_s1_outputPayload_selValid_78) || _zz_s1_outputPayload_selValid_80) || _zz_s1_outputPayload_selValid_82) || _zz_s1_outputPayload_selValid_84) || _zz_s1_outputPayload_selValid_86) || _zz_s1_outputPayload_selValid_88) || _zz_s1_outputPayload_selValid_90) || _zz_s1_outputPayload_selValid_92);
  assign _zz_s1_outputPayload_sel_2_1 = (((((((((((((((_zz_s1_outputPayload_selValid_63 || _zz_s1_outputPayload_selValid_64) || _zz_s1_outputPayload_selValid_67) || _zz_s1_outputPayload_selValid_68) || _zz_s1_outputPayload_selValid_71) || _zz_s1_outputPayload_selValid_72) || _zz_s1_outputPayload_selValid_75) || _zz_s1_outputPayload_selValid_76) || _zz_s1_outputPayload_selValid_79) || _zz_s1_outputPayload_selValid_80) || _zz_s1_outputPayload_selValid_83) || _zz_s1_outputPayload_selValid_84) || _zz_s1_outputPayload_selValid_87) || _zz_s1_outputPayload_selValid_88) || _zz_s1_outputPayload_selValid_91) || _zz_s1_outputPayload_selValid_92);
  assign _zz_s1_outputPayload_sel_2_2 = (((((((((((((((_zz_s1_outputPayload_selValid_65 || _zz_s1_outputPayload_selValid_66) || _zz_s1_outputPayload_selValid_67) || _zz_s1_outputPayload_selValid_68) || _zz_s1_outputPayload_selValid_73) || _zz_s1_outputPayload_selValid_74) || _zz_s1_outputPayload_selValid_75) || _zz_s1_outputPayload_selValid_76) || _zz_s1_outputPayload_selValid_81) || _zz_s1_outputPayload_selValid_82) || _zz_s1_outputPayload_selValid_83) || _zz_s1_outputPayload_selValid_84) || _zz_s1_outputPayload_selValid_89) || _zz_s1_outputPayload_selValid_90) || _zz_s1_outputPayload_selValid_91) || _zz_s1_outputPayload_selValid_92);
  assign _zz_s1_outputPayload_sel_2_3 = (((((((((((((((_zz_s1_outputPayload_selValid_69 || _zz_s1_outputPayload_selValid_70) || _zz_s1_outputPayload_selValid_71) || _zz_s1_outputPayload_selValid_72) || _zz_s1_outputPayload_selValid_73) || _zz_s1_outputPayload_selValid_74) || _zz_s1_outputPayload_selValid_75) || _zz_s1_outputPayload_selValid_76) || _zz_s1_outputPayload_selValid_85) || _zz_s1_outputPayload_selValid_86) || _zz_s1_outputPayload_selValid_87) || _zz_s1_outputPayload_selValid_88) || _zz_s1_outputPayload_selValid_89) || _zz_s1_outputPayload_selValid_90) || _zz_s1_outputPayload_selValid_91) || _zz_s1_outputPayload_selValid_92);
  assign _zz_s1_outputPayload_sel_2_4 = (((((((((((((((_zz_s1_outputPayload_selValid_77 || _zz_s1_outputPayload_selValid_78) || _zz_s1_outputPayload_selValid_79) || _zz_s1_outputPayload_selValid_80) || _zz_s1_outputPayload_selValid_81) || _zz_s1_outputPayload_selValid_82) || _zz_s1_outputPayload_selValid_83) || _zz_s1_outputPayload_selValid_84) || _zz_s1_outputPayload_selValid_85) || _zz_s1_outputPayload_selValid_86) || _zz_s1_outputPayload_selValid_87) || _zz_s1_outputPayload_selValid_88) || _zz_s1_outputPayload_selValid_89) || _zz_s1_outputPayload_selValid_90) || _zz_s1_outputPayload_selValid_91) || _zz_s1_outputPayload_selValid_92);
  assign s1_outputPayload_sel_2 = {_zz_s1_outputPayload_sel_2_4,{_zz_s1_outputPayload_sel_2_3,{_zz_s1_outputPayload_sel_2_2,{_zz_s1_outputPayload_sel_2_1,_zz_s1_outputPayload_sel_2}}}};
  assign _zz_s1_outputPayload_selValid_93 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h03));
  assign _zz_s1_outputPayload_selValid_94 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h03));
  assign _zz_s1_outputPayload_selValid_95 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h03));
  assign _zz_s1_outputPayload_selValid_96 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h03));
  assign _zz_s1_outputPayload_selValid_97 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h03));
  assign _zz_s1_outputPayload_selValid_98 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h03));
  assign _zz_s1_outputPayload_selValid_99 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h03));
  assign _zz_s1_outputPayload_selValid_100 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h03));
  assign _zz_s1_outputPayload_selValid_101 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h03));
  assign _zz_s1_outputPayload_selValid_102 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h03));
  assign _zz_s1_outputPayload_selValid_103 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h03));
  assign _zz_s1_outputPayload_selValid_104 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h03));
  assign _zz_s1_outputPayload_selValid_105 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h03));
  assign _zz_s1_outputPayload_selValid_106 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h03));
  assign _zz_s1_outputPayload_selValid_107 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h03));
  assign _zz_s1_outputPayload_selValid_108 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h03));
  assign _zz_s1_outputPayload_selValid_109 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h03));
  assign _zz_s1_outputPayload_selValid_110 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h03));
  assign _zz_s1_outputPayload_selValid_111 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h03));
  assign _zz_s1_outputPayload_selValid_112 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h03));
  assign _zz_s1_outputPayload_selValid_113 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h03));
  assign _zz_s1_outputPayload_selValid_114 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h03));
  assign _zz_s1_outputPayload_selValid_115 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h03));
  assign _zz_s1_outputPayload_selValid_116 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h03));
  assign _zz_s1_outputPayload_selValid_117 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h03));
  assign _zz_s1_outputPayload_selValid_118 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h03));
  assign _zz_s1_outputPayload_selValid_119 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h03));
  assign _zz_s1_outputPayload_selValid_120 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h03));
  assign _zz_s1_outputPayload_selValid_121 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h03));
  assign _zz_s1_outputPayload_selValid_122 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h03));
  assign _zz_s1_outputPayload_selValid_123 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h03));
  assign _zz_s1_outputPayload_sel_3 = (((((((((((((((_zz_s1_outputPayload_selValid_93 || _zz_s1_outputPayload_selValid_95) || _zz_s1_outputPayload_selValid_97) || _zz_s1_outputPayload_selValid_99) || _zz_s1_outputPayload_selValid_101) || _zz_s1_outputPayload_selValid_103) || _zz_s1_outputPayload_selValid_105) || _zz_s1_outputPayload_selValid_107) || _zz_s1_outputPayload_selValid_109) || _zz_s1_outputPayload_selValid_111) || _zz_s1_outputPayload_selValid_113) || _zz_s1_outputPayload_selValid_115) || _zz_s1_outputPayload_selValid_117) || _zz_s1_outputPayload_selValid_119) || _zz_s1_outputPayload_selValid_121) || _zz_s1_outputPayload_selValid_123);
  assign _zz_s1_outputPayload_sel_3_1 = (((((((((((((((_zz_s1_outputPayload_selValid_94 || _zz_s1_outputPayload_selValid_95) || _zz_s1_outputPayload_selValid_98) || _zz_s1_outputPayload_selValid_99) || _zz_s1_outputPayload_selValid_102) || _zz_s1_outputPayload_selValid_103) || _zz_s1_outputPayload_selValid_106) || _zz_s1_outputPayload_selValid_107) || _zz_s1_outputPayload_selValid_110) || _zz_s1_outputPayload_selValid_111) || _zz_s1_outputPayload_selValid_114) || _zz_s1_outputPayload_selValid_115) || _zz_s1_outputPayload_selValid_118) || _zz_s1_outputPayload_selValid_119) || _zz_s1_outputPayload_selValid_122) || _zz_s1_outputPayload_selValid_123);
  assign _zz_s1_outputPayload_sel_3_2 = (((((((((((((((_zz_s1_outputPayload_selValid_96 || _zz_s1_outputPayload_selValid_97) || _zz_s1_outputPayload_selValid_98) || _zz_s1_outputPayload_selValid_99) || _zz_s1_outputPayload_selValid_104) || _zz_s1_outputPayload_selValid_105) || _zz_s1_outputPayload_selValid_106) || _zz_s1_outputPayload_selValid_107) || _zz_s1_outputPayload_selValid_112) || _zz_s1_outputPayload_selValid_113) || _zz_s1_outputPayload_selValid_114) || _zz_s1_outputPayload_selValid_115) || _zz_s1_outputPayload_selValid_120) || _zz_s1_outputPayload_selValid_121) || _zz_s1_outputPayload_selValid_122) || _zz_s1_outputPayload_selValid_123);
  assign _zz_s1_outputPayload_sel_3_3 = (((((((((((((((_zz_s1_outputPayload_selValid_100 || _zz_s1_outputPayload_selValid_101) || _zz_s1_outputPayload_selValid_102) || _zz_s1_outputPayload_selValid_103) || _zz_s1_outputPayload_selValid_104) || _zz_s1_outputPayload_selValid_105) || _zz_s1_outputPayload_selValid_106) || _zz_s1_outputPayload_selValid_107) || _zz_s1_outputPayload_selValid_116) || _zz_s1_outputPayload_selValid_117) || _zz_s1_outputPayload_selValid_118) || _zz_s1_outputPayload_selValid_119) || _zz_s1_outputPayload_selValid_120) || _zz_s1_outputPayload_selValid_121) || _zz_s1_outputPayload_selValid_122) || _zz_s1_outputPayload_selValid_123);
  assign _zz_s1_outputPayload_sel_3_4 = (((((((((((((((_zz_s1_outputPayload_selValid_108 || _zz_s1_outputPayload_selValid_109) || _zz_s1_outputPayload_selValid_110) || _zz_s1_outputPayload_selValid_111) || _zz_s1_outputPayload_selValid_112) || _zz_s1_outputPayload_selValid_113) || _zz_s1_outputPayload_selValid_114) || _zz_s1_outputPayload_selValid_115) || _zz_s1_outputPayload_selValid_116) || _zz_s1_outputPayload_selValid_117) || _zz_s1_outputPayload_selValid_118) || _zz_s1_outputPayload_selValid_119) || _zz_s1_outputPayload_selValid_120) || _zz_s1_outputPayload_selValid_121) || _zz_s1_outputPayload_selValid_122) || _zz_s1_outputPayload_selValid_123);
  assign s1_outputPayload_sel_3 = {_zz_s1_outputPayload_sel_3_4,{_zz_s1_outputPayload_sel_3_3,{_zz_s1_outputPayload_sel_3_2,{_zz_s1_outputPayload_sel_3_1,_zz_s1_outputPayload_sel_3}}}};
  assign _zz_s1_outputPayload_selValid_124 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h04));
  assign _zz_s1_outputPayload_selValid_125 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h04));
  assign _zz_s1_outputPayload_selValid_126 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h04));
  assign _zz_s1_outputPayload_selValid_127 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h04));
  assign _zz_s1_outputPayload_selValid_128 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h04));
  assign _zz_s1_outputPayload_selValid_129 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h04));
  assign _zz_s1_outputPayload_selValid_130 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h04));
  assign _zz_s1_outputPayload_selValid_131 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h04));
  assign _zz_s1_outputPayload_selValid_132 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h04));
  assign _zz_s1_outputPayload_selValid_133 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h04));
  assign _zz_s1_outputPayload_selValid_134 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h04));
  assign _zz_s1_outputPayload_selValid_135 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h04));
  assign _zz_s1_outputPayload_selValid_136 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h04));
  assign _zz_s1_outputPayload_selValid_137 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h04));
  assign _zz_s1_outputPayload_selValid_138 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h04));
  assign _zz_s1_outputPayload_selValid_139 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h04));
  assign _zz_s1_outputPayload_selValid_140 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h04));
  assign _zz_s1_outputPayload_selValid_141 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h04));
  assign _zz_s1_outputPayload_selValid_142 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h04));
  assign _zz_s1_outputPayload_selValid_143 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h04));
  assign _zz_s1_outputPayload_selValid_144 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h04));
  assign _zz_s1_outputPayload_selValid_145 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h04));
  assign _zz_s1_outputPayload_selValid_146 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h04));
  assign _zz_s1_outputPayload_selValid_147 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h04));
  assign _zz_s1_outputPayload_selValid_148 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h04));
  assign _zz_s1_outputPayload_selValid_149 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h04));
  assign _zz_s1_outputPayload_selValid_150 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h04));
  assign _zz_s1_outputPayload_selValid_151 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h04));
  assign _zz_s1_outputPayload_selValid_152 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h04));
  assign _zz_s1_outputPayload_selValid_153 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h04));
  assign _zz_s1_outputPayload_selValid_154 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h04));
  assign _zz_s1_outputPayload_sel_4 = (((((((((((((((_zz_s1_outputPayload_selValid_124 || _zz_s1_outputPayload_selValid_126) || _zz_s1_outputPayload_selValid_128) || _zz_s1_outputPayload_selValid_130) || _zz_s1_outputPayload_selValid_132) || _zz_s1_outputPayload_selValid_134) || _zz_s1_outputPayload_selValid_136) || _zz_s1_outputPayload_selValid_138) || _zz_s1_outputPayload_selValid_140) || _zz_s1_outputPayload_selValid_142) || _zz_s1_outputPayload_selValid_144) || _zz_s1_outputPayload_selValid_146) || _zz_s1_outputPayload_selValid_148) || _zz_s1_outputPayload_selValid_150) || _zz_s1_outputPayload_selValid_152) || _zz_s1_outputPayload_selValid_154);
  assign _zz_s1_outputPayload_sel_4_1 = (((((((((((((((_zz_s1_outputPayload_selValid_125 || _zz_s1_outputPayload_selValid_126) || _zz_s1_outputPayload_selValid_129) || _zz_s1_outputPayload_selValid_130) || _zz_s1_outputPayload_selValid_133) || _zz_s1_outputPayload_selValid_134) || _zz_s1_outputPayload_selValid_137) || _zz_s1_outputPayload_selValid_138) || _zz_s1_outputPayload_selValid_141) || _zz_s1_outputPayload_selValid_142) || _zz_s1_outputPayload_selValid_145) || _zz_s1_outputPayload_selValid_146) || _zz_s1_outputPayload_selValid_149) || _zz_s1_outputPayload_selValid_150) || _zz_s1_outputPayload_selValid_153) || _zz_s1_outputPayload_selValid_154);
  assign _zz_s1_outputPayload_sel_4_2 = (((((((((((((((_zz_s1_outputPayload_selValid_127 || _zz_s1_outputPayload_selValid_128) || _zz_s1_outputPayload_selValid_129) || _zz_s1_outputPayload_selValid_130) || _zz_s1_outputPayload_selValid_135) || _zz_s1_outputPayload_selValid_136) || _zz_s1_outputPayload_selValid_137) || _zz_s1_outputPayload_selValid_138) || _zz_s1_outputPayload_selValid_143) || _zz_s1_outputPayload_selValid_144) || _zz_s1_outputPayload_selValid_145) || _zz_s1_outputPayload_selValid_146) || _zz_s1_outputPayload_selValid_151) || _zz_s1_outputPayload_selValid_152) || _zz_s1_outputPayload_selValid_153) || _zz_s1_outputPayload_selValid_154);
  assign _zz_s1_outputPayload_sel_4_3 = (((((((((((((((_zz_s1_outputPayload_selValid_131 || _zz_s1_outputPayload_selValid_132) || _zz_s1_outputPayload_selValid_133) || _zz_s1_outputPayload_selValid_134) || _zz_s1_outputPayload_selValid_135) || _zz_s1_outputPayload_selValid_136) || _zz_s1_outputPayload_selValid_137) || _zz_s1_outputPayload_selValid_138) || _zz_s1_outputPayload_selValid_147) || _zz_s1_outputPayload_selValid_148) || _zz_s1_outputPayload_selValid_149) || _zz_s1_outputPayload_selValid_150) || _zz_s1_outputPayload_selValid_151) || _zz_s1_outputPayload_selValid_152) || _zz_s1_outputPayload_selValid_153) || _zz_s1_outputPayload_selValid_154);
  assign _zz_s1_outputPayload_sel_4_4 = (((((((((((((((_zz_s1_outputPayload_selValid_139 || _zz_s1_outputPayload_selValid_140) || _zz_s1_outputPayload_selValid_141) || _zz_s1_outputPayload_selValid_142) || _zz_s1_outputPayload_selValid_143) || _zz_s1_outputPayload_selValid_144) || _zz_s1_outputPayload_selValid_145) || _zz_s1_outputPayload_selValid_146) || _zz_s1_outputPayload_selValid_147) || _zz_s1_outputPayload_selValid_148) || _zz_s1_outputPayload_selValid_149) || _zz_s1_outputPayload_selValid_150) || _zz_s1_outputPayload_selValid_151) || _zz_s1_outputPayload_selValid_152) || _zz_s1_outputPayload_selValid_153) || _zz_s1_outputPayload_selValid_154);
  assign s1_outputPayload_sel_4 = {_zz_s1_outputPayload_sel_4_4,{_zz_s1_outputPayload_sel_4_3,{_zz_s1_outputPayload_sel_4_2,{_zz_s1_outputPayload_sel_4_1,_zz_s1_outputPayload_sel_4}}}};
  assign _zz_s1_outputPayload_selValid_155 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h05));
  assign _zz_s1_outputPayload_selValid_156 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h05));
  assign _zz_s1_outputPayload_selValid_157 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h05));
  assign _zz_s1_outputPayload_selValid_158 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h05));
  assign _zz_s1_outputPayload_selValid_159 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h05));
  assign _zz_s1_outputPayload_selValid_160 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h05));
  assign _zz_s1_outputPayload_selValid_161 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h05));
  assign _zz_s1_outputPayload_selValid_162 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h05));
  assign _zz_s1_outputPayload_selValid_163 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h05));
  assign _zz_s1_outputPayload_selValid_164 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h05));
  assign _zz_s1_outputPayload_selValid_165 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h05));
  assign _zz_s1_outputPayload_selValid_166 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h05));
  assign _zz_s1_outputPayload_selValid_167 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h05));
  assign _zz_s1_outputPayload_selValid_168 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h05));
  assign _zz_s1_outputPayload_selValid_169 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h05));
  assign _zz_s1_outputPayload_selValid_170 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h05));
  assign _zz_s1_outputPayload_selValid_171 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h05));
  assign _zz_s1_outputPayload_selValid_172 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h05));
  assign _zz_s1_outputPayload_selValid_173 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h05));
  assign _zz_s1_outputPayload_selValid_174 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h05));
  assign _zz_s1_outputPayload_selValid_175 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h05));
  assign _zz_s1_outputPayload_selValid_176 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h05));
  assign _zz_s1_outputPayload_selValid_177 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h05));
  assign _zz_s1_outputPayload_selValid_178 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h05));
  assign _zz_s1_outputPayload_selValid_179 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h05));
  assign _zz_s1_outputPayload_selValid_180 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h05));
  assign _zz_s1_outputPayload_selValid_181 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h05));
  assign _zz_s1_outputPayload_selValid_182 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h05));
  assign _zz_s1_outputPayload_selValid_183 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h05));
  assign _zz_s1_outputPayload_selValid_184 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h05));
  assign _zz_s1_outputPayload_selValid_185 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h05));
  assign _zz_s1_outputPayload_sel_5 = (((((((((((((((_zz_s1_outputPayload_selValid_155 || _zz_s1_outputPayload_selValid_157) || _zz_s1_outputPayload_selValid_159) || _zz_s1_outputPayload_selValid_161) || _zz_s1_outputPayload_selValid_163) || _zz_s1_outputPayload_selValid_165) || _zz_s1_outputPayload_selValid_167) || _zz_s1_outputPayload_selValid_169) || _zz_s1_outputPayload_selValid_171) || _zz_s1_outputPayload_selValid_173) || _zz_s1_outputPayload_selValid_175) || _zz_s1_outputPayload_selValid_177) || _zz_s1_outputPayload_selValid_179) || _zz_s1_outputPayload_selValid_181) || _zz_s1_outputPayload_selValid_183) || _zz_s1_outputPayload_selValid_185);
  assign _zz_s1_outputPayload_sel_5_1 = (((((((((((((((_zz_s1_outputPayload_selValid_156 || _zz_s1_outputPayload_selValid_157) || _zz_s1_outputPayload_selValid_160) || _zz_s1_outputPayload_selValid_161) || _zz_s1_outputPayload_selValid_164) || _zz_s1_outputPayload_selValid_165) || _zz_s1_outputPayload_selValid_168) || _zz_s1_outputPayload_selValid_169) || _zz_s1_outputPayload_selValid_172) || _zz_s1_outputPayload_selValid_173) || _zz_s1_outputPayload_selValid_176) || _zz_s1_outputPayload_selValid_177) || _zz_s1_outputPayload_selValid_180) || _zz_s1_outputPayload_selValid_181) || _zz_s1_outputPayload_selValid_184) || _zz_s1_outputPayload_selValid_185);
  assign _zz_s1_outputPayload_sel_5_2 = (((((((((((((((_zz_s1_outputPayload_selValid_158 || _zz_s1_outputPayload_selValid_159) || _zz_s1_outputPayload_selValid_160) || _zz_s1_outputPayload_selValid_161) || _zz_s1_outputPayload_selValid_166) || _zz_s1_outputPayload_selValid_167) || _zz_s1_outputPayload_selValid_168) || _zz_s1_outputPayload_selValid_169) || _zz_s1_outputPayload_selValid_174) || _zz_s1_outputPayload_selValid_175) || _zz_s1_outputPayload_selValid_176) || _zz_s1_outputPayload_selValid_177) || _zz_s1_outputPayload_selValid_182) || _zz_s1_outputPayload_selValid_183) || _zz_s1_outputPayload_selValid_184) || _zz_s1_outputPayload_selValid_185);
  assign _zz_s1_outputPayload_sel_5_3 = (((((((((((((((_zz_s1_outputPayload_selValid_162 || _zz_s1_outputPayload_selValid_163) || _zz_s1_outputPayload_selValid_164) || _zz_s1_outputPayload_selValid_165) || _zz_s1_outputPayload_selValid_166) || _zz_s1_outputPayload_selValid_167) || _zz_s1_outputPayload_selValid_168) || _zz_s1_outputPayload_selValid_169) || _zz_s1_outputPayload_selValid_178) || _zz_s1_outputPayload_selValid_179) || _zz_s1_outputPayload_selValid_180) || _zz_s1_outputPayload_selValid_181) || _zz_s1_outputPayload_selValid_182) || _zz_s1_outputPayload_selValid_183) || _zz_s1_outputPayload_selValid_184) || _zz_s1_outputPayload_selValid_185);
  assign _zz_s1_outputPayload_sel_5_4 = (((((((((((((((_zz_s1_outputPayload_selValid_170 || _zz_s1_outputPayload_selValid_171) || _zz_s1_outputPayload_selValid_172) || _zz_s1_outputPayload_selValid_173) || _zz_s1_outputPayload_selValid_174) || _zz_s1_outputPayload_selValid_175) || _zz_s1_outputPayload_selValid_176) || _zz_s1_outputPayload_selValid_177) || _zz_s1_outputPayload_selValid_178) || _zz_s1_outputPayload_selValid_179) || _zz_s1_outputPayload_selValid_180) || _zz_s1_outputPayload_selValid_181) || _zz_s1_outputPayload_selValid_182) || _zz_s1_outputPayload_selValid_183) || _zz_s1_outputPayload_selValid_184) || _zz_s1_outputPayload_selValid_185);
  assign s1_outputPayload_sel_5 = {_zz_s1_outputPayload_sel_5_4,{_zz_s1_outputPayload_sel_5_3,{_zz_s1_outputPayload_sel_5_2,{_zz_s1_outputPayload_sel_5_1,_zz_s1_outputPayload_sel_5}}}};
  assign _zz_s1_outputPayload_selValid_186 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h06));
  assign _zz_s1_outputPayload_selValid_187 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h06));
  assign _zz_s1_outputPayload_selValid_188 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h06));
  assign _zz_s1_outputPayload_selValid_189 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h06));
  assign _zz_s1_outputPayload_selValid_190 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h06));
  assign _zz_s1_outputPayload_selValid_191 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h06));
  assign _zz_s1_outputPayload_selValid_192 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h06));
  assign _zz_s1_outputPayload_selValid_193 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h06));
  assign _zz_s1_outputPayload_selValid_194 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h06));
  assign _zz_s1_outputPayload_selValid_195 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h06));
  assign _zz_s1_outputPayload_selValid_196 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h06));
  assign _zz_s1_outputPayload_selValid_197 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h06));
  assign _zz_s1_outputPayload_selValid_198 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h06));
  assign _zz_s1_outputPayload_selValid_199 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h06));
  assign _zz_s1_outputPayload_selValid_200 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h06));
  assign _zz_s1_outputPayload_selValid_201 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h06));
  assign _zz_s1_outputPayload_selValid_202 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h06));
  assign _zz_s1_outputPayload_selValid_203 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h06));
  assign _zz_s1_outputPayload_selValid_204 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h06));
  assign _zz_s1_outputPayload_selValid_205 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h06));
  assign _zz_s1_outputPayload_selValid_206 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h06));
  assign _zz_s1_outputPayload_selValid_207 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h06));
  assign _zz_s1_outputPayload_selValid_208 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h06));
  assign _zz_s1_outputPayload_selValid_209 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h06));
  assign _zz_s1_outputPayload_selValid_210 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h06));
  assign _zz_s1_outputPayload_selValid_211 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h06));
  assign _zz_s1_outputPayload_selValid_212 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h06));
  assign _zz_s1_outputPayload_selValid_213 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h06));
  assign _zz_s1_outputPayload_selValid_214 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h06));
  assign _zz_s1_outputPayload_selValid_215 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h06));
  assign _zz_s1_outputPayload_selValid_216 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h06));
  assign _zz_s1_outputPayload_sel_6 = (((((((((((((((_zz_s1_outputPayload_selValid_186 || _zz_s1_outputPayload_selValid_188) || _zz_s1_outputPayload_selValid_190) || _zz_s1_outputPayload_selValid_192) || _zz_s1_outputPayload_selValid_194) || _zz_s1_outputPayload_selValid_196) || _zz_s1_outputPayload_selValid_198) || _zz_s1_outputPayload_selValid_200) || _zz_s1_outputPayload_selValid_202) || _zz_s1_outputPayload_selValid_204) || _zz_s1_outputPayload_selValid_206) || _zz_s1_outputPayload_selValid_208) || _zz_s1_outputPayload_selValid_210) || _zz_s1_outputPayload_selValid_212) || _zz_s1_outputPayload_selValid_214) || _zz_s1_outputPayload_selValid_216);
  assign _zz_s1_outputPayload_sel_6_1 = (((((((((((((((_zz_s1_outputPayload_selValid_187 || _zz_s1_outputPayload_selValid_188) || _zz_s1_outputPayload_selValid_191) || _zz_s1_outputPayload_selValid_192) || _zz_s1_outputPayload_selValid_195) || _zz_s1_outputPayload_selValid_196) || _zz_s1_outputPayload_selValid_199) || _zz_s1_outputPayload_selValid_200) || _zz_s1_outputPayload_selValid_203) || _zz_s1_outputPayload_selValid_204) || _zz_s1_outputPayload_selValid_207) || _zz_s1_outputPayload_selValid_208) || _zz_s1_outputPayload_selValid_211) || _zz_s1_outputPayload_selValid_212) || _zz_s1_outputPayload_selValid_215) || _zz_s1_outputPayload_selValid_216);
  assign _zz_s1_outputPayload_sel_6_2 = (((((((((((((((_zz_s1_outputPayload_selValid_189 || _zz_s1_outputPayload_selValid_190) || _zz_s1_outputPayload_selValid_191) || _zz_s1_outputPayload_selValid_192) || _zz_s1_outputPayload_selValid_197) || _zz_s1_outputPayload_selValid_198) || _zz_s1_outputPayload_selValid_199) || _zz_s1_outputPayload_selValid_200) || _zz_s1_outputPayload_selValid_205) || _zz_s1_outputPayload_selValid_206) || _zz_s1_outputPayload_selValid_207) || _zz_s1_outputPayload_selValid_208) || _zz_s1_outputPayload_selValid_213) || _zz_s1_outputPayload_selValid_214) || _zz_s1_outputPayload_selValid_215) || _zz_s1_outputPayload_selValid_216);
  assign _zz_s1_outputPayload_sel_6_3 = (((((((((((((((_zz_s1_outputPayload_selValid_193 || _zz_s1_outputPayload_selValid_194) || _zz_s1_outputPayload_selValid_195) || _zz_s1_outputPayload_selValid_196) || _zz_s1_outputPayload_selValid_197) || _zz_s1_outputPayload_selValid_198) || _zz_s1_outputPayload_selValid_199) || _zz_s1_outputPayload_selValid_200) || _zz_s1_outputPayload_selValid_209) || _zz_s1_outputPayload_selValid_210) || _zz_s1_outputPayload_selValid_211) || _zz_s1_outputPayload_selValid_212) || _zz_s1_outputPayload_selValid_213) || _zz_s1_outputPayload_selValid_214) || _zz_s1_outputPayload_selValid_215) || _zz_s1_outputPayload_selValid_216);
  assign _zz_s1_outputPayload_sel_6_4 = (((((((((((((((_zz_s1_outputPayload_selValid_201 || _zz_s1_outputPayload_selValid_202) || _zz_s1_outputPayload_selValid_203) || _zz_s1_outputPayload_selValid_204) || _zz_s1_outputPayload_selValid_205) || _zz_s1_outputPayload_selValid_206) || _zz_s1_outputPayload_selValid_207) || _zz_s1_outputPayload_selValid_208) || _zz_s1_outputPayload_selValid_209) || _zz_s1_outputPayload_selValid_210) || _zz_s1_outputPayload_selValid_211) || _zz_s1_outputPayload_selValid_212) || _zz_s1_outputPayload_selValid_213) || _zz_s1_outputPayload_selValid_214) || _zz_s1_outputPayload_selValid_215) || _zz_s1_outputPayload_selValid_216);
  assign s1_outputPayload_sel_6 = {_zz_s1_outputPayload_sel_6_4,{_zz_s1_outputPayload_sel_6_3,{_zz_s1_outputPayload_sel_6_2,{_zz_s1_outputPayload_sel_6_1,_zz_s1_outputPayload_sel_6}}}};
  assign _zz_s1_outputPayload_selValid_217 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h07));
  assign _zz_s1_outputPayload_selValid_218 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h07));
  assign _zz_s1_outputPayload_selValid_219 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h07));
  assign _zz_s1_outputPayload_selValid_220 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h07));
  assign _zz_s1_outputPayload_selValid_221 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h07));
  assign _zz_s1_outputPayload_selValid_222 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h07));
  assign _zz_s1_outputPayload_selValid_223 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h07));
  assign _zz_s1_outputPayload_selValid_224 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h07));
  assign _zz_s1_outputPayload_selValid_225 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h07));
  assign _zz_s1_outputPayload_selValid_226 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h07));
  assign _zz_s1_outputPayload_selValid_227 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h07));
  assign _zz_s1_outputPayload_selValid_228 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h07));
  assign _zz_s1_outputPayload_selValid_229 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h07));
  assign _zz_s1_outputPayload_selValid_230 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h07));
  assign _zz_s1_outputPayload_selValid_231 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h07));
  assign _zz_s1_outputPayload_selValid_232 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h07));
  assign _zz_s1_outputPayload_selValid_233 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h07));
  assign _zz_s1_outputPayload_selValid_234 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h07));
  assign _zz_s1_outputPayload_selValid_235 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h07));
  assign _zz_s1_outputPayload_selValid_236 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h07));
  assign _zz_s1_outputPayload_selValid_237 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h07));
  assign _zz_s1_outputPayload_selValid_238 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h07));
  assign _zz_s1_outputPayload_selValid_239 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h07));
  assign _zz_s1_outputPayload_selValid_240 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h07));
  assign _zz_s1_outputPayload_selValid_241 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h07));
  assign _zz_s1_outputPayload_selValid_242 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h07));
  assign _zz_s1_outputPayload_selValid_243 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h07));
  assign _zz_s1_outputPayload_selValid_244 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h07));
  assign _zz_s1_outputPayload_selValid_245 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h07));
  assign _zz_s1_outputPayload_selValid_246 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h07));
  assign _zz_s1_outputPayload_selValid_247 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h07));
  assign _zz_s1_outputPayload_sel_7 = (((((((((((((((_zz_s1_outputPayload_selValid_217 || _zz_s1_outputPayload_selValid_219) || _zz_s1_outputPayload_selValid_221) || _zz_s1_outputPayload_selValid_223) || _zz_s1_outputPayload_selValid_225) || _zz_s1_outputPayload_selValid_227) || _zz_s1_outputPayload_selValid_229) || _zz_s1_outputPayload_selValid_231) || _zz_s1_outputPayload_selValid_233) || _zz_s1_outputPayload_selValid_235) || _zz_s1_outputPayload_selValid_237) || _zz_s1_outputPayload_selValid_239) || _zz_s1_outputPayload_selValid_241) || _zz_s1_outputPayload_selValid_243) || _zz_s1_outputPayload_selValid_245) || _zz_s1_outputPayload_selValid_247);
  assign _zz_s1_outputPayload_sel_7_1 = (((((((((((((((_zz_s1_outputPayload_selValid_218 || _zz_s1_outputPayload_selValid_219) || _zz_s1_outputPayload_selValid_222) || _zz_s1_outputPayload_selValid_223) || _zz_s1_outputPayload_selValid_226) || _zz_s1_outputPayload_selValid_227) || _zz_s1_outputPayload_selValid_230) || _zz_s1_outputPayload_selValid_231) || _zz_s1_outputPayload_selValid_234) || _zz_s1_outputPayload_selValid_235) || _zz_s1_outputPayload_selValid_238) || _zz_s1_outputPayload_selValid_239) || _zz_s1_outputPayload_selValid_242) || _zz_s1_outputPayload_selValid_243) || _zz_s1_outputPayload_selValid_246) || _zz_s1_outputPayload_selValid_247);
  assign _zz_s1_outputPayload_sel_7_2 = (((((((((((((((_zz_s1_outputPayload_selValid_220 || _zz_s1_outputPayload_selValid_221) || _zz_s1_outputPayload_selValid_222) || _zz_s1_outputPayload_selValid_223) || _zz_s1_outputPayload_selValid_228) || _zz_s1_outputPayload_selValid_229) || _zz_s1_outputPayload_selValid_230) || _zz_s1_outputPayload_selValid_231) || _zz_s1_outputPayload_selValid_236) || _zz_s1_outputPayload_selValid_237) || _zz_s1_outputPayload_selValid_238) || _zz_s1_outputPayload_selValid_239) || _zz_s1_outputPayload_selValid_244) || _zz_s1_outputPayload_selValid_245) || _zz_s1_outputPayload_selValid_246) || _zz_s1_outputPayload_selValid_247);
  assign _zz_s1_outputPayload_sel_7_3 = (((((((((((((((_zz_s1_outputPayload_selValid_224 || _zz_s1_outputPayload_selValid_225) || _zz_s1_outputPayload_selValid_226) || _zz_s1_outputPayload_selValid_227) || _zz_s1_outputPayload_selValid_228) || _zz_s1_outputPayload_selValid_229) || _zz_s1_outputPayload_selValid_230) || _zz_s1_outputPayload_selValid_231) || _zz_s1_outputPayload_selValid_240) || _zz_s1_outputPayload_selValid_241) || _zz_s1_outputPayload_selValid_242) || _zz_s1_outputPayload_selValid_243) || _zz_s1_outputPayload_selValid_244) || _zz_s1_outputPayload_selValid_245) || _zz_s1_outputPayload_selValid_246) || _zz_s1_outputPayload_selValid_247);
  assign _zz_s1_outputPayload_sel_7_4 = (((((((((((((((_zz_s1_outputPayload_selValid_232 || _zz_s1_outputPayload_selValid_233) || _zz_s1_outputPayload_selValid_234) || _zz_s1_outputPayload_selValid_235) || _zz_s1_outputPayload_selValid_236) || _zz_s1_outputPayload_selValid_237) || _zz_s1_outputPayload_selValid_238) || _zz_s1_outputPayload_selValid_239) || _zz_s1_outputPayload_selValid_240) || _zz_s1_outputPayload_selValid_241) || _zz_s1_outputPayload_selValid_242) || _zz_s1_outputPayload_selValid_243) || _zz_s1_outputPayload_selValid_244) || _zz_s1_outputPayload_selValid_245) || _zz_s1_outputPayload_selValid_246) || _zz_s1_outputPayload_selValid_247);
  assign s1_outputPayload_sel_7 = {_zz_s1_outputPayload_sel_7_4,{_zz_s1_outputPayload_sel_7_3,{_zz_s1_outputPayload_sel_7_2,{_zz_s1_outputPayload_sel_7_1,_zz_s1_outputPayload_sel_7}}}};
  assign _zz_s1_outputPayload_selValid_248 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h08));
  assign _zz_s1_outputPayload_selValid_249 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h08));
  assign _zz_s1_outputPayload_selValid_250 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h08));
  assign _zz_s1_outputPayload_selValid_251 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h08));
  assign _zz_s1_outputPayload_selValid_252 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h08));
  assign _zz_s1_outputPayload_selValid_253 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h08));
  assign _zz_s1_outputPayload_selValid_254 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h08));
  assign _zz_s1_outputPayload_selValid_255 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h08));
  assign _zz_s1_outputPayload_selValid_256 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h08));
  assign _zz_s1_outputPayload_selValid_257 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h08));
  assign _zz_s1_outputPayload_selValid_258 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h08));
  assign _zz_s1_outputPayload_selValid_259 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h08));
  assign _zz_s1_outputPayload_selValid_260 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h08));
  assign _zz_s1_outputPayload_selValid_261 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h08));
  assign _zz_s1_outputPayload_selValid_262 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h08));
  assign _zz_s1_outputPayload_selValid_263 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h08));
  assign _zz_s1_outputPayload_selValid_264 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h08));
  assign _zz_s1_outputPayload_selValid_265 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h08));
  assign _zz_s1_outputPayload_selValid_266 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h08));
  assign _zz_s1_outputPayload_selValid_267 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h08));
  assign _zz_s1_outputPayload_selValid_268 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h08));
  assign _zz_s1_outputPayload_selValid_269 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h08));
  assign _zz_s1_outputPayload_selValid_270 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h08));
  assign _zz_s1_outputPayload_selValid_271 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h08));
  assign _zz_s1_outputPayload_selValid_272 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h08));
  assign _zz_s1_outputPayload_selValid_273 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h08));
  assign _zz_s1_outputPayload_selValid_274 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h08));
  assign _zz_s1_outputPayload_selValid_275 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h08));
  assign _zz_s1_outputPayload_selValid_276 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h08));
  assign _zz_s1_outputPayload_selValid_277 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h08));
  assign _zz_s1_outputPayload_selValid_278 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h08));
  assign _zz_s1_outputPayload_sel_8 = (((((((((((((((_zz_s1_outputPayload_selValid_248 || _zz_s1_outputPayload_selValid_250) || _zz_s1_outputPayload_selValid_252) || _zz_s1_outputPayload_selValid_254) || _zz_s1_outputPayload_selValid_256) || _zz_s1_outputPayload_selValid_258) || _zz_s1_outputPayload_selValid_260) || _zz_s1_outputPayload_selValid_262) || _zz_s1_outputPayload_selValid_264) || _zz_s1_outputPayload_selValid_266) || _zz_s1_outputPayload_selValid_268) || _zz_s1_outputPayload_selValid_270) || _zz_s1_outputPayload_selValid_272) || _zz_s1_outputPayload_selValid_274) || _zz_s1_outputPayload_selValid_276) || _zz_s1_outputPayload_selValid_278);
  assign _zz_s1_outputPayload_sel_8_1 = (((((((((((((((_zz_s1_outputPayload_selValid_249 || _zz_s1_outputPayload_selValid_250) || _zz_s1_outputPayload_selValid_253) || _zz_s1_outputPayload_selValid_254) || _zz_s1_outputPayload_selValid_257) || _zz_s1_outputPayload_selValid_258) || _zz_s1_outputPayload_selValid_261) || _zz_s1_outputPayload_selValid_262) || _zz_s1_outputPayload_selValid_265) || _zz_s1_outputPayload_selValid_266) || _zz_s1_outputPayload_selValid_269) || _zz_s1_outputPayload_selValid_270) || _zz_s1_outputPayload_selValid_273) || _zz_s1_outputPayload_selValid_274) || _zz_s1_outputPayload_selValid_277) || _zz_s1_outputPayload_selValid_278);
  assign _zz_s1_outputPayload_sel_8_2 = (((((((((((((((_zz_s1_outputPayload_selValid_251 || _zz_s1_outputPayload_selValid_252) || _zz_s1_outputPayload_selValid_253) || _zz_s1_outputPayload_selValid_254) || _zz_s1_outputPayload_selValid_259) || _zz_s1_outputPayload_selValid_260) || _zz_s1_outputPayload_selValid_261) || _zz_s1_outputPayload_selValid_262) || _zz_s1_outputPayload_selValid_267) || _zz_s1_outputPayload_selValid_268) || _zz_s1_outputPayload_selValid_269) || _zz_s1_outputPayload_selValid_270) || _zz_s1_outputPayload_selValid_275) || _zz_s1_outputPayload_selValid_276) || _zz_s1_outputPayload_selValid_277) || _zz_s1_outputPayload_selValid_278);
  assign _zz_s1_outputPayload_sel_8_3 = (((((((((((((((_zz_s1_outputPayload_selValid_255 || _zz_s1_outputPayload_selValid_256) || _zz_s1_outputPayload_selValid_257) || _zz_s1_outputPayload_selValid_258) || _zz_s1_outputPayload_selValid_259) || _zz_s1_outputPayload_selValid_260) || _zz_s1_outputPayload_selValid_261) || _zz_s1_outputPayload_selValid_262) || _zz_s1_outputPayload_selValid_271) || _zz_s1_outputPayload_selValid_272) || _zz_s1_outputPayload_selValid_273) || _zz_s1_outputPayload_selValid_274) || _zz_s1_outputPayload_selValid_275) || _zz_s1_outputPayload_selValid_276) || _zz_s1_outputPayload_selValid_277) || _zz_s1_outputPayload_selValid_278);
  assign _zz_s1_outputPayload_sel_8_4 = (((((((((((((((_zz_s1_outputPayload_selValid_263 || _zz_s1_outputPayload_selValid_264) || _zz_s1_outputPayload_selValid_265) || _zz_s1_outputPayload_selValid_266) || _zz_s1_outputPayload_selValid_267) || _zz_s1_outputPayload_selValid_268) || _zz_s1_outputPayload_selValid_269) || _zz_s1_outputPayload_selValid_270) || _zz_s1_outputPayload_selValid_271) || _zz_s1_outputPayload_selValid_272) || _zz_s1_outputPayload_selValid_273) || _zz_s1_outputPayload_selValid_274) || _zz_s1_outputPayload_selValid_275) || _zz_s1_outputPayload_selValid_276) || _zz_s1_outputPayload_selValid_277) || _zz_s1_outputPayload_selValid_278);
  assign s1_outputPayload_sel_8 = {_zz_s1_outputPayload_sel_8_4,{_zz_s1_outputPayload_sel_8_3,{_zz_s1_outputPayload_sel_8_2,{_zz_s1_outputPayload_sel_8_1,_zz_s1_outputPayload_sel_8}}}};
  assign _zz_s1_outputPayload_selValid_279 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h09));
  assign _zz_s1_outputPayload_selValid_280 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h09));
  assign _zz_s1_outputPayload_selValid_281 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h09));
  assign _zz_s1_outputPayload_selValid_282 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h09));
  assign _zz_s1_outputPayload_selValid_283 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h09));
  assign _zz_s1_outputPayload_selValid_284 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h09));
  assign _zz_s1_outputPayload_selValid_285 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h09));
  assign _zz_s1_outputPayload_selValid_286 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h09));
  assign _zz_s1_outputPayload_selValid_287 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h09));
  assign _zz_s1_outputPayload_selValid_288 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h09));
  assign _zz_s1_outputPayload_selValid_289 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h09));
  assign _zz_s1_outputPayload_selValid_290 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h09));
  assign _zz_s1_outputPayload_selValid_291 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h09));
  assign _zz_s1_outputPayload_selValid_292 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h09));
  assign _zz_s1_outputPayload_selValid_293 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h09));
  assign _zz_s1_outputPayload_selValid_294 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h09));
  assign _zz_s1_outputPayload_selValid_295 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h09));
  assign _zz_s1_outputPayload_selValid_296 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h09));
  assign _zz_s1_outputPayload_selValid_297 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h09));
  assign _zz_s1_outputPayload_selValid_298 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h09));
  assign _zz_s1_outputPayload_selValid_299 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h09));
  assign _zz_s1_outputPayload_selValid_300 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h09));
  assign _zz_s1_outputPayload_selValid_301 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h09));
  assign _zz_s1_outputPayload_selValid_302 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h09));
  assign _zz_s1_outputPayload_selValid_303 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h09));
  assign _zz_s1_outputPayload_selValid_304 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h09));
  assign _zz_s1_outputPayload_selValid_305 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h09));
  assign _zz_s1_outputPayload_selValid_306 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h09));
  assign _zz_s1_outputPayload_selValid_307 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h09));
  assign _zz_s1_outputPayload_selValid_308 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h09));
  assign _zz_s1_outputPayload_selValid_309 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h09));
  assign _zz_s1_outputPayload_sel_9 = (((((((((((((((_zz_s1_outputPayload_selValid_279 || _zz_s1_outputPayload_selValid_281) || _zz_s1_outputPayload_selValid_283) || _zz_s1_outputPayload_selValid_285) || _zz_s1_outputPayload_selValid_287) || _zz_s1_outputPayload_selValid_289) || _zz_s1_outputPayload_selValid_291) || _zz_s1_outputPayload_selValid_293) || _zz_s1_outputPayload_selValid_295) || _zz_s1_outputPayload_selValid_297) || _zz_s1_outputPayload_selValid_299) || _zz_s1_outputPayload_selValid_301) || _zz_s1_outputPayload_selValid_303) || _zz_s1_outputPayload_selValid_305) || _zz_s1_outputPayload_selValid_307) || _zz_s1_outputPayload_selValid_309);
  assign _zz_s1_outputPayload_sel_9_1 = (((((((((((((((_zz_s1_outputPayload_selValid_280 || _zz_s1_outputPayload_selValid_281) || _zz_s1_outputPayload_selValid_284) || _zz_s1_outputPayload_selValid_285) || _zz_s1_outputPayload_selValid_288) || _zz_s1_outputPayload_selValid_289) || _zz_s1_outputPayload_selValid_292) || _zz_s1_outputPayload_selValid_293) || _zz_s1_outputPayload_selValid_296) || _zz_s1_outputPayload_selValid_297) || _zz_s1_outputPayload_selValid_300) || _zz_s1_outputPayload_selValid_301) || _zz_s1_outputPayload_selValid_304) || _zz_s1_outputPayload_selValid_305) || _zz_s1_outputPayload_selValid_308) || _zz_s1_outputPayload_selValid_309);
  assign _zz_s1_outputPayload_sel_9_2 = (((((((((((((((_zz_s1_outputPayload_selValid_282 || _zz_s1_outputPayload_selValid_283) || _zz_s1_outputPayload_selValid_284) || _zz_s1_outputPayload_selValid_285) || _zz_s1_outputPayload_selValid_290) || _zz_s1_outputPayload_selValid_291) || _zz_s1_outputPayload_selValid_292) || _zz_s1_outputPayload_selValid_293) || _zz_s1_outputPayload_selValid_298) || _zz_s1_outputPayload_selValid_299) || _zz_s1_outputPayload_selValid_300) || _zz_s1_outputPayload_selValid_301) || _zz_s1_outputPayload_selValid_306) || _zz_s1_outputPayload_selValid_307) || _zz_s1_outputPayload_selValid_308) || _zz_s1_outputPayload_selValid_309);
  assign _zz_s1_outputPayload_sel_9_3 = (((((((((((((((_zz_s1_outputPayload_selValid_286 || _zz_s1_outputPayload_selValid_287) || _zz_s1_outputPayload_selValid_288) || _zz_s1_outputPayload_selValid_289) || _zz_s1_outputPayload_selValid_290) || _zz_s1_outputPayload_selValid_291) || _zz_s1_outputPayload_selValid_292) || _zz_s1_outputPayload_selValid_293) || _zz_s1_outputPayload_selValid_302) || _zz_s1_outputPayload_selValid_303) || _zz_s1_outputPayload_selValid_304) || _zz_s1_outputPayload_selValid_305) || _zz_s1_outputPayload_selValid_306) || _zz_s1_outputPayload_selValid_307) || _zz_s1_outputPayload_selValid_308) || _zz_s1_outputPayload_selValid_309);
  assign _zz_s1_outputPayload_sel_9_4 = (((((((((((((((_zz_s1_outputPayload_selValid_294 || _zz_s1_outputPayload_selValid_295) || _zz_s1_outputPayload_selValid_296) || _zz_s1_outputPayload_selValid_297) || _zz_s1_outputPayload_selValid_298) || _zz_s1_outputPayload_selValid_299) || _zz_s1_outputPayload_selValid_300) || _zz_s1_outputPayload_selValid_301) || _zz_s1_outputPayload_selValid_302) || _zz_s1_outputPayload_selValid_303) || _zz_s1_outputPayload_selValid_304) || _zz_s1_outputPayload_selValid_305) || _zz_s1_outputPayload_selValid_306) || _zz_s1_outputPayload_selValid_307) || _zz_s1_outputPayload_selValid_308) || _zz_s1_outputPayload_selValid_309);
  assign s1_outputPayload_sel_9 = {_zz_s1_outputPayload_sel_9_4,{_zz_s1_outputPayload_sel_9_3,{_zz_s1_outputPayload_sel_9_2,{_zz_s1_outputPayload_sel_9_1,_zz_s1_outputPayload_sel_9}}}};
  assign _zz_s1_outputPayload_selValid_310 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_311 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_312 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_313 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_314 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_315 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_316 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_317 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_318 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_319 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_320 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_321 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_322 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_323 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_324 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_325 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_326 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_327 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_328 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_329 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_330 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_331 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_332 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_333 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_334 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_335 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_336 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_337 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_338 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_339 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h0a));
  assign _zz_s1_outputPayload_selValid_340 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h0a));
  assign _zz_s1_outputPayload_sel_10 = (((((((((((((((_zz_s1_outputPayload_selValid_310 || _zz_s1_outputPayload_selValid_312) || _zz_s1_outputPayload_selValid_314) || _zz_s1_outputPayload_selValid_316) || _zz_s1_outputPayload_selValid_318) || _zz_s1_outputPayload_selValid_320) || _zz_s1_outputPayload_selValid_322) || _zz_s1_outputPayload_selValid_324) || _zz_s1_outputPayload_selValid_326) || _zz_s1_outputPayload_selValid_328) || _zz_s1_outputPayload_selValid_330) || _zz_s1_outputPayload_selValid_332) || _zz_s1_outputPayload_selValid_334) || _zz_s1_outputPayload_selValid_336) || _zz_s1_outputPayload_selValid_338) || _zz_s1_outputPayload_selValid_340);
  assign _zz_s1_outputPayload_sel_10_1 = (((((((((((((((_zz_s1_outputPayload_selValid_311 || _zz_s1_outputPayload_selValid_312) || _zz_s1_outputPayload_selValid_315) || _zz_s1_outputPayload_selValid_316) || _zz_s1_outputPayload_selValid_319) || _zz_s1_outputPayload_selValid_320) || _zz_s1_outputPayload_selValid_323) || _zz_s1_outputPayload_selValid_324) || _zz_s1_outputPayload_selValid_327) || _zz_s1_outputPayload_selValid_328) || _zz_s1_outputPayload_selValid_331) || _zz_s1_outputPayload_selValid_332) || _zz_s1_outputPayload_selValid_335) || _zz_s1_outputPayload_selValid_336) || _zz_s1_outputPayload_selValid_339) || _zz_s1_outputPayload_selValid_340);
  assign _zz_s1_outputPayload_sel_10_2 = (((((((((((((((_zz_s1_outputPayload_selValid_313 || _zz_s1_outputPayload_selValid_314) || _zz_s1_outputPayload_selValid_315) || _zz_s1_outputPayload_selValid_316) || _zz_s1_outputPayload_selValid_321) || _zz_s1_outputPayload_selValid_322) || _zz_s1_outputPayload_selValid_323) || _zz_s1_outputPayload_selValid_324) || _zz_s1_outputPayload_selValid_329) || _zz_s1_outputPayload_selValid_330) || _zz_s1_outputPayload_selValid_331) || _zz_s1_outputPayload_selValid_332) || _zz_s1_outputPayload_selValid_337) || _zz_s1_outputPayload_selValid_338) || _zz_s1_outputPayload_selValid_339) || _zz_s1_outputPayload_selValid_340);
  assign _zz_s1_outputPayload_sel_10_3 = (((((((((((((((_zz_s1_outputPayload_selValid_317 || _zz_s1_outputPayload_selValid_318) || _zz_s1_outputPayload_selValid_319) || _zz_s1_outputPayload_selValid_320) || _zz_s1_outputPayload_selValid_321) || _zz_s1_outputPayload_selValid_322) || _zz_s1_outputPayload_selValid_323) || _zz_s1_outputPayload_selValid_324) || _zz_s1_outputPayload_selValid_333) || _zz_s1_outputPayload_selValid_334) || _zz_s1_outputPayload_selValid_335) || _zz_s1_outputPayload_selValid_336) || _zz_s1_outputPayload_selValid_337) || _zz_s1_outputPayload_selValid_338) || _zz_s1_outputPayload_selValid_339) || _zz_s1_outputPayload_selValid_340);
  assign _zz_s1_outputPayload_sel_10_4 = (((((((((((((((_zz_s1_outputPayload_selValid_325 || _zz_s1_outputPayload_selValid_326) || _zz_s1_outputPayload_selValid_327) || _zz_s1_outputPayload_selValid_328) || _zz_s1_outputPayload_selValid_329) || _zz_s1_outputPayload_selValid_330) || _zz_s1_outputPayload_selValid_331) || _zz_s1_outputPayload_selValid_332) || _zz_s1_outputPayload_selValid_333) || _zz_s1_outputPayload_selValid_334) || _zz_s1_outputPayload_selValid_335) || _zz_s1_outputPayload_selValid_336) || _zz_s1_outputPayload_selValid_337) || _zz_s1_outputPayload_selValid_338) || _zz_s1_outputPayload_selValid_339) || _zz_s1_outputPayload_selValid_340);
  assign s1_outputPayload_sel_10 = {_zz_s1_outputPayload_sel_10_4,{_zz_s1_outputPayload_sel_10_3,{_zz_s1_outputPayload_sel_10_2,{_zz_s1_outputPayload_sel_10_1,_zz_s1_outputPayload_sel_10}}}};
  assign _zz_s1_outputPayload_selValid_341 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_342 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_343 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_344 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_345 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_346 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_347 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_348 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_349 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_350 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_351 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_352 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_353 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_354 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_355 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_356 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_357 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_358 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_359 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_360 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_361 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_362 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_363 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_364 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_365 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_366 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_367 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_368 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_369 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_370 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h0b));
  assign _zz_s1_outputPayload_selValid_371 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h0b));
  assign _zz_s1_outputPayload_sel_11 = (((((((((((((((_zz_s1_outputPayload_selValid_341 || _zz_s1_outputPayload_selValid_343) || _zz_s1_outputPayload_selValid_345) || _zz_s1_outputPayload_selValid_347) || _zz_s1_outputPayload_selValid_349) || _zz_s1_outputPayload_selValid_351) || _zz_s1_outputPayload_selValid_353) || _zz_s1_outputPayload_selValid_355) || _zz_s1_outputPayload_selValid_357) || _zz_s1_outputPayload_selValid_359) || _zz_s1_outputPayload_selValid_361) || _zz_s1_outputPayload_selValid_363) || _zz_s1_outputPayload_selValid_365) || _zz_s1_outputPayload_selValid_367) || _zz_s1_outputPayload_selValid_369) || _zz_s1_outputPayload_selValid_371);
  assign _zz_s1_outputPayload_sel_11_1 = (((((((((((((((_zz_s1_outputPayload_selValid_342 || _zz_s1_outputPayload_selValid_343) || _zz_s1_outputPayload_selValid_346) || _zz_s1_outputPayload_selValid_347) || _zz_s1_outputPayload_selValid_350) || _zz_s1_outputPayload_selValid_351) || _zz_s1_outputPayload_selValid_354) || _zz_s1_outputPayload_selValid_355) || _zz_s1_outputPayload_selValid_358) || _zz_s1_outputPayload_selValid_359) || _zz_s1_outputPayload_selValid_362) || _zz_s1_outputPayload_selValid_363) || _zz_s1_outputPayload_selValid_366) || _zz_s1_outputPayload_selValid_367) || _zz_s1_outputPayload_selValid_370) || _zz_s1_outputPayload_selValid_371);
  assign _zz_s1_outputPayload_sel_11_2 = (((((((((((((((_zz_s1_outputPayload_selValid_344 || _zz_s1_outputPayload_selValid_345) || _zz_s1_outputPayload_selValid_346) || _zz_s1_outputPayload_selValid_347) || _zz_s1_outputPayload_selValid_352) || _zz_s1_outputPayload_selValid_353) || _zz_s1_outputPayload_selValid_354) || _zz_s1_outputPayload_selValid_355) || _zz_s1_outputPayload_selValid_360) || _zz_s1_outputPayload_selValid_361) || _zz_s1_outputPayload_selValid_362) || _zz_s1_outputPayload_selValid_363) || _zz_s1_outputPayload_selValid_368) || _zz_s1_outputPayload_selValid_369) || _zz_s1_outputPayload_selValid_370) || _zz_s1_outputPayload_selValid_371);
  assign _zz_s1_outputPayload_sel_11_3 = (((((((((((((((_zz_s1_outputPayload_selValid_348 || _zz_s1_outputPayload_selValid_349) || _zz_s1_outputPayload_selValid_350) || _zz_s1_outputPayload_selValid_351) || _zz_s1_outputPayload_selValid_352) || _zz_s1_outputPayload_selValid_353) || _zz_s1_outputPayload_selValid_354) || _zz_s1_outputPayload_selValid_355) || _zz_s1_outputPayload_selValid_364) || _zz_s1_outputPayload_selValid_365) || _zz_s1_outputPayload_selValid_366) || _zz_s1_outputPayload_selValid_367) || _zz_s1_outputPayload_selValid_368) || _zz_s1_outputPayload_selValid_369) || _zz_s1_outputPayload_selValid_370) || _zz_s1_outputPayload_selValid_371);
  assign _zz_s1_outputPayload_sel_11_4 = (((((((((((((((_zz_s1_outputPayload_selValid_356 || _zz_s1_outputPayload_selValid_357) || _zz_s1_outputPayload_selValid_358) || _zz_s1_outputPayload_selValid_359) || _zz_s1_outputPayload_selValid_360) || _zz_s1_outputPayload_selValid_361) || _zz_s1_outputPayload_selValid_362) || _zz_s1_outputPayload_selValid_363) || _zz_s1_outputPayload_selValid_364) || _zz_s1_outputPayload_selValid_365) || _zz_s1_outputPayload_selValid_366) || _zz_s1_outputPayload_selValid_367) || _zz_s1_outputPayload_selValid_368) || _zz_s1_outputPayload_selValid_369) || _zz_s1_outputPayload_selValid_370) || _zz_s1_outputPayload_selValid_371);
  assign s1_outputPayload_sel_11 = {_zz_s1_outputPayload_sel_11_4,{_zz_s1_outputPayload_sel_11_3,{_zz_s1_outputPayload_sel_11_2,{_zz_s1_outputPayload_sel_11_1,_zz_s1_outputPayload_sel_11}}}};
  assign _zz_s1_outputPayload_selValid_372 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_373 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_374 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_375 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_376 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_377 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_378 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_379 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_380 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_381 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_382 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_383 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_384 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_385 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_386 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_387 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_388 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_389 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_390 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_391 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_392 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_393 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_394 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_395 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_396 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_397 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_398 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_399 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_400 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_401 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h0c));
  assign _zz_s1_outputPayload_selValid_402 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h0c));
  assign _zz_s1_outputPayload_sel_12 = (((((((((((((((_zz_s1_outputPayload_selValid_372 || _zz_s1_outputPayload_selValid_374) || _zz_s1_outputPayload_selValid_376) || _zz_s1_outputPayload_selValid_378) || _zz_s1_outputPayload_selValid_380) || _zz_s1_outputPayload_selValid_382) || _zz_s1_outputPayload_selValid_384) || _zz_s1_outputPayload_selValid_386) || _zz_s1_outputPayload_selValid_388) || _zz_s1_outputPayload_selValid_390) || _zz_s1_outputPayload_selValid_392) || _zz_s1_outputPayload_selValid_394) || _zz_s1_outputPayload_selValid_396) || _zz_s1_outputPayload_selValid_398) || _zz_s1_outputPayload_selValid_400) || _zz_s1_outputPayload_selValid_402);
  assign _zz_s1_outputPayload_sel_12_1 = (((((((((((((((_zz_s1_outputPayload_selValid_373 || _zz_s1_outputPayload_selValid_374) || _zz_s1_outputPayload_selValid_377) || _zz_s1_outputPayload_selValid_378) || _zz_s1_outputPayload_selValid_381) || _zz_s1_outputPayload_selValid_382) || _zz_s1_outputPayload_selValid_385) || _zz_s1_outputPayload_selValid_386) || _zz_s1_outputPayload_selValid_389) || _zz_s1_outputPayload_selValid_390) || _zz_s1_outputPayload_selValid_393) || _zz_s1_outputPayload_selValid_394) || _zz_s1_outputPayload_selValid_397) || _zz_s1_outputPayload_selValid_398) || _zz_s1_outputPayload_selValid_401) || _zz_s1_outputPayload_selValid_402);
  assign _zz_s1_outputPayload_sel_12_2 = (((((((((((((((_zz_s1_outputPayload_selValid_375 || _zz_s1_outputPayload_selValid_376) || _zz_s1_outputPayload_selValid_377) || _zz_s1_outputPayload_selValid_378) || _zz_s1_outputPayload_selValid_383) || _zz_s1_outputPayload_selValid_384) || _zz_s1_outputPayload_selValid_385) || _zz_s1_outputPayload_selValid_386) || _zz_s1_outputPayload_selValid_391) || _zz_s1_outputPayload_selValid_392) || _zz_s1_outputPayload_selValid_393) || _zz_s1_outputPayload_selValid_394) || _zz_s1_outputPayload_selValid_399) || _zz_s1_outputPayload_selValid_400) || _zz_s1_outputPayload_selValid_401) || _zz_s1_outputPayload_selValid_402);
  assign _zz_s1_outputPayload_sel_12_3 = (((((((((((((((_zz_s1_outputPayload_selValid_379 || _zz_s1_outputPayload_selValid_380) || _zz_s1_outputPayload_selValid_381) || _zz_s1_outputPayload_selValid_382) || _zz_s1_outputPayload_selValid_383) || _zz_s1_outputPayload_selValid_384) || _zz_s1_outputPayload_selValid_385) || _zz_s1_outputPayload_selValid_386) || _zz_s1_outputPayload_selValid_395) || _zz_s1_outputPayload_selValid_396) || _zz_s1_outputPayload_selValid_397) || _zz_s1_outputPayload_selValid_398) || _zz_s1_outputPayload_selValid_399) || _zz_s1_outputPayload_selValid_400) || _zz_s1_outputPayload_selValid_401) || _zz_s1_outputPayload_selValid_402);
  assign _zz_s1_outputPayload_sel_12_4 = (((((((((((((((_zz_s1_outputPayload_selValid_387 || _zz_s1_outputPayload_selValid_388) || _zz_s1_outputPayload_selValid_389) || _zz_s1_outputPayload_selValid_390) || _zz_s1_outputPayload_selValid_391) || _zz_s1_outputPayload_selValid_392) || _zz_s1_outputPayload_selValid_393) || _zz_s1_outputPayload_selValid_394) || _zz_s1_outputPayload_selValid_395) || _zz_s1_outputPayload_selValid_396) || _zz_s1_outputPayload_selValid_397) || _zz_s1_outputPayload_selValid_398) || _zz_s1_outputPayload_selValid_399) || _zz_s1_outputPayload_selValid_400) || _zz_s1_outputPayload_selValid_401) || _zz_s1_outputPayload_selValid_402);
  assign s1_outputPayload_sel_12 = {_zz_s1_outputPayload_sel_12_4,{_zz_s1_outputPayload_sel_12_3,{_zz_s1_outputPayload_sel_12_2,{_zz_s1_outputPayload_sel_12_1,_zz_s1_outputPayload_sel_12}}}};
  assign _zz_s1_outputPayload_selValid_403 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_404 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_405 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_406 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_407 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_408 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_409 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_410 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_411 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_412 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_413 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_414 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_415 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_416 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_417 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_418 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_419 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_420 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_421 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_422 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_423 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_424 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_425 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_426 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_427 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_428 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_429 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_430 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_431 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_432 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h0d));
  assign _zz_s1_outputPayload_selValid_433 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h0d));
  assign _zz_s1_outputPayload_sel_13 = (((((((((((((((_zz_s1_outputPayload_selValid_403 || _zz_s1_outputPayload_selValid_405) || _zz_s1_outputPayload_selValid_407) || _zz_s1_outputPayload_selValid_409) || _zz_s1_outputPayload_selValid_411) || _zz_s1_outputPayload_selValid_413) || _zz_s1_outputPayload_selValid_415) || _zz_s1_outputPayload_selValid_417) || _zz_s1_outputPayload_selValid_419) || _zz_s1_outputPayload_selValid_421) || _zz_s1_outputPayload_selValid_423) || _zz_s1_outputPayload_selValid_425) || _zz_s1_outputPayload_selValid_427) || _zz_s1_outputPayload_selValid_429) || _zz_s1_outputPayload_selValid_431) || _zz_s1_outputPayload_selValid_433);
  assign _zz_s1_outputPayload_sel_13_1 = (((((((((((((((_zz_s1_outputPayload_selValid_404 || _zz_s1_outputPayload_selValid_405) || _zz_s1_outputPayload_selValid_408) || _zz_s1_outputPayload_selValid_409) || _zz_s1_outputPayload_selValid_412) || _zz_s1_outputPayload_selValid_413) || _zz_s1_outputPayload_selValid_416) || _zz_s1_outputPayload_selValid_417) || _zz_s1_outputPayload_selValid_420) || _zz_s1_outputPayload_selValid_421) || _zz_s1_outputPayload_selValid_424) || _zz_s1_outputPayload_selValid_425) || _zz_s1_outputPayload_selValid_428) || _zz_s1_outputPayload_selValid_429) || _zz_s1_outputPayload_selValid_432) || _zz_s1_outputPayload_selValid_433);
  assign _zz_s1_outputPayload_sel_13_2 = (((((((((((((((_zz_s1_outputPayload_selValid_406 || _zz_s1_outputPayload_selValid_407) || _zz_s1_outputPayload_selValid_408) || _zz_s1_outputPayload_selValid_409) || _zz_s1_outputPayload_selValid_414) || _zz_s1_outputPayload_selValid_415) || _zz_s1_outputPayload_selValid_416) || _zz_s1_outputPayload_selValid_417) || _zz_s1_outputPayload_selValid_422) || _zz_s1_outputPayload_selValid_423) || _zz_s1_outputPayload_selValid_424) || _zz_s1_outputPayload_selValid_425) || _zz_s1_outputPayload_selValid_430) || _zz_s1_outputPayload_selValid_431) || _zz_s1_outputPayload_selValid_432) || _zz_s1_outputPayload_selValid_433);
  assign _zz_s1_outputPayload_sel_13_3 = (((((((((((((((_zz_s1_outputPayload_selValid_410 || _zz_s1_outputPayload_selValid_411) || _zz_s1_outputPayload_selValid_412) || _zz_s1_outputPayload_selValid_413) || _zz_s1_outputPayload_selValid_414) || _zz_s1_outputPayload_selValid_415) || _zz_s1_outputPayload_selValid_416) || _zz_s1_outputPayload_selValid_417) || _zz_s1_outputPayload_selValid_426) || _zz_s1_outputPayload_selValid_427) || _zz_s1_outputPayload_selValid_428) || _zz_s1_outputPayload_selValid_429) || _zz_s1_outputPayload_selValid_430) || _zz_s1_outputPayload_selValid_431) || _zz_s1_outputPayload_selValid_432) || _zz_s1_outputPayload_selValid_433);
  assign _zz_s1_outputPayload_sel_13_4 = (((((((((((((((_zz_s1_outputPayload_selValid_418 || _zz_s1_outputPayload_selValid_419) || _zz_s1_outputPayload_selValid_420) || _zz_s1_outputPayload_selValid_421) || _zz_s1_outputPayload_selValid_422) || _zz_s1_outputPayload_selValid_423) || _zz_s1_outputPayload_selValid_424) || _zz_s1_outputPayload_selValid_425) || _zz_s1_outputPayload_selValid_426) || _zz_s1_outputPayload_selValid_427) || _zz_s1_outputPayload_selValid_428) || _zz_s1_outputPayload_selValid_429) || _zz_s1_outputPayload_selValid_430) || _zz_s1_outputPayload_selValid_431) || _zz_s1_outputPayload_selValid_432) || _zz_s1_outputPayload_selValid_433);
  assign s1_outputPayload_sel_13 = {_zz_s1_outputPayload_sel_13_4,{_zz_s1_outputPayload_sel_13_3,{_zz_s1_outputPayload_sel_13_2,{_zz_s1_outputPayload_sel_13_1,_zz_s1_outputPayload_sel_13}}}};
  assign _zz_s1_outputPayload_selValid_434 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_435 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_436 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_437 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_438 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_439 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_440 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_441 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_442 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_443 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_444 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_445 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_446 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_447 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_448 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_449 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_450 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_451 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_452 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_453 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_454 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_455 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_456 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_457 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_458 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_459 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_460 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_461 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_462 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_463 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h0e));
  assign _zz_s1_outputPayload_selValid_464 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h0e));
  assign _zz_s1_outputPayload_sel_14 = (((((((((((((((_zz_s1_outputPayload_selValid_434 || _zz_s1_outputPayload_selValid_436) || _zz_s1_outputPayload_selValid_438) || _zz_s1_outputPayload_selValid_440) || _zz_s1_outputPayload_selValid_442) || _zz_s1_outputPayload_selValid_444) || _zz_s1_outputPayload_selValid_446) || _zz_s1_outputPayload_selValid_448) || _zz_s1_outputPayload_selValid_450) || _zz_s1_outputPayload_selValid_452) || _zz_s1_outputPayload_selValid_454) || _zz_s1_outputPayload_selValid_456) || _zz_s1_outputPayload_selValid_458) || _zz_s1_outputPayload_selValid_460) || _zz_s1_outputPayload_selValid_462) || _zz_s1_outputPayload_selValid_464);
  assign _zz_s1_outputPayload_sel_14_1 = (((((((((((((((_zz_s1_outputPayload_selValid_435 || _zz_s1_outputPayload_selValid_436) || _zz_s1_outputPayload_selValid_439) || _zz_s1_outputPayload_selValid_440) || _zz_s1_outputPayload_selValid_443) || _zz_s1_outputPayload_selValid_444) || _zz_s1_outputPayload_selValid_447) || _zz_s1_outputPayload_selValid_448) || _zz_s1_outputPayload_selValid_451) || _zz_s1_outputPayload_selValid_452) || _zz_s1_outputPayload_selValid_455) || _zz_s1_outputPayload_selValid_456) || _zz_s1_outputPayload_selValid_459) || _zz_s1_outputPayload_selValid_460) || _zz_s1_outputPayload_selValid_463) || _zz_s1_outputPayload_selValid_464);
  assign _zz_s1_outputPayload_sel_14_2 = (((((((((((((((_zz_s1_outputPayload_selValid_437 || _zz_s1_outputPayload_selValid_438) || _zz_s1_outputPayload_selValid_439) || _zz_s1_outputPayload_selValid_440) || _zz_s1_outputPayload_selValid_445) || _zz_s1_outputPayload_selValid_446) || _zz_s1_outputPayload_selValid_447) || _zz_s1_outputPayload_selValid_448) || _zz_s1_outputPayload_selValid_453) || _zz_s1_outputPayload_selValid_454) || _zz_s1_outputPayload_selValid_455) || _zz_s1_outputPayload_selValid_456) || _zz_s1_outputPayload_selValid_461) || _zz_s1_outputPayload_selValid_462) || _zz_s1_outputPayload_selValid_463) || _zz_s1_outputPayload_selValid_464);
  assign _zz_s1_outputPayload_sel_14_3 = (((((((((((((((_zz_s1_outputPayload_selValid_441 || _zz_s1_outputPayload_selValid_442) || _zz_s1_outputPayload_selValid_443) || _zz_s1_outputPayload_selValid_444) || _zz_s1_outputPayload_selValid_445) || _zz_s1_outputPayload_selValid_446) || _zz_s1_outputPayload_selValid_447) || _zz_s1_outputPayload_selValid_448) || _zz_s1_outputPayload_selValid_457) || _zz_s1_outputPayload_selValid_458) || _zz_s1_outputPayload_selValid_459) || _zz_s1_outputPayload_selValid_460) || _zz_s1_outputPayload_selValid_461) || _zz_s1_outputPayload_selValid_462) || _zz_s1_outputPayload_selValid_463) || _zz_s1_outputPayload_selValid_464);
  assign _zz_s1_outputPayload_sel_14_4 = (((((((((((((((_zz_s1_outputPayload_selValid_449 || _zz_s1_outputPayload_selValid_450) || _zz_s1_outputPayload_selValid_451) || _zz_s1_outputPayload_selValid_452) || _zz_s1_outputPayload_selValid_453) || _zz_s1_outputPayload_selValid_454) || _zz_s1_outputPayload_selValid_455) || _zz_s1_outputPayload_selValid_456) || _zz_s1_outputPayload_selValid_457) || _zz_s1_outputPayload_selValid_458) || _zz_s1_outputPayload_selValid_459) || _zz_s1_outputPayload_selValid_460) || _zz_s1_outputPayload_selValid_461) || _zz_s1_outputPayload_selValid_462) || _zz_s1_outputPayload_selValid_463) || _zz_s1_outputPayload_selValid_464);
  assign s1_outputPayload_sel_14 = {_zz_s1_outputPayload_sel_14_4,{_zz_s1_outputPayload_sel_14_3,{_zz_s1_outputPayload_sel_14_2,{_zz_s1_outputPayload_sel_14_1,_zz_s1_outputPayload_sel_14}}}};
  assign _zz_s1_outputPayload_selValid_465 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_466 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_467 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_468 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_469 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_470 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_471 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_472 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_473 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_474 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_475 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_476 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_477 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_478 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_479 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_480 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_481 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_482 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_483 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_484 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_485 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_486 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_487 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_488 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_489 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_490 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_491 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_492 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_493 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_494 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h0f));
  assign _zz_s1_outputPayload_selValid_495 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h0f));
  assign _zz_s1_outputPayload_sel_15 = (((((((((((((((_zz_s1_outputPayload_selValid_465 || _zz_s1_outputPayload_selValid_467) || _zz_s1_outputPayload_selValid_469) || _zz_s1_outputPayload_selValid_471) || _zz_s1_outputPayload_selValid_473) || _zz_s1_outputPayload_selValid_475) || _zz_s1_outputPayload_selValid_477) || _zz_s1_outputPayload_selValid_479) || _zz_s1_outputPayload_selValid_481) || _zz_s1_outputPayload_selValid_483) || _zz_s1_outputPayload_selValid_485) || _zz_s1_outputPayload_selValid_487) || _zz_s1_outputPayload_selValid_489) || _zz_s1_outputPayload_selValid_491) || _zz_s1_outputPayload_selValid_493) || _zz_s1_outputPayload_selValid_495);
  assign _zz_s1_outputPayload_sel_15_1 = (((((((((((((((_zz_s1_outputPayload_selValid_466 || _zz_s1_outputPayload_selValid_467) || _zz_s1_outputPayload_selValid_470) || _zz_s1_outputPayload_selValid_471) || _zz_s1_outputPayload_selValid_474) || _zz_s1_outputPayload_selValid_475) || _zz_s1_outputPayload_selValid_478) || _zz_s1_outputPayload_selValid_479) || _zz_s1_outputPayload_selValid_482) || _zz_s1_outputPayload_selValid_483) || _zz_s1_outputPayload_selValid_486) || _zz_s1_outputPayload_selValid_487) || _zz_s1_outputPayload_selValid_490) || _zz_s1_outputPayload_selValid_491) || _zz_s1_outputPayload_selValid_494) || _zz_s1_outputPayload_selValid_495);
  assign _zz_s1_outputPayload_sel_15_2 = (((((((((((((((_zz_s1_outputPayload_selValid_468 || _zz_s1_outputPayload_selValid_469) || _zz_s1_outputPayload_selValid_470) || _zz_s1_outputPayload_selValid_471) || _zz_s1_outputPayload_selValid_476) || _zz_s1_outputPayload_selValid_477) || _zz_s1_outputPayload_selValid_478) || _zz_s1_outputPayload_selValid_479) || _zz_s1_outputPayload_selValid_484) || _zz_s1_outputPayload_selValid_485) || _zz_s1_outputPayload_selValid_486) || _zz_s1_outputPayload_selValid_487) || _zz_s1_outputPayload_selValid_492) || _zz_s1_outputPayload_selValid_493) || _zz_s1_outputPayload_selValid_494) || _zz_s1_outputPayload_selValid_495);
  assign _zz_s1_outputPayload_sel_15_3 = (((((((((((((((_zz_s1_outputPayload_selValid_472 || _zz_s1_outputPayload_selValid_473) || _zz_s1_outputPayload_selValid_474) || _zz_s1_outputPayload_selValid_475) || _zz_s1_outputPayload_selValid_476) || _zz_s1_outputPayload_selValid_477) || _zz_s1_outputPayload_selValid_478) || _zz_s1_outputPayload_selValid_479) || _zz_s1_outputPayload_selValid_488) || _zz_s1_outputPayload_selValid_489) || _zz_s1_outputPayload_selValid_490) || _zz_s1_outputPayload_selValid_491) || _zz_s1_outputPayload_selValid_492) || _zz_s1_outputPayload_selValid_493) || _zz_s1_outputPayload_selValid_494) || _zz_s1_outputPayload_selValid_495);
  assign _zz_s1_outputPayload_sel_15_4 = (((((((((((((((_zz_s1_outputPayload_selValid_480 || _zz_s1_outputPayload_selValid_481) || _zz_s1_outputPayload_selValid_482) || _zz_s1_outputPayload_selValid_483) || _zz_s1_outputPayload_selValid_484) || _zz_s1_outputPayload_selValid_485) || _zz_s1_outputPayload_selValid_486) || _zz_s1_outputPayload_selValid_487) || _zz_s1_outputPayload_selValid_488) || _zz_s1_outputPayload_selValid_489) || _zz_s1_outputPayload_selValid_490) || _zz_s1_outputPayload_selValid_491) || _zz_s1_outputPayload_selValid_492) || _zz_s1_outputPayload_selValid_493) || _zz_s1_outputPayload_selValid_494) || _zz_s1_outputPayload_selValid_495);
  assign s1_outputPayload_sel_15 = {_zz_s1_outputPayload_sel_15_4,{_zz_s1_outputPayload_sel_15_3,{_zz_s1_outputPayload_sel_15_2,{_zz_s1_outputPayload_sel_15_1,_zz_s1_outputPayload_sel_15}}}};
  assign _zz_s1_outputPayload_selValid_496 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h10));
  assign _zz_s1_outputPayload_selValid_497 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h10));
  assign _zz_s1_outputPayload_selValid_498 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h10));
  assign _zz_s1_outputPayload_selValid_499 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h10));
  assign _zz_s1_outputPayload_selValid_500 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h10));
  assign _zz_s1_outputPayload_selValid_501 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h10));
  assign _zz_s1_outputPayload_selValid_502 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h10));
  assign _zz_s1_outputPayload_selValid_503 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h10));
  assign _zz_s1_outputPayload_selValid_504 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h10));
  assign _zz_s1_outputPayload_selValid_505 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h10));
  assign _zz_s1_outputPayload_selValid_506 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h10));
  assign _zz_s1_outputPayload_selValid_507 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h10));
  assign _zz_s1_outputPayload_selValid_508 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h10));
  assign _zz_s1_outputPayload_selValid_509 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h10));
  assign _zz_s1_outputPayload_selValid_510 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h10));
  assign _zz_s1_outputPayload_selValid_511 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h10));
  assign _zz_s1_outputPayload_selValid_512 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h10));
  assign _zz_s1_outputPayload_selValid_513 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h10));
  assign _zz_s1_outputPayload_selValid_514 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h10));
  assign _zz_s1_outputPayload_selValid_515 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h10));
  assign _zz_s1_outputPayload_selValid_516 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h10));
  assign _zz_s1_outputPayload_selValid_517 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h10));
  assign _zz_s1_outputPayload_selValid_518 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h10));
  assign _zz_s1_outputPayload_selValid_519 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h10));
  assign _zz_s1_outputPayload_selValid_520 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h10));
  assign _zz_s1_outputPayload_selValid_521 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h10));
  assign _zz_s1_outputPayload_selValid_522 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h10));
  assign _zz_s1_outputPayload_selValid_523 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h10));
  assign _zz_s1_outputPayload_selValid_524 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h10));
  assign _zz_s1_outputPayload_selValid_525 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h10));
  assign _zz_s1_outputPayload_selValid_526 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h10));
  assign _zz_s1_outputPayload_sel_16 = (((((((((((((((_zz_s1_outputPayload_selValid_496 || _zz_s1_outputPayload_selValid_498) || _zz_s1_outputPayload_selValid_500) || _zz_s1_outputPayload_selValid_502) || _zz_s1_outputPayload_selValid_504) || _zz_s1_outputPayload_selValid_506) || _zz_s1_outputPayload_selValid_508) || _zz_s1_outputPayload_selValid_510) || _zz_s1_outputPayload_selValid_512) || _zz_s1_outputPayload_selValid_514) || _zz_s1_outputPayload_selValid_516) || _zz_s1_outputPayload_selValid_518) || _zz_s1_outputPayload_selValid_520) || _zz_s1_outputPayload_selValid_522) || _zz_s1_outputPayload_selValid_524) || _zz_s1_outputPayload_selValid_526);
  assign _zz_s1_outputPayload_sel_16_1 = (((((((((((((((_zz_s1_outputPayload_selValid_497 || _zz_s1_outputPayload_selValid_498) || _zz_s1_outputPayload_selValid_501) || _zz_s1_outputPayload_selValid_502) || _zz_s1_outputPayload_selValid_505) || _zz_s1_outputPayload_selValid_506) || _zz_s1_outputPayload_selValid_509) || _zz_s1_outputPayload_selValid_510) || _zz_s1_outputPayload_selValid_513) || _zz_s1_outputPayload_selValid_514) || _zz_s1_outputPayload_selValid_517) || _zz_s1_outputPayload_selValid_518) || _zz_s1_outputPayload_selValid_521) || _zz_s1_outputPayload_selValid_522) || _zz_s1_outputPayload_selValid_525) || _zz_s1_outputPayload_selValid_526);
  assign _zz_s1_outputPayload_sel_16_2 = (((((((((((((((_zz_s1_outputPayload_selValid_499 || _zz_s1_outputPayload_selValid_500) || _zz_s1_outputPayload_selValid_501) || _zz_s1_outputPayload_selValid_502) || _zz_s1_outputPayload_selValid_507) || _zz_s1_outputPayload_selValid_508) || _zz_s1_outputPayload_selValid_509) || _zz_s1_outputPayload_selValid_510) || _zz_s1_outputPayload_selValid_515) || _zz_s1_outputPayload_selValid_516) || _zz_s1_outputPayload_selValid_517) || _zz_s1_outputPayload_selValid_518) || _zz_s1_outputPayload_selValid_523) || _zz_s1_outputPayload_selValid_524) || _zz_s1_outputPayload_selValid_525) || _zz_s1_outputPayload_selValid_526);
  assign _zz_s1_outputPayload_sel_16_3 = (((((((((((((((_zz_s1_outputPayload_selValid_503 || _zz_s1_outputPayload_selValid_504) || _zz_s1_outputPayload_selValid_505) || _zz_s1_outputPayload_selValid_506) || _zz_s1_outputPayload_selValid_507) || _zz_s1_outputPayload_selValid_508) || _zz_s1_outputPayload_selValid_509) || _zz_s1_outputPayload_selValid_510) || _zz_s1_outputPayload_selValid_519) || _zz_s1_outputPayload_selValid_520) || _zz_s1_outputPayload_selValid_521) || _zz_s1_outputPayload_selValid_522) || _zz_s1_outputPayload_selValid_523) || _zz_s1_outputPayload_selValid_524) || _zz_s1_outputPayload_selValid_525) || _zz_s1_outputPayload_selValid_526);
  assign _zz_s1_outputPayload_sel_16_4 = (((((((((((((((_zz_s1_outputPayload_selValid_511 || _zz_s1_outputPayload_selValid_512) || _zz_s1_outputPayload_selValid_513) || _zz_s1_outputPayload_selValid_514) || _zz_s1_outputPayload_selValid_515) || _zz_s1_outputPayload_selValid_516) || _zz_s1_outputPayload_selValid_517) || _zz_s1_outputPayload_selValid_518) || _zz_s1_outputPayload_selValid_519) || _zz_s1_outputPayload_selValid_520) || _zz_s1_outputPayload_selValid_521) || _zz_s1_outputPayload_selValid_522) || _zz_s1_outputPayload_selValid_523) || _zz_s1_outputPayload_selValid_524) || _zz_s1_outputPayload_selValid_525) || _zz_s1_outputPayload_selValid_526);
  assign s1_outputPayload_sel_16 = {_zz_s1_outputPayload_sel_16_4,{_zz_s1_outputPayload_sel_16_3,{_zz_s1_outputPayload_sel_16_2,{_zz_s1_outputPayload_sel_16_1,_zz_s1_outputPayload_sel_16}}}};
  assign _zz_s1_outputPayload_selValid_527 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h11));
  assign _zz_s1_outputPayload_selValid_528 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h11));
  assign _zz_s1_outputPayload_selValid_529 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h11));
  assign _zz_s1_outputPayload_selValid_530 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h11));
  assign _zz_s1_outputPayload_selValid_531 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h11));
  assign _zz_s1_outputPayload_selValid_532 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h11));
  assign _zz_s1_outputPayload_selValid_533 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h11));
  assign _zz_s1_outputPayload_selValid_534 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h11));
  assign _zz_s1_outputPayload_selValid_535 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h11));
  assign _zz_s1_outputPayload_selValid_536 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h11));
  assign _zz_s1_outputPayload_selValid_537 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h11));
  assign _zz_s1_outputPayload_selValid_538 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h11));
  assign _zz_s1_outputPayload_selValid_539 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h11));
  assign _zz_s1_outputPayload_selValid_540 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h11));
  assign _zz_s1_outputPayload_selValid_541 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h11));
  assign _zz_s1_outputPayload_selValid_542 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h11));
  assign _zz_s1_outputPayload_selValid_543 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h11));
  assign _zz_s1_outputPayload_selValid_544 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h11));
  assign _zz_s1_outputPayload_selValid_545 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h11));
  assign _zz_s1_outputPayload_selValid_546 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h11));
  assign _zz_s1_outputPayload_selValid_547 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h11));
  assign _zz_s1_outputPayload_selValid_548 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h11));
  assign _zz_s1_outputPayload_selValid_549 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h11));
  assign _zz_s1_outputPayload_selValid_550 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h11));
  assign _zz_s1_outputPayload_selValid_551 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h11));
  assign _zz_s1_outputPayload_selValid_552 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h11));
  assign _zz_s1_outputPayload_selValid_553 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h11));
  assign _zz_s1_outputPayload_selValid_554 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h11));
  assign _zz_s1_outputPayload_selValid_555 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h11));
  assign _zz_s1_outputPayload_selValid_556 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h11));
  assign _zz_s1_outputPayload_selValid_557 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h11));
  assign _zz_s1_outputPayload_sel_17 = (((((((((((((((_zz_s1_outputPayload_selValid_527 || _zz_s1_outputPayload_selValid_529) || _zz_s1_outputPayload_selValid_531) || _zz_s1_outputPayload_selValid_533) || _zz_s1_outputPayload_selValid_535) || _zz_s1_outputPayload_selValid_537) || _zz_s1_outputPayload_selValid_539) || _zz_s1_outputPayload_selValid_541) || _zz_s1_outputPayload_selValid_543) || _zz_s1_outputPayload_selValid_545) || _zz_s1_outputPayload_selValid_547) || _zz_s1_outputPayload_selValid_549) || _zz_s1_outputPayload_selValid_551) || _zz_s1_outputPayload_selValid_553) || _zz_s1_outputPayload_selValid_555) || _zz_s1_outputPayload_selValid_557);
  assign _zz_s1_outputPayload_sel_17_1 = (((((((((((((((_zz_s1_outputPayload_selValid_528 || _zz_s1_outputPayload_selValid_529) || _zz_s1_outputPayload_selValid_532) || _zz_s1_outputPayload_selValid_533) || _zz_s1_outputPayload_selValid_536) || _zz_s1_outputPayload_selValid_537) || _zz_s1_outputPayload_selValid_540) || _zz_s1_outputPayload_selValid_541) || _zz_s1_outputPayload_selValid_544) || _zz_s1_outputPayload_selValid_545) || _zz_s1_outputPayload_selValid_548) || _zz_s1_outputPayload_selValid_549) || _zz_s1_outputPayload_selValid_552) || _zz_s1_outputPayload_selValid_553) || _zz_s1_outputPayload_selValid_556) || _zz_s1_outputPayload_selValid_557);
  assign _zz_s1_outputPayload_sel_17_2 = (((((((((((((((_zz_s1_outputPayload_selValid_530 || _zz_s1_outputPayload_selValid_531) || _zz_s1_outputPayload_selValid_532) || _zz_s1_outputPayload_selValid_533) || _zz_s1_outputPayload_selValid_538) || _zz_s1_outputPayload_selValid_539) || _zz_s1_outputPayload_selValid_540) || _zz_s1_outputPayload_selValid_541) || _zz_s1_outputPayload_selValid_546) || _zz_s1_outputPayload_selValid_547) || _zz_s1_outputPayload_selValid_548) || _zz_s1_outputPayload_selValid_549) || _zz_s1_outputPayload_selValid_554) || _zz_s1_outputPayload_selValid_555) || _zz_s1_outputPayload_selValid_556) || _zz_s1_outputPayload_selValid_557);
  assign _zz_s1_outputPayload_sel_17_3 = (((((((((((((((_zz_s1_outputPayload_selValid_534 || _zz_s1_outputPayload_selValid_535) || _zz_s1_outputPayload_selValid_536) || _zz_s1_outputPayload_selValid_537) || _zz_s1_outputPayload_selValid_538) || _zz_s1_outputPayload_selValid_539) || _zz_s1_outputPayload_selValid_540) || _zz_s1_outputPayload_selValid_541) || _zz_s1_outputPayload_selValid_550) || _zz_s1_outputPayload_selValid_551) || _zz_s1_outputPayload_selValid_552) || _zz_s1_outputPayload_selValid_553) || _zz_s1_outputPayload_selValid_554) || _zz_s1_outputPayload_selValid_555) || _zz_s1_outputPayload_selValid_556) || _zz_s1_outputPayload_selValid_557);
  assign _zz_s1_outputPayload_sel_17_4 = (((((((((((((((_zz_s1_outputPayload_selValid_542 || _zz_s1_outputPayload_selValid_543) || _zz_s1_outputPayload_selValid_544) || _zz_s1_outputPayload_selValid_545) || _zz_s1_outputPayload_selValid_546) || _zz_s1_outputPayload_selValid_547) || _zz_s1_outputPayload_selValid_548) || _zz_s1_outputPayload_selValid_549) || _zz_s1_outputPayload_selValid_550) || _zz_s1_outputPayload_selValid_551) || _zz_s1_outputPayload_selValid_552) || _zz_s1_outputPayload_selValid_553) || _zz_s1_outputPayload_selValid_554) || _zz_s1_outputPayload_selValid_555) || _zz_s1_outputPayload_selValid_556) || _zz_s1_outputPayload_selValid_557);
  assign s1_outputPayload_sel_17 = {_zz_s1_outputPayload_sel_17_4,{_zz_s1_outputPayload_sel_17_3,{_zz_s1_outputPayload_sel_17_2,{_zz_s1_outputPayload_sel_17_1,_zz_s1_outputPayload_sel_17}}}};
  assign _zz_s1_outputPayload_selValid_558 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h12));
  assign _zz_s1_outputPayload_selValid_559 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h12));
  assign _zz_s1_outputPayload_selValid_560 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h12));
  assign _zz_s1_outputPayload_selValid_561 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h12));
  assign _zz_s1_outputPayload_selValid_562 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h12));
  assign _zz_s1_outputPayload_selValid_563 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h12));
  assign _zz_s1_outputPayload_selValid_564 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h12));
  assign _zz_s1_outputPayload_selValid_565 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h12));
  assign _zz_s1_outputPayload_selValid_566 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h12));
  assign _zz_s1_outputPayload_selValid_567 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h12));
  assign _zz_s1_outputPayload_selValid_568 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h12));
  assign _zz_s1_outputPayload_selValid_569 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h12));
  assign _zz_s1_outputPayload_selValid_570 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h12));
  assign _zz_s1_outputPayload_selValid_571 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h12));
  assign _zz_s1_outputPayload_selValid_572 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h12));
  assign _zz_s1_outputPayload_selValid_573 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h12));
  assign _zz_s1_outputPayload_selValid_574 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h12));
  assign _zz_s1_outputPayload_selValid_575 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h12));
  assign _zz_s1_outputPayload_selValid_576 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h12));
  assign _zz_s1_outputPayload_selValid_577 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h12));
  assign _zz_s1_outputPayload_selValid_578 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h12));
  assign _zz_s1_outputPayload_selValid_579 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h12));
  assign _zz_s1_outputPayload_selValid_580 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h12));
  assign _zz_s1_outputPayload_selValid_581 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h12));
  assign _zz_s1_outputPayload_selValid_582 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h12));
  assign _zz_s1_outputPayload_selValid_583 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h12));
  assign _zz_s1_outputPayload_selValid_584 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h12));
  assign _zz_s1_outputPayload_selValid_585 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h12));
  assign _zz_s1_outputPayload_selValid_586 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h12));
  assign _zz_s1_outputPayload_selValid_587 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h12));
  assign _zz_s1_outputPayload_selValid_588 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h12));
  assign _zz_s1_outputPayload_sel_18 = (((((((((((((((_zz_s1_outputPayload_selValid_558 || _zz_s1_outputPayload_selValid_560) || _zz_s1_outputPayload_selValid_562) || _zz_s1_outputPayload_selValid_564) || _zz_s1_outputPayload_selValid_566) || _zz_s1_outputPayload_selValid_568) || _zz_s1_outputPayload_selValid_570) || _zz_s1_outputPayload_selValid_572) || _zz_s1_outputPayload_selValid_574) || _zz_s1_outputPayload_selValid_576) || _zz_s1_outputPayload_selValid_578) || _zz_s1_outputPayload_selValid_580) || _zz_s1_outputPayload_selValid_582) || _zz_s1_outputPayload_selValid_584) || _zz_s1_outputPayload_selValid_586) || _zz_s1_outputPayload_selValid_588);
  assign _zz_s1_outputPayload_sel_18_1 = (((((((((((((((_zz_s1_outputPayload_selValid_559 || _zz_s1_outputPayload_selValid_560) || _zz_s1_outputPayload_selValid_563) || _zz_s1_outputPayload_selValid_564) || _zz_s1_outputPayload_selValid_567) || _zz_s1_outputPayload_selValid_568) || _zz_s1_outputPayload_selValid_571) || _zz_s1_outputPayload_selValid_572) || _zz_s1_outputPayload_selValid_575) || _zz_s1_outputPayload_selValid_576) || _zz_s1_outputPayload_selValid_579) || _zz_s1_outputPayload_selValid_580) || _zz_s1_outputPayload_selValid_583) || _zz_s1_outputPayload_selValid_584) || _zz_s1_outputPayload_selValid_587) || _zz_s1_outputPayload_selValid_588);
  assign _zz_s1_outputPayload_sel_18_2 = (((((((((((((((_zz_s1_outputPayload_selValid_561 || _zz_s1_outputPayload_selValid_562) || _zz_s1_outputPayload_selValid_563) || _zz_s1_outputPayload_selValid_564) || _zz_s1_outputPayload_selValid_569) || _zz_s1_outputPayload_selValid_570) || _zz_s1_outputPayload_selValid_571) || _zz_s1_outputPayload_selValid_572) || _zz_s1_outputPayload_selValid_577) || _zz_s1_outputPayload_selValid_578) || _zz_s1_outputPayload_selValid_579) || _zz_s1_outputPayload_selValid_580) || _zz_s1_outputPayload_selValid_585) || _zz_s1_outputPayload_selValid_586) || _zz_s1_outputPayload_selValid_587) || _zz_s1_outputPayload_selValid_588);
  assign _zz_s1_outputPayload_sel_18_3 = (((((((((((((((_zz_s1_outputPayload_selValid_565 || _zz_s1_outputPayload_selValid_566) || _zz_s1_outputPayload_selValid_567) || _zz_s1_outputPayload_selValid_568) || _zz_s1_outputPayload_selValid_569) || _zz_s1_outputPayload_selValid_570) || _zz_s1_outputPayload_selValid_571) || _zz_s1_outputPayload_selValid_572) || _zz_s1_outputPayload_selValid_581) || _zz_s1_outputPayload_selValid_582) || _zz_s1_outputPayload_selValid_583) || _zz_s1_outputPayload_selValid_584) || _zz_s1_outputPayload_selValid_585) || _zz_s1_outputPayload_selValid_586) || _zz_s1_outputPayload_selValid_587) || _zz_s1_outputPayload_selValid_588);
  assign _zz_s1_outputPayload_sel_18_4 = (((((((((((((((_zz_s1_outputPayload_selValid_573 || _zz_s1_outputPayload_selValid_574) || _zz_s1_outputPayload_selValid_575) || _zz_s1_outputPayload_selValid_576) || _zz_s1_outputPayload_selValid_577) || _zz_s1_outputPayload_selValid_578) || _zz_s1_outputPayload_selValid_579) || _zz_s1_outputPayload_selValid_580) || _zz_s1_outputPayload_selValid_581) || _zz_s1_outputPayload_selValid_582) || _zz_s1_outputPayload_selValid_583) || _zz_s1_outputPayload_selValid_584) || _zz_s1_outputPayload_selValid_585) || _zz_s1_outputPayload_selValid_586) || _zz_s1_outputPayload_selValid_587) || _zz_s1_outputPayload_selValid_588);
  assign s1_outputPayload_sel_18 = {_zz_s1_outputPayload_sel_18_4,{_zz_s1_outputPayload_sel_18_3,{_zz_s1_outputPayload_sel_18_2,{_zz_s1_outputPayload_sel_18_1,_zz_s1_outputPayload_sel_18}}}};
  assign _zz_s1_outputPayload_selValid_589 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h13));
  assign _zz_s1_outputPayload_selValid_590 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h13));
  assign _zz_s1_outputPayload_selValid_591 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h13));
  assign _zz_s1_outputPayload_selValid_592 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h13));
  assign _zz_s1_outputPayload_selValid_593 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h13));
  assign _zz_s1_outputPayload_selValid_594 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h13));
  assign _zz_s1_outputPayload_selValid_595 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h13));
  assign _zz_s1_outputPayload_selValid_596 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h13));
  assign _zz_s1_outputPayload_selValid_597 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h13));
  assign _zz_s1_outputPayload_selValid_598 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h13));
  assign _zz_s1_outputPayload_selValid_599 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h13));
  assign _zz_s1_outputPayload_selValid_600 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h13));
  assign _zz_s1_outputPayload_selValid_601 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h13));
  assign _zz_s1_outputPayload_selValid_602 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h13));
  assign _zz_s1_outputPayload_selValid_603 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h13));
  assign _zz_s1_outputPayload_selValid_604 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h13));
  assign _zz_s1_outputPayload_selValid_605 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h13));
  assign _zz_s1_outputPayload_selValid_606 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h13));
  assign _zz_s1_outputPayload_selValid_607 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h13));
  assign _zz_s1_outputPayload_selValid_608 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h13));
  assign _zz_s1_outputPayload_selValid_609 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h13));
  assign _zz_s1_outputPayload_selValid_610 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h13));
  assign _zz_s1_outputPayload_selValid_611 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h13));
  assign _zz_s1_outputPayload_selValid_612 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h13));
  assign _zz_s1_outputPayload_selValid_613 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h13));
  assign _zz_s1_outputPayload_selValid_614 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h13));
  assign _zz_s1_outputPayload_selValid_615 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h13));
  assign _zz_s1_outputPayload_selValid_616 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h13));
  assign _zz_s1_outputPayload_selValid_617 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h13));
  assign _zz_s1_outputPayload_selValid_618 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h13));
  assign _zz_s1_outputPayload_selValid_619 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h13));
  assign _zz_s1_outputPayload_sel_19 = (((((((((((((((_zz_s1_outputPayload_selValid_589 || _zz_s1_outputPayload_selValid_591) || _zz_s1_outputPayload_selValid_593) || _zz_s1_outputPayload_selValid_595) || _zz_s1_outputPayload_selValid_597) || _zz_s1_outputPayload_selValid_599) || _zz_s1_outputPayload_selValid_601) || _zz_s1_outputPayload_selValid_603) || _zz_s1_outputPayload_selValid_605) || _zz_s1_outputPayload_selValid_607) || _zz_s1_outputPayload_selValid_609) || _zz_s1_outputPayload_selValid_611) || _zz_s1_outputPayload_selValid_613) || _zz_s1_outputPayload_selValid_615) || _zz_s1_outputPayload_selValid_617) || _zz_s1_outputPayload_selValid_619);
  assign _zz_s1_outputPayload_sel_19_1 = (((((((((((((((_zz_s1_outputPayload_selValid_590 || _zz_s1_outputPayload_selValid_591) || _zz_s1_outputPayload_selValid_594) || _zz_s1_outputPayload_selValid_595) || _zz_s1_outputPayload_selValid_598) || _zz_s1_outputPayload_selValid_599) || _zz_s1_outputPayload_selValid_602) || _zz_s1_outputPayload_selValid_603) || _zz_s1_outputPayload_selValid_606) || _zz_s1_outputPayload_selValid_607) || _zz_s1_outputPayload_selValid_610) || _zz_s1_outputPayload_selValid_611) || _zz_s1_outputPayload_selValid_614) || _zz_s1_outputPayload_selValid_615) || _zz_s1_outputPayload_selValid_618) || _zz_s1_outputPayload_selValid_619);
  assign _zz_s1_outputPayload_sel_19_2 = (((((((((((((((_zz_s1_outputPayload_selValid_592 || _zz_s1_outputPayload_selValid_593) || _zz_s1_outputPayload_selValid_594) || _zz_s1_outputPayload_selValid_595) || _zz_s1_outputPayload_selValid_600) || _zz_s1_outputPayload_selValid_601) || _zz_s1_outputPayload_selValid_602) || _zz_s1_outputPayload_selValid_603) || _zz_s1_outputPayload_selValid_608) || _zz_s1_outputPayload_selValid_609) || _zz_s1_outputPayload_selValid_610) || _zz_s1_outputPayload_selValid_611) || _zz_s1_outputPayload_selValid_616) || _zz_s1_outputPayload_selValid_617) || _zz_s1_outputPayload_selValid_618) || _zz_s1_outputPayload_selValid_619);
  assign _zz_s1_outputPayload_sel_19_3 = (((((((((((((((_zz_s1_outputPayload_selValid_596 || _zz_s1_outputPayload_selValid_597) || _zz_s1_outputPayload_selValid_598) || _zz_s1_outputPayload_selValid_599) || _zz_s1_outputPayload_selValid_600) || _zz_s1_outputPayload_selValid_601) || _zz_s1_outputPayload_selValid_602) || _zz_s1_outputPayload_selValid_603) || _zz_s1_outputPayload_selValid_612) || _zz_s1_outputPayload_selValid_613) || _zz_s1_outputPayload_selValid_614) || _zz_s1_outputPayload_selValid_615) || _zz_s1_outputPayload_selValid_616) || _zz_s1_outputPayload_selValid_617) || _zz_s1_outputPayload_selValid_618) || _zz_s1_outputPayload_selValid_619);
  assign _zz_s1_outputPayload_sel_19_4 = (((((((((((((((_zz_s1_outputPayload_selValid_604 || _zz_s1_outputPayload_selValid_605) || _zz_s1_outputPayload_selValid_606) || _zz_s1_outputPayload_selValid_607) || _zz_s1_outputPayload_selValid_608) || _zz_s1_outputPayload_selValid_609) || _zz_s1_outputPayload_selValid_610) || _zz_s1_outputPayload_selValid_611) || _zz_s1_outputPayload_selValid_612) || _zz_s1_outputPayload_selValid_613) || _zz_s1_outputPayload_selValid_614) || _zz_s1_outputPayload_selValid_615) || _zz_s1_outputPayload_selValid_616) || _zz_s1_outputPayload_selValid_617) || _zz_s1_outputPayload_selValid_618) || _zz_s1_outputPayload_selValid_619);
  assign s1_outputPayload_sel_19 = {_zz_s1_outputPayload_sel_19_4,{_zz_s1_outputPayload_sel_19_3,{_zz_s1_outputPayload_sel_19_2,{_zz_s1_outputPayload_sel_19_1,_zz_s1_outputPayload_sel_19}}}};
  assign _zz_s1_outputPayload_selValid_620 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h14));
  assign _zz_s1_outputPayload_selValid_621 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h14));
  assign _zz_s1_outputPayload_selValid_622 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h14));
  assign _zz_s1_outputPayload_selValid_623 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h14));
  assign _zz_s1_outputPayload_selValid_624 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h14));
  assign _zz_s1_outputPayload_selValid_625 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h14));
  assign _zz_s1_outputPayload_selValid_626 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h14));
  assign _zz_s1_outputPayload_selValid_627 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h14));
  assign _zz_s1_outputPayload_selValid_628 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h14));
  assign _zz_s1_outputPayload_selValid_629 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h14));
  assign _zz_s1_outputPayload_selValid_630 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h14));
  assign _zz_s1_outputPayload_selValid_631 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h14));
  assign _zz_s1_outputPayload_selValid_632 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h14));
  assign _zz_s1_outputPayload_selValid_633 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h14));
  assign _zz_s1_outputPayload_selValid_634 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h14));
  assign _zz_s1_outputPayload_selValid_635 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h14));
  assign _zz_s1_outputPayload_selValid_636 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h14));
  assign _zz_s1_outputPayload_selValid_637 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h14));
  assign _zz_s1_outputPayload_selValid_638 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h14));
  assign _zz_s1_outputPayload_selValid_639 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h14));
  assign _zz_s1_outputPayload_selValid_640 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h14));
  assign _zz_s1_outputPayload_selValid_641 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h14));
  assign _zz_s1_outputPayload_selValid_642 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h14));
  assign _zz_s1_outputPayload_selValid_643 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h14));
  assign _zz_s1_outputPayload_selValid_644 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h14));
  assign _zz_s1_outputPayload_selValid_645 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h14));
  assign _zz_s1_outputPayload_selValid_646 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h14));
  assign _zz_s1_outputPayload_selValid_647 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h14));
  assign _zz_s1_outputPayload_selValid_648 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h14));
  assign _zz_s1_outputPayload_selValid_649 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h14));
  assign _zz_s1_outputPayload_selValid_650 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h14));
  assign _zz_s1_outputPayload_sel_20 = (((((((((((((((_zz_s1_outputPayload_selValid_620 || _zz_s1_outputPayload_selValid_622) || _zz_s1_outputPayload_selValid_624) || _zz_s1_outputPayload_selValid_626) || _zz_s1_outputPayload_selValid_628) || _zz_s1_outputPayload_selValid_630) || _zz_s1_outputPayload_selValid_632) || _zz_s1_outputPayload_selValid_634) || _zz_s1_outputPayload_selValid_636) || _zz_s1_outputPayload_selValid_638) || _zz_s1_outputPayload_selValid_640) || _zz_s1_outputPayload_selValid_642) || _zz_s1_outputPayload_selValid_644) || _zz_s1_outputPayload_selValid_646) || _zz_s1_outputPayload_selValid_648) || _zz_s1_outputPayload_selValid_650);
  assign _zz_s1_outputPayload_sel_20_1 = (((((((((((((((_zz_s1_outputPayload_selValid_621 || _zz_s1_outputPayload_selValid_622) || _zz_s1_outputPayload_selValid_625) || _zz_s1_outputPayload_selValid_626) || _zz_s1_outputPayload_selValid_629) || _zz_s1_outputPayload_selValid_630) || _zz_s1_outputPayload_selValid_633) || _zz_s1_outputPayload_selValid_634) || _zz_s1_outputPayload_selValid_637) || _zz_s1_outputPayload_selValid_638) || _zz_s1_outputPayload_selValid_641) || _zz_s1_outputPayload_selValid_642) || _zz_s1_outputPayload_selValid_645) || _zz_s1_outputPayload_selValid_646) || _zz_s1_outputPayload_selValid_649) || _zz_s1_outputPayload_selValid_650);
  assign _zz_s1_outputPayload_sel_20_2 = (((((((((((((((_zz_s1_outputPayload_selValid_623 || _zz_s1_outputPayload_selValid_624) || _zz_s1_outputPayload_selValid_625) || _zz_s1_outputPayload_selValid_626) || _zz_s1_outputPayload_selValid_631) || _zz_s1_outputPayload_selValid_632) || _zz_s1_outputPayload_selValid_633) || _zz_s1_outputPayload_selValid_634) || _zz_s1_outputPayload_selValid_639) || _zz_s1_outputPayload_selValid_640) || _zz_s1_outputPayload_selValid_641) || _zz_s1_outputPayload_selValid_642) || _zz_s1_outputPayload_selValid_647) || _zz_s1_outputPayload_selValid_648) || _zz_s1_outputPayload_selValid_649) || _zz_s1_outputPayload_selValid_650);
  assign _zz_s1_outputPayload_sel_20_3 = (((((((((((((((_zz_s1_outputPayload_selValid_627 || _zz_s1_outputPayload_selValid_628) || _zz_s1_outputPayload_selValid_629) || _zz_s1_outputPayload_selValid_630) || _zz_s1_outputPayload_selValid_631) || _zz_s1_outputPayload_selValid_632) || _zz_s1_outputPayload_selValid_633) || _zz_s1_outputPayload_selValid_634) || _zz_s1_outputPayload_selValid_643) || _zz_s1_outputPayload_selValid_644) || _zz_s1_outputPayload_selValid_645) || _zz_s1_outputPayload_selValid_646) || _zz_s1_outputPayload_selValid_647) || _zz_s1_outputPayload_selValid_648) || _zz_s1_outputPayload_selValid_649) || _zz_s1_outputPayload_selValid_650);
  assign _zz_s1_outputPayload_sel_20_4 = (((((((((((((((_zz_s1_outputPayload_selValid_635 || _zz_s1_outputPayload_selValid_636) || _zz_s1_outputPayload_selValid_637) || _zz_s1_outputPayload_selValid_638) || _zz_s1_outputPayload_selValid_639) || _zz_s1_outputPayload_selValid_640) || _zz_s1_outputPayload_selValid_641) || _zz_s1_outputPayload_selValid_642) || _zz_s1_outputPayload_selValid_643) || _zz_s1_outputPayload_selValid_644) || _zz_s1_outputPayload_selValid_645) || _zz_s1_outputPayload_selValid_646) || _zz_s1_outputPayload_selValid_647) || _zz_s1_outputPayload_selValid_648) || _zz_s1_outputPayload_selValid_649) || _zz_s1_outputPayload_selValid_650);
  assign s1_outputPayload_sel_20 = {_zz_s1_outputPayload_sel_20_4,{_zz_s1_outputPayload_sel_20_3,{_zz_s1_outputPayload_sel_20_2,{_zz_s1_outputPayload_sel_20_1,_zz_s1_outputPayload_sel_20}}}};
  assign _zz_s1_outputPayload_selValid_651 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h15));
  assign _zz_s1_outputPayload_selValid_652 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h15));
  assign _zz_s1_outputPayload_selValid_653 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h15));
  assign _zz_s1_outputPayload_selValid_654 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h15));
  assign _zz_s1_outputPayload_selValid_655 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h15));
  assign _zz_s1_outputPayload_selValid_656 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h15));
  assign _zz_s1_outputPayload_selValid_657 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h15));
  assign _zz_s1_outputPayload_selValid_658 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h15));
  assign _zz_s1_outputPayload_selValid_659 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h15));
  assign _zz_s1_outputPayload_selValid_660 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h15));
  assign _zz_s1_outputPayload_selValid_661 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h15));
  assign _zz_s1_outputPayload_selValid_662 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h15));
  assign _zz_s1_outputPayload_selValid_663 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h15));
  assign _zz_s1_outputPayload_selValid_664 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h15));
  assign _zz_s1_outputPayload_selValid_665 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h15));
  assign _zz_s1_outputPayload_selValid_666 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h15));
  assign _zz_s1_outputPayload_selValid_667 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h15));
  assign _zz_s1_outputPayload_selValid_668 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h15));
  assign _zz_s1_outputPayload_selValid_669 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h15));
  assign _zz_s1_outputPayload_selValid_670 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h15));
  assign _zz_s1_outputPayload_selValid_671 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h15));
  assign _zz_s1_outputPayload_selValid_672 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h15));
  assign _zz_s1_outputPayload_selValid_673 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h15));
  assign _zz_s1_outputPayload_selValid_674 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h15));
  assign _zz_s1_outputPayload_selValid_675 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h15));
  assign _zz_s1_outputPayload_selValid_676 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h15));
  assign _zz_s1_outputPayload_selValid_677 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h15));
  assign _zz_s1_outputPayload_selValid_678 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h15));
  assign _zz_s1_outputPayload_selValid_679 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h15));
  assign _zz_s1_outputPayload_selValid_680 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h15));
  assign _zz_s1_outputPayload_selValid_681 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h15));
  assign _zz_s1_outputPayload_sel_21 = (((((((((((((((_zz_s1_outputPayload_selValid_651 || _zz_s1_outputPayload_selValid_653) || _zz_s1_outputPayload_selValid_655) || _zz_s1_outputPayload_selValid_657) || _zz_s1_outputPayload_selValid_659) || _zz_s1_outputPayload_selValid_661) || _zz_s1_outputPayload_selValid_663) || _zz_s1_outputPayload_selValid_665) || _zz_s1_outputPayload_selValid_667) || _zz_s1_outputPayload_selValid_669) || _zz_s1_outputPayload_selValid_671) || _zz_s1_outputPayload_selValid_673) || _zz_s1_outputPayload_selValid_675) || _zz_s1_outputPayload_selValid_677) || _zz_s1_outputPayload_selValid_679) || _zz_s1_outputPayload_selValid_681);
  assign _zz_s1_outputPayload_sel_21_1 = (((((((((((((((_zz_s1_outputPayload_selValid_652 || _zz_s1_outputPayload_selValid_653) || _zz_s1_outputPayload_selValid_656) || _zz_s1_outputPayload_selValid_657) || _zz_s1_outputPayload_selValid_660) || _zz_s1_outputPayload_selValid_661) || _zz_s1_outputPayload_selValid_664) || _zz_s1_outputPayload_selValid_665) || _zz_s1_outputPayload_selValid_668) || _zz_s1_outputPayload_selValid_669) || _zz_s1_outputPayload_selValid_672) || _zz_s1_outputPayload_selValid_673) || _zz_s1_outputPayload_selValid_676) || _zz_s1_outputPayload_selValid_677) || _zz_s1_outputPayload_selValid_680) || _zz_s1_outputPayload_selValid_681);
  assign _zz_s1_outputPayload_sel_21_2 = (((((((((((((((_zz_s1_outputPayload_selValid_654 || _zz_s1_outputPayload_selValid_655) || _zz_s1_outputPayload_selValid_656) || _zz_s1_outputPayload_selValid_657) || _zz_s1_outputPayload_selValid_662) || _zz_s1_outputPayload_selValid_663) || _zz_s1_outputPayload_selValid_664) || _zz_s1_outputPayload_selValid_665) || _zz_s1_outputPayload_selValid_670) || _zz_s1_outputPayload_selValid_671) || _zz_s1_outputPayload_selValid_672) || _zz_s1_outputPayload_selValid_673) || _zz_s1_outputPayload_selValid_678) || _zz_s1_outputPayload_selValid_679) || _zz_s1_outputPayload_selValid_680) || _zz_s1_outputPayload_selValid_681);
  assign _zz_s1_outputPayload_sel_21_3 = (((((((((((((((_zz_s1_outputPayload_selValid_658 || _zz_s1_outputPayload_selValid_659) || _zz_s1_outputPayload_selValid_660) || _zz_s1_outputPayload_selValid_661) || _zz_s1_outputPayload_selValid_662) || _zz_s1_outputPayload_selValid_663) || _zz_s1_outputPayload_selValid_664) || _zz_s1_outputPayload_selValid_665) || _zz_s1_outputPayload_selValid_674) || _zz_s1_outputPayload_selValid_675) || _zz_s1_outputPayload_selValid_676) || _zz_s1_outputPayload_selValid_677) || _zz_s1_outputPayload_selValid_678) || _zz_s1_outputPayload_selValid_679) || _zz_s1_outputPayload_selValid_680) || _zz_s1_outputPayload_selValid_681);
  assign _zz_s1_outputPayload_sel_21_4 = (((((((((((((((_zz_s1_outputPayload_selValid_666 || _zz_s1_outputPayload_selValid_667) || _zz_s1_outputPayload_selValid_668) || _zz_s1_outputPayload_selValid_669) || _zz_s1_outputPayload_selValid_670) || _zz_s1_outputPayload_selValid_671) || _zz_s1_outputPayload_selValid_672) || _zz_s1_outputPayload_selValid_673) || _zz_s1_outputPayload_selValid_674) || _zz_s1_outputPayload_selValid_675) || _zz_s1_outputPayload_selValid_676) || _zz_s1_outputPayload_selValid_677) || _zz_s1_outputPayload_selValid_678) || _zz_s1_outputPayload_selValid_679) || _zz_s1_outputPayload_selValid_680) || _zz_s1_outputPayload_selValid_681);
  assign s1_outputPayload_sel_21 = {_zz_s1_outputPayload_sel_21_4,{_zz_s1_outputPayload_sel_21_3,{_zz_s1_outputPayload_sel_21_2,{_zz_s1_outputPayload_sel_21_1,_zz_s1_outputPayload_sel_21}}}};
  assign _zz_s1_outputPayload_selValid_682 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h16));
  assign _zz_s1_outputPayload_selValid_683 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h16));
  assign _zz_s1_outputPayload_selValid_684 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h16));
  assign _zz_s1_outputPayload_selValid_685 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h16));
  assign _zz_s1_outputPayload_selValid_686 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h16));
  assign _zz_s1_outputPayload_selValid_687 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h16));
  assign _zz_s1_outputPayload_selValid_688 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h16));
  assign _zz_s1_outputPayload_selValid_689 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h16));
  assign _zz_s1_outputPayload_selValid_690 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h16));
  assign _zz_s1_outputPayload_selValid_691 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h16));
  assign _zz_s1_outputPayload_selValid_692 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h16));
  assign _zz_s1_outputPayload_selValid_693 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h16));
  assign _zz_s1_outputPayload_selValid_694 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h16));
  assign _zz_s1_outputPayload_selValid_695 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h16));
  assign _zz_s1_outputPayload_selValid_696 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h16));
  assign _zz_s1_outputPayload_selValid_697 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h16));
  assign _zz_s1_outputPayload_selValid_698 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h16));
  assign _zz_s1_outputPayload_selValid_699 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h16));
  assign _zz_s1_outputPayload_selValid_700 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h16));
  assign _zz_s1_outputPayload_selValid_701 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h16));
  assign _zz_s1_outputPayload_selValid_702 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h16));
  assign _zz_s1_outputPayload_selValid_703 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h16));
  assign _zz_s1_outputPayload_selValid_704 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h16));
  assign _zz_s1_outputPayload_selValid_705 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h16));
  assign _zz_s1_outputPayload_selValid_706 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h16));
  assign _zz_s1_outputPayload_selValid_707 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h16));
  assign _zz_s1_outputPayload_selValid_708 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h16));
  assign _zz_s1_outputPayload_selValid_709 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h16));
  assign _zz_s1_outputPayload_selValid_710 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h16));
  assign _zz_s1_outputPayload_selValid_711 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h16));
  assign _zz_s1_outputPayload_selValid_712 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h16));
  assign _zz_s1_outputPayload_sel_22 = (((((((((((((((_zz_s1_outputPayload_selValid_682 || _zz_s1_outputPayload_selValid_684) || _zz_s1_outputPayload_selValid_686) || _zz_s1_outputPayload_selValid_688) || _zz_s1_outputPayload_selValid_690) || _zz_s1_outputPayload_selValid_692) || _zz_s1_outputPayload_selValid_694) || _zz_s1_outputPayload_selValid_696) || _zz_s1_outputPayload_selValid_698) || _zz_s1_outputPayload_selValid_700) || _zz_s1_outputPayload_selValid_702) || _zz_s1_outputPayload_selValid_704) || _zz_s1_outputPayload_selValid_706) || _zz_s1_outputPayload_selValid_708) || _zz_s1_outputPayload_selValid_710) || _zz_s1_outputPayload_selValid_712);
  assign _zz_s1_outputPayload_sel_22_1 = (((((((((((((((_zz_s1_outputPayload_selValid_683 || _zz_s1_outputPayload_selValid_684) || _zz_s1_outputPayload_selValid_687) || _zz_s1_outputPayload_selValid_688) || _zz_s1_outputPayload_selValid_691) || _zz_s1_outputPayload_selValid_692) || _zz_s1_outputPayload_selValid_695) || _zz_s1_outputPayload_selValid_696) || _zz_s1_outputPayload_selValid_699) || _zz_s1_outputPayload_selValid_700) || _zz_s1_outputPayload_selValid_703) || _zz_s1_outputPayload_selValid_704) || _zz_s1_outputPayload_selValid_707) || _zz_s1_outputPayload_selValid_708) || _zz_s1_outputPayload_selValid_711) || _zz_s1_outputPayload_selValid_712);
  assign _zz_s1_outputPayload_sel_22_2 = (((((((((((((((_zz_s1_outputPayload_selValid_685 || _zz_s1_outputPayload_selValid_686) || _zz_s1_outputPayload_selValid_687) || _zz_s1_outputPayload_selValid_688) || _zz_s1_outputPayload_selValid_693) || _zz_s1_outputPayload_selValid_694) || _zz_s1_outputPayload_selValid_695) || _zz_s1_outputPayload_selValid_696) || _zz_s1_outputPayload_selValid_701) || _zz_s1_outputPayload_selValid_702) || _zz_s1_outputPayload_selValid_703) || _zz_s1_outputPayload_selValid_704) || _zz_s1_outputPayload_selValid_709) || _zz_s1_outputPayload_selValid_710) || _zz_s1_outputPayload_selValid_711) || _zz_s1_outputPayload_selValid_712);
  assign _zz_s1_outputPayload_sel_22_3 = (((((((((((((((_zz_s1_outputPayload_selValid_689 || _zz_s1_outputPayload_selValid_690) || _zz_s1_outputPayload_selValid_691) || _zz_s1_outputPayload_selValid_692) || _zz_s1_outputPayload_selValid_693) || _zz_s1_outputPayload_selValid_694) || _zz_s1_outputPayload_selValid_695) || _zz_s1_outputPayload_selValid_696) || _zz_s1_outputPayload_selValid_705) || _zz_s1_outputPayload_selValid_706) || _zz_s1_outputPayload_selValid_707) || _zz_s1_outputPayload_selValid_708) || _zz_s1_outputPayload_selValid_709) || _zz_s1_outputPayload_selValid_710) || _zz_s1_outputPayload_selValid_711) || _zz_s1_outputPayload_selValid_712);
  assign _zz_s1_outputPayload_sel_22_4 = (((((((((((((((_zz_s1_outputPayload_selValid_697 || _zz_s1_outputPayload_selValid_698) || _zz_s1_outputPayload_selValid_699) || _zz_s1_outputPayload_selValid_700) || _zz_s1_outputPayload_selValid_701) || _zz_s1_outputPayload_selValid_702) || _zz_s1_outputPayload_selValid_703) || _zz_s1_outputPayload_selValid_704) || _zz_s1_outputPayload_selValid_705) || _zz_s1_outputPayload_selValid_706) || _zz_s1_outputPayload_selValid_707) || _zz_s1_outputPayload_selValid_708) || _zz_s1_outputPayload_selValid_709) || _zz_s1_outputPayload_selValid_710) || _zz_s1_outputPayload_selValid_711) || _zz_s1_outputPayload_selValid_712);
  assign s1_outputPayload_sel_22 = {_zz_s1_outputPayload_sel_22_4,{_zz_s1_outputPayload_sel_22_3,{_zz_s1_outputPayload_sel_22_2,{_zz_s1_outputPayload_sel_22_1,_zz_s1_outputPayload_sel_22}}}};
  assign _zz_s1_outputPayload_selValid_713 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h17));
  assign _zz_s1_outputPayload_selValid_714 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h17));
  assign _zz_s1_outputPayload_selValid_715 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h17));
  assign _zz_s1_outputPayload_selValid_716 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h17));
  assign _zz_s1_outputPayload_selValid_717 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h17));
  assign _zz_s1_outputPayload_selValid_718 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h17));
  assign _zz_s1_outputPayload_selValid_719 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h17));
  assign _zz_s1_outputPayload_selValid_720 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h17));
  assign _zz_s1_outputPayload_selValid_721 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h17));
  assign _zz_s1_outputPayload_selValid_722 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h17));
  assign _zz_s1_outputPayload_selValid_723 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h17));
  assign _zz_s1_outputPayload_selValid_724 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h17));
  assign _zz_s1_outputPayload_selValid_725 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h17));
  assign _zz_s1_outputPayload_selValid_726 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h17));
  assign _zz_s1_outputPayload_selValid_727 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h17));
  assign _zz_s1_outputPayload_selValid_728 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h17));
  assign _zz_s1_outputPayload_selValid_729 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h17));
  assign _zz_s1_outputPayload_selValid_730 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h17));
  assign _zz_s1_outputPayload_selValid_731 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h17));
  assign _zz_s1_outputPayload_selValid_732 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h17));
  assign _zz_s1_outputPayload_selValid_733 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h17));
  assign _zz_s1_outputPayload_selValid_734 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h17));
  assign _zz_s1_outputPayload_selValid_735 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h17));
  assign _zz_s1_outputPayload_selValid_736 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h17));
  assign _zz_s1_outputPayload_selValid_737 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h17));
  assign _zz_s1_outputPayload_selValid_738 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h17));
  assign _zz_s1_outputPayload_selValid_739 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h17));
  assign _zz_s1_outputPayload_selValid_740 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h17));
  assign _zz_s1_outputPayload_selValid_741 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h17));
  assign _zz_s1_outputPayload_selValid_742 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h17));
  assign _zz_s1_outputPayload_selValid_743 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h17));
  assign _zz_s1_outputPayload_sel_23 = (((((((((((((((_zz_s1_outputPayload_selValid_713 || _zz_s1_outputPayload_selValid_715) || _zz_s1_outputPayload_selValid_717) || _zz_s1_outputPayload_selValid_719) || _zz_s1_outputPayload_selValid_721) || _zz_s1_outputPayload_selValid_723) || _zz_s1_outputPayload_selValid_725) || _zz_s1_outputPayload_selValid_727) || _zz_s1_outputPayload_selValid_729) || _zz_s1_outputPayload_selValid_731) || _zz_s1_outputPayload_selValid_733) || _zz_s1_outputPayload_selValid_735) || _zz_s1_outputPayload_selValid_737) || _zz_s1_outputPayload_selValid_739) || _zz_s1_outputPayload_selValid_741) || _zz_s1_outputPayload_selValid_743);
  assign _zz_s1_outputPayload_sel_23_1 = (((((((((((((((_zz_s1_outputPayload_selValid_714 || _zz_s1_outputPayload_selValid_715) || _zz_s1_outputPayload_selValid_718) || _zz_s1_outputPayload_selValid_719) || _zz_s1_outputPayload_selValid_722) || _zz_s1_outputPayload_selValid_723) || _zz_s1_outputPayload_selValid_726) || _zz_s1_outputPayload_selValid_727) || _zz_s1_outputPayload_selValid_730) || _zz_s1_outputPayload_selValid_731) || _zz_s1_outputPayload_selValid_734) || _zz_s1_outputPayload_selValid_735) || _zz_s1_outputPayload_selValid_738) || _zz_s1_outputPayload_selValid_739) || _zz_s1_outputPayload_selValid_742) || _zz_s1_outputPayload_selValid_743);
  assign _zz_s1_outputPayload_sel_23_2 = (((((((((((((((_zz_s1_outputPayload_selValid_716 || _zz_s1_outputPayload_selValid_717) || _zz_s1_outputPayload_selValid_718) || _zz_s1_outputPayload_selValid_719) || _zz_s1_outputPayload_selValid_724) || _zz_s1_outputPayload_selValid_725) || _zz_s1_outputPayload_selValid_726) || _zz_s1_outputPayload_selValid_727) || _zz_s1_outputPayload_selValid_732) || _zz_s1_outputPayload_selValid_733) || _zz_s1_outputPayload_selValid_734) || _zz_s1_outputPayload_selValid_735) || _zz_s1_outputPayload_selValid_740) || _zz_s1_outputPayload_selValid_741) || _zz_s1_outputPayload_selValid_742) || _zz_s1_outputPayload_selValid_743);
  assign _zz_s1_outputPayload_sel_23_3 = (((((((((((((((_zz_s1_outputPayload_selValid_720 || _zz_s1_outputPayload_selValid_721) || _zz_s1_outputPayload_selValid_722) || _zz_s1_outputPayload_selValid_723) || _zz_s1_outputPayload_selValid_724) || _zz_s1_outputPayload_selValid_725) || _zz_s1_outputPayload_selValid_726) || _zz_s1_outputPayload_selValid_727) || _zz_s1_outputPayload_selValid_736) || _zz_s1_outputPayload_selValid_737) || _zz_s1_outputPayload_selValid_738) || _zz_s1_outputPayload_selValid_739) || _zz_s1_outputPayload_selValid_740) || _zz_s1_outputPayload_selValid_741) || _zz_s1_outputPayload_selValid_742) || _zz_s1_outputPayload_selValid_743);
  assign _zz_s1_outputPayload_sel_23_4 = (((((((((((((((_zz_s1_outputPayload_selValid_728 || _zz_s1_outputPayload_selValid_729) || _zz_s1_outputPayload_selValid_730) || _zz_s1_outputPayload_selValid_731) || _zz_s1_outputPayload_selValid_732) || _zz_s1_outputPayload_selValid_733) || _zz_s1_outputPayload_selValid_734) || _zz_s1_outputPayload_selValid_735) || _zz_s1_outputPayload_selValid_736) || _zz_s1_outputPayload_selValid_737) || _zz_s1_outputPayload_selValid_738) || _zz_s1_outputPayload_selValid_739) || _zz_s1_outputPayload_selValid_740) || _zz_s1_outputPayload_selValid_741) || _zz_s1_outputPayload_selValid_742) || _zz_s1_outputPayload_selValid_743);
  assign s1_outputPayload_sel_23 = {_zz_s1_outputPayload_sel_23_4,{_zz_s1_outputPayload_sel_23_3,{_zz_s1_outputPayload_sel_23_2,{_zz_s1_outputPayload_sel_23_1,_zz_s1_outputPayload_sel_23}}}};
  assign _zz_s1_outputPayload_selValid_744 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h18));
  assign _zz_s1_outputPayload_selValid_745 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h18));
  assign _zz_s1_outputPayload_selValid_746 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h18));
  assign _zz_s1_outputPayload_selValid_747 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h18));
  assign _zz_s1_outputPayload_selValid_748 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h18));
  assign _zz_s1_outputPayload_selValid_749 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h18));
  assign _zz_s1_outputPayload_selValid_750 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h18));
  assign _zz_s1_outputPayload_selValid_751 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h18));
  assign _zz_s1_outputPayload_selValid_752 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h18));
  assign _zz_s1_outputPayload_selValid_753 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h18));
  assign _zz_s1_outputPayload_selValid_754 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h18));
  assign _zz_s1_outputPayload_selValid_755 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h18));
  assign _zz_s1_outputPayload_selValid_756 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h18));
  assign _zz_s1_outputPayload_selValid_757 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h18));
  assign _zz_s1_outputPayload_selValid_758 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h18));
  assign _zz_s1_outputPayload_selValid_759 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h18));
  assign _zz_s1_outputPayload_selValid_760 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h18));
  assign _zz_s1_outputPayload_selValid_761 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h18));
  assign _zz_s1_outputPayload_selValid_762 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h18));
  assign _zz_s1_outputPayload_selValid_763 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h18));
  assign _zz_s1_outputPayload_selValid_764 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h18));
  assign _zz_s1_outputPayload_selValid_765 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h18));
  assign _zz_s1_outputPayload_selValid_766 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h18));
  assign _zz_s1_outputPayload_selValid_767 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h18));
  assign _zz_s1_outputPayload_selValid_768 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h18));
  assign _zz_s1_outputPayload_selValid_769 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h18));
  assign _zz_s1_outputPayload_selValid_770 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h18));
  assign _zz_s1_outputPayload_selValid_771 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h18));
  assign _zz_s1_outputPayload_selValid_772 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h18));
  assign _zz_s1_outputPayload_selValid_773 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h18));
  assign _zz_s1_outputPayload_selValid_774 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h18));
  assign _zz_s1_outputPayload_sel_24 = (((((((((((((((_zz_s1_outputPayload_selValid_744 || _zz_s1_outputPayload_selValid_746) || _zz_s1_outputPayload_selValid_748) || _zz_s1_outputPayload_selValid_750) || _zz_s1_outputPayload_selValid_752) || _zz_s1_outputPayload_selValid_754) || _zz_s1_outputPayload_selValid_756) || _zz_s1_outputPayload_selValid_758) || _zz_s1_outputPayload_selValid_760) || _zz_s1_outputPayload_selValid_762) || _zz_s1_outputPayload_selValid_764) || _zz_s1_outputPayload_selValid_766) || _zz_s1_outputPayload_selValid_768) || _zz_s1_outputPayload_selValid_770) || _zz_s1_outputPayload_selValid_772) || _zz_s1_outputPayload_selValid_774);
  assign _zz_s1_outputPayload_sel_24_1 = (((((((((((((((_zz_s1_outputPayload_selValid_745 || _zz_s1_outputPayload_selValid_746) || _zz_s1_outputPayload_selValid_749) || _zz_s1_outputPayload_selValid_750) || _zz_s1_outputPayload_selValid_753) || _zz_s1_outputPayload_selValid_754) || _zz_s1_outputPayload_selValid_757) || _zz_s1_outputPayload_selValid_758) || _zz_s1_outputPayload_selValid_761) || _zz_s1_outputPayload_selValid_762) || _zz_s1_outputPayload_selValid_765) || _zz_s1_outputPayload_selValid_766) || _zz_s1_outputPayload_selValid_769) || _zz_s1_outputPayload_selValid_770) || _zz_s1_outputPayload_selValid_773) || _zz_s1_outputPayload_selValid_774);
  assign _zz_s1_outputPayload_sel_24_2 = (((((((((((((((_zz_s1_outputPayload_selValid_747 || _zz_s1_outputPayload_selValid_748) || _zz_s1_outputPayload_selValid_749) || _zz_s1_outputPayload_selValid_750) || _zz_s1_outputPayload_selValid_755) || _zz_s1_outputPayload_selValid_756) || _zz_s1_outputPayload_selValid_757) || _zz_s1_outputPayload_selValid_758) || _zz_s1_outputPayload_selValid_763) || _zz_s1_outputPayload_selValid_764) || _zz_s1_outputPayload_selValid_765) || _zz_s1_outputPayload_selValid_766) || _zz_s1_outputPayload_selValid_771) || _zz_s1_outputPayload_selValid_772) || _zz_s1_outputPayload_selValid_773) || _zz_s1_outputPayload_selValid_774);
  assign _zz_s1_outputPayload_sel_24_3 = (((((((((((((((_zz_s1_outputPayload_selValid_751 || _zz_s1_outputPayload_selValid_752) || _zz_s1_outputPayload_selValid_753) || _zz_s1_outputPayload_selValid_754) || _zz_s1_outputPayload_selValid_755) || _zz_s1_outputPayload_selValid_756) || _zz_s1_outputPayload_selValid_757) || _zz_s1_outputPayload_selValid_758) || _zz_s1_outputPayload_selValid_767) || _zz_s1_outputPayload_selValid_768) || _zz_s1_outputPayload_selValid_769) || _zz_s1_outputPayload_selValid_770) || _zz_s1_outputPayload_selValid_771) || _zz_s1_outputPayload_selValid_772) || _zz_s1_outputPayload_selValid_773) || _zz_s1_outputPayload_selValid_774);
  assign _zz_s1_outputPayload_sel_24_4 = (((((((((((((((_zz_s1_outputPayload_selValid_759 || _zz_s1_outputPayload_selValid_760) || _zz_s1_outputPayload_selValid_761) || _zz_s1_outputPayload_selValid_762) || _zz_s1_outputPayload_selValid_763) || _zz_s1_outputPayload_selValid_764) || _zz_s1_outputPayload_selValid_765) || _zz_s1_outputPayload_selValid_766) || _zz_s1_outputPayload_selValid_767) || _zz_s1_outputPayload_selValid_768) || _zz_s1_outputPayload_selValid_769) || _zz_s1_outputPayload_selValid_770) || _zz_s1_outputPayload_selValid_771) || _zz_s1_outputPayload_selValid_772) || _zz_s1_outputPayload_selValid_773) || _zz_s1_outputPayload_selValid_774);
  assign s1_outputPayload_sel_24 = {_zz_s1_outputPayload_sel_24_4,{_zz_s1_outputPayload_sel_24_3,{_zz_s1_outputPayload_sel_24_2,{_zz_s1_outputPayload_sel_24_1,_zz_s1_outputPayload_sel_24}}}};
  assign _zz_s1_outputPayload_selValid_775 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h19));
  assign _zz_s1_outputPayload_selValid_776 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h19));
  assign _zz_s1_outputPayload_selValid_777 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h19));
  assign _zz_s1_outputPayload_selValid_778 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h19));
  assign _zz_s1_outputPayload_selValid_779 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h19));
  assign _zz_s1_outputPayload_selValid_780 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h19));
  assign _zz_s1_outputPayload_selValid_781 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h19));
  assign _zz_s1_outputPayload_selValid_782 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h19));
  assign _zz_s1_outputPayload_selValid_783 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h19));
  assign _zz_s1_outputPayload_selValid_784 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h19));
  assign _zz_s1_outputPayload_selValid_785 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h19));
  assign _zz_s1_outputPayload_selValid_786 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h19));
  assign _zz_s1_outputPayload_selValid_787 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h19));
  assign _zz_s1_outputPayload_selValid_788 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h19));
  assign _zz_s1_outputPayload_selValid_789 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h19));
  assign _zz_s1_outputPayload_selValid_790 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h19));
  assign _zz_s1_outputPayload_selValid_791 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h19));
  assign _zz_s1_outputPayload_selValid_792 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h19));
  assign _zz_s1_outputPayload_selValid_793 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h19));
  assign _zz_s1_outputPayload_selValid_794 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h19));
  assign _zz_s1_outputPayload_selValid_795 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h19));
  assign _zz_s1_outputPayload_selValid_796 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h19));
  assign _zz_s1_outputPayload_selValid_797 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h19));
  assign _zz_s1_outputPayload_selValid_798 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h19));
  assign _zz_s1_outputPayload_selValid_799 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h19));
  assign _zz_s1_outputPayload_selValid_800 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h19));
  assign _zz_s1_outputPayload_selValid_801 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h19));
  assign _zz_s1_outputPayload_selValid_802 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h19));
  assign _zz_s1_outputPayload_selValid_803 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h19));
  assign _zz_s1_outputPayload_selValid_804 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h19));
  assign _zz_s1_outputPayload_selValid_805 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h19));
  assign _zz_s1_outputPayload_sel_25 = (((((((((((((((_zz_s1_outputPayload_selValid_775 || _zz_s1_outputPayload_selValid_777) || _zz_s1_outputPayload_selValid_779) || _zz_s1_outputPayload_selValid_781) || _zz_s1_outputPayload_selValid_783) || _zz_s1_outputPayload_selValid_785) || _zz_s1_outputPayload_selValid_787) || _zz_s1_outputPayload_selValid_789) || _zz_s1_outputPayload_selValid_791) || _zz_s1_outputPayload_selValid_793) || _zz_s1_outputPayload_selValid_795) || _zz_s1_outputPayload_selValid_797) || _zz_s1_outputPayload_selValid_799) || _zz_s1_outputPayload_selValid_801) || _zz_s1_outputPayload_selValid_803) || _zz_s1_outputPayload_selValid_805);
  assign _zz_s1_outputPayload_sel_25_1 = (((((((((((((((_zz_s1_outputPayload_selValid_776 || _zz_s1_outputPayload_selValid_777) || _zz_s1_outputPayload_selValid_780) || _zz_s1_outputPayload_selValid_781) || _zz_s1_outputPayload_selValid_784) || _zz_s1_outputPayload_selValid_785) || _zz_s1_outputPayload_selValid_788) || _zz_s1_outputPayload_selValid_789) || _zz_s1_outputPayload_selValid_792) || _zz_s1_outputPayload_selValid_793) || _zz_s1_outputPayload_selValid_796) || _zz_s1_outputPayload_selValid_797) || _zz_s1_outputPayload_selValid_800) || _zz_s1_outputPayload_selValid_801) || _zz_s1_outputPayload_selValid_804) || _zz_s1_outputPayload_selValid_805);
  assign _zz_s1_outputPayload_sel_25_2 = (((((((((((((((_zz_s1_outputPayload_selValid_778 || _zz_s1_outputPayload_selValid_779) || _zz_s1_outputPayload_selValid_780) || _zz_s1_outputPayload_selValid_781) || _zz_s1_outputPayload_selValid_786) || _zz_s1_outputPayload_selValid_787) || _zz_s1_outputPayload_selValid_788) || _zz_s1_outputPayload_selValid_789) || _zz_s1_outputPayload_selValid_794) || _zz_s1_outputPayload_selValid_795) || _zz_s1_outputPayload_selValid_796) || _zz_s1_outputPayload_selValid_797) || _zz_s1_outputPayload_selValid_802) || _zz_s1_outputPayload_selValid_803) || _zz_s1_outputPayload_selValid_804) || _zz_s1_outputPayload_selValid_805);
  assign _zz_s1_outputPayload_sel_25_3 = (((((((((((((((_zz_s1_outputPayload_selValid_782 || _zz_s1_outputPayload_selValid_783) || _zz_s1_outputPayload_selValid_784) || _zz_s1_outputPayload_selValid_785) || _zz_s1_outputPayload_selValid_786) || _zz_s1_outputPayload_selValid_787) || _zz_s1_outputPayload_selValid_788) || _zz_s1_outputPayload_selValid_789) || _zz_s1_outputPayload_selValid_798) || _zz_s1_outputPayload_selValid_799) || _zz_s1_outputPayload_selValid_800) || _zz_s1_outputPayload_selValid_801) || _zz_s1_outputPayload_selValid_802) || _zz_s1_outputPayload_selValid_803) || _zz_s1_outputPayload_selValid_804) || _zz_s1_outputPayload_selValid_805);
  assign _zz_s1_outputPayload_sel_25_4 = (((((((((((((((_zz_s1_outputPayload_selValid_790 || _zz_s1_outputPayload_selValid_791) || _zz_s1_outputPayload_selValid_792) || _zz_s1_outputPayload_selValid_793) || _zz_s1_outputPayload_selValid_794) || _zz_s1_outputPayload_selValid_795) || _zz_s1_outputPayload_selValid_796) || _zz_s1_outputPayload_selValid_797) || _zz_s1_outputPayload_selValid_798) || _zz_s1_outputPayload_selValid_799) || _zz_s1_outputPayload_selValid_800) || _zz_s1_outputPayload_selValid_801) || _zz_s1_outputPayload_selValid_802) || _zz_s1_outputPayload_selValid_803) || _zz_s1_outputPayload_selValid_804) || _zz_s1_outputPayload_selValid_805);
  assign s1_outputPayload_sel_25 = {_zz_s1_outputPayload_sel_25_4,{_zz_s1_outputPayload_sel_25_3,{_zz_s1_outputPayload_sel_25_2,{_zz_s1_outputPayload_sel_25_1,_zz_s1_outputPayload_sel_25}}}};
  assign _zz_s1_outputPayload_selValid_806 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_807 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_808 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_809 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_810 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_811 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_812 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_813 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_814 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_815 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_816 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_817 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_818 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_819 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_820 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_821 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_822 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_823 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_824 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_825 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_826 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_827 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_828 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_829 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_830 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_831 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_832 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_833 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_834 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_835 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h1a));
  assign _zz_s1_outputPayload_selValid_836 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h1a));
  assign _zz_s1_outputPayload_sel_26 = (((((((((((((((_zz_s1_outputPayload_selValid_806 || _zz_s1_outputPayload_selValid_808) || _zz_s1_outputPayload_selValid_810) || _zz_s1_outputPayload_selValid_812) || _zz_s1_outputPayload_selValid_814) || _zz_s1_outputPayload_selValid_816) || _zz_s1_outputPayload_selValid_818) || _zz_s1_outputPayload_selValid_820) || _zz_s1_outputPayload_selValid_822) || _zz_s1_outputPayload_selValid_824) || _zz_s1_outputPayload_selValid_826) || _zz_s1_outputPayload_selValid_828) || _zz_s1_outputPayload_selValid_830) || _zz_s1_outputPayload_selValid_832) || _zz_s1_outputPayload_selValid_834) || _zz_s1_outputPayload_selValid_836);
  assign _zz_s1_outputPayload_sel_26_1 = (((((((((((((((_zz_s1_outputPayload_selValid_807 || _zz_s1_outputPayload_selValid_808) || _zz_s1_outputPayload_selValid_811) || _zz_s1_outputPayload_selValid_812) || _zz_s1_outputPayload_selValid_815) || _zz_s1_outputPayload_selValid_816) || _zz_s1_outputPayload_selValid_819) || _zz_s1_outputPayload_selValid_820) || _zz_s1_outputPayload_selValid_823) || _zz_s1_outputPayload_selValid_824) || _zz_s1_outputPayload_selValid_827) || _zz_s1_outputPayload_selValid_828) || _zz_s1_outputPayload_selValid_831) || _zz_s1_outputPayload_selValid_832) || _zz_s1_outputPayload_selValid_835) || _zz_s1_outputPayload_selValid_836);
  assign _zz_s1_outputPayload_sel_26_2 = (((((((((((((((_zz_s1_outputPayload_selValid_809 || _zz_s1_outputPayload_selValid_810) || _zz_s1_outputPayload_selValid_811) || _zz_s1_outputPayload_selValid_812) || _zz_s1_outputPayload_selValid_817) || _zz_s1_outputPayload_selValid_818) || _zz_s1_outputPayload_selValid_819) || _zz_s1_outputPayload_selValid_820) || _zz_s1_outputPayload_selValid_825) || _zz_s1_outputPayload_selValid_826) || _zz_s1_outputPayload_selValid_827) || _zz_s1_outputPayload_selValid_828) || _zz_s1_outputPayload_selValid_833) || _zz_s1_outputPayload_selValid_834) || _zz_s1_outputPayload_selValid_835) || _zz_s1_outputPayload_selValid_836);
  assign _zz_s1_outputPayload_sel_26_3 = (((((((((((((((_zz_s1_outputPayload_selValid_813 || _zz_s1_outputPayload_selValid_814) || _zz_s1_outputPayload_selValid_815) || _zz_s1_outputPayload_selValid_816) || _zz_s1_outputPayload_selValid_817) || _zz_s1_outputPayload_selValid_818) || _zz_s1_outputPayload_selValid_819) || _zz_s1_outputPayload_selValid_820) || _zz_s1_outputPayload_selValid_829) || _zz_s1_outputPayload_selValid_830) || _zz_s1_outputPayload_selValid_831) || _zz_s1_outputPayload_selValid_832) || _zz_s1_outputPayload_selValid_833) || _zz_s1_outputPayload_selValid_834) || _zz_s1_outputPayload_selValid_835) || _zz_s1_outputPayload_selValid_836);
  assign _zz_s1_outputPayload_sel_26_4 = (((((((((((((((_zz_s1_outputPayload_selValid_821 || _zz_s1_outputPayload_selValid_822) || _zz_s1_outputPayload_selValid_823) || _zz_s1_outputPayload_selValid_824) || _zz_s1_outputPayload_selValid_825) || _zz_s1_outputPayload_selValid_826) || _zz_s1_outputPayload_selValid_827) || _zz_s1_outputPayload_selValid_828) || _zz_s1_outputPayload_selValid_829) || _zz_s1_outputPayload_selValid_830) || _zz_s1_outputPayload_selValid_831) || _zz_s1_outputPayload_selValid_832) || _zz_s1_outputPayload_selValid_833) || _zz_s1_outputPayload_selValid_834) || _zz_s1_outputPayload_selValid_835) || _zz_s1_outputPayload_selValid_836);
  assign s1_outputPayload_sel_26 = {_zz_s1_outputPayload_sel_26_4,{_zz_s1_outputPayload_sel_26_3,{_zz_s1_outputPayload_sel_26_2,{_zz_s1_outputPayload_sel_26_1,_zz_s1_outputPayload_sel_26}}}};
  assign _zz_s1_outputPayload_selValid_837 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_838 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_839 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_840 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_841 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_842 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_843 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_844 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_845 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_846 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_847 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_848 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_849 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_850 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_851 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_852 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_853 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_854 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_855 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_856 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_857 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_858 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_859 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_860 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_861 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_862 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_863 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_864 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_865 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_866 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h1b));
  assign _zz_s1_outputPayload_selValid_867 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h1b));
  assign _zz_s1_outputPayload_sel_27 = (((((((((((((((_zz_s1_outputPayload_selValid_837 || _zz_s1_outputPayload_selValid_839) || _zz_s1_outputPayload_selValid_841) || _zz_s1_outputPayload_selValid_843) || _zz_s1_outputPayload_selValid_845) || _zz_s1_outputPayload_selValid_847) || _zz_s1_outputPayload_selValid_849) || _zz_s1_outputPayload_selValid_851) || _zz_s1_outputPayload_selValid_853) || _zz_s1_outputPayload_selValid_855) || _zz_s1_outputPayload_selValid_857) || _zz_s1_outputPayload_selValid_859) || _zz_s1_outputPayload_selValid_861) || _zz_s1_outputPayload_selValid_863) || _zz_s1_outputPayload_selValid_865) || _zz_s1_outputPayload_selValid_867);
  assign _zz_s1_outputPayload_sel_27_1 = (((((((((((((((_zz_s1_outputPayload_selValid_838 || _zz_s1_outputPayload_selValid_839) || _zz_s1_outputPayload_selValid_842) || _zz_s1_outputPayload_selValid_843) || _zz_s1_outputPayload_selValid_846) || _zz_s1_outputPayload_selValid_847) || _zz_s1_outputPayload_selValid_850) || _zz_s1_outputPayload_selValid_851) || _zz_s1_outputPayload_selValid_854) || _zz_s1_outputPayload_selValid_855) || _zz_s1_outputPayload_selValid_858) || _zz_s1_outputPayload_selValid_859) || _zz_s1_outputPayload_selValid_862) || _zz_s1_outputPayload_selValid_863) || _zz_s1_outputPayload_selValid_866) || _zz_s1_outputPayload_selValid_867);
  assign _zz_s1_outputPayload_sel_27_2 = (((((((((((((((_zz_s1_outputPayload_selValid_840 || _zz_s1_outputPayload_selValid_841) || _zz_s1_outputPayload_selValid_842) || _zz_s1_outputPayload_selValid_843) || _zz_s1_outputPayload_selValid_848) || _zz_s1_outputPayload_selValid_849) || _zz_s1_outputPayload_selValid_850) || _zz_s1_outputPayload_selValid_851) || _zz_s1_outputPayload_selValid_856) || _zz_s1_outputPayload_selValid_857) || _zz_s1_outputPayload_selValid_858) || _zz_s1_outputPayload_selValid_859) || _zz_s1_outputPayload_selValid_864) || _zz_s1_outputPayload_selValid_865) || _zz_s1_outputPayload_selValid_866) || _zz_s1_outputPayload_selValid_867);
  assign _zz_s1_outputPayload_sel_27_3 = (((((((((((((((_zz_s1_outputPayload_selValid_844 || _zz_s1_outputPayload_selValid_845) || _zz_s1_outputPayload_selValid_846) || _zz_s1_outputPayload_selValid_847) || _zz_s1_outputPayload_selValid_848) || _zz_s1_outputPayload_selValid_849) || _zz_s1_outputPayload_selValid_850) || _zz_s1_outputPayload_selValid_851) || _zz_s1_outputPayload_selValid_860) || _zz_s1_outputPayload_selValid_861) || _zz_s1_outputPayload_selValid_862) || _zz_s1_outputPayload_selValid_863) || _zz_s1_outputPayload_selValid_864) || _zz_s1_outputPayload_selValid_865) || _zz_s1_outputPayload_selValid_866) || _zz_s1_outputPayload_selValid_867);
  assign _zz_s1_outputPayload_sel_27_4 = (((((((((((((((_zz_s1_outputPayload_selValid_852 || _zz_s1_outputPayload_selValid_853) || _zz_s1_outputPayload_selValid_854) || _zz_s1_outputPayload_selValid_855) || _zz_s1_outputPayload_selValid_856) || _zz_s1_outputPayload_selValid_857) || _zz_s1_outputPayload_selValid_858) || _zz_s1_outputPayload_selValid_859) || _zz_s1_outputPayload_selValid_860) || _zz_s1_outputPayload_selValid_861) || _zz_s1_outputPayload_selValid_862) || _zz_s1_outputPayload_selValid_863) || _zz_s1_outputPayload_selValid_864) || _zz_s1_outputPayload_selValid_865) || _zz_s1_outputPayload_selValid_866) || _zz_s1_outputPayload_selValid_867);
  assign s1_outputPayload_sel_27 = {_zz_s1_outputPayload_sel_27_4,{_zz_s1_outputPayload_sel_27_3,{_zz_s1_outputPayload_sel_27_2,{_zz_s1_outputPayload_sel_27_1,_zz_s1_outputPayload_sel_27}}}};
  assign _zz_s1_outputPayload_selValid_868 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_869 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_870 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_871 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_872 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_873 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_874 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_875 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_876 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_877 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_878 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_879 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_880 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_881 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_882 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_883 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_884 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_885 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_886 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_887 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_888 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_889 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_890 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_891 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_892 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_893 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_894 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_895 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_896 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_897 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h1c));
  assign _zz_s1_outputPayload_selValid_898 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h1c));
  assign _zz_s1_outputPayload_sel_28 = (((((((((((((((_zz_s1_outputPayload_selValid_868 || _zz_s1_outputPayload_selValid_870) || _zz_s1_outputPayload_selValid_872) || _zz_s1_outputPayload_selValid_874) || _zz_s1_outputPayload_selValid_876) || _zz_s1_outputPayload_selValid_878) || _zz_s1_outputPayload_selValid_880) || _zz_s1_outputPayload_selValid_882) || _zz_s1_outputPayload_selValid_884) || _zz_s1_outputPayload_selValid_886) || _zz_s1_outputPayload_selValid_888) || _zz_s1_outputPayload_selValid_890) || _zz_s1_outputPayload_selValid_892) || _zz_s1_outputPayload_selValid_894) || _zz_s1_outputPayload_selValid_896) || _zz_s1_outputPayload_selValid_898);
  assign _zz_s1_outputPayload_sel_28_1 = (((((((((((((((_zz_s1_outputPayload_selValid_869 || _zz_s1_outputPayload_selValid_870) || _zz_s1_outputPayload_selValid_873) || _zz_s1_outputPayload_selValid_874) || _zz_s1_outputPayload_selValid_877) || _zz_s1_outputPayload_selValid_878) || _zz_s1_outputPayload_selValid_881) || _zz_s1_outputPayload_selValid_882) || _zz_s1_outputPayload_selValid_885) || _zz_s1_outputPayload_selValid_886) || _zz_s1_outputPayload_selValid_889) || _zz_s1_outputPayload_selValid_890) || _zz_s1_outputPayload_selValid_893) || _zz_s1_outputPayload_selValid_894) || _zz_s1_outputPayload_selValid_897) || _zz_s1_outputPayload_selValid_898);
  assign _zz_s1_outputPayload_sel_28_2 = (((((((((((((((_zz_s1_outputPayload_selValid_871 || _zz_s1_outputPayload_selValid_872) || _zz_s1_outputPayload_selValid_873) || _zz_s1_outputPayload_selValid_874) || _zz_s1_outputPayload_selValid_879) || _zz_s1_outputPayload_selValid_880) || _zz_s1_outputPayload_selValid_881) || _zz_s1_outputPayload_selValid_882) || _zz_s1_outputPayload_selValid_887) || _zz_s1_outputPayload_selValid_888) || _zz_s1_outputPayload_selValid_889) || _zz_s1_outputPayload_selValid_890) || _zz_s1_outputPayload_selValid_895) || _zz_s1_outputPayload_selValid_896) || _zz_s1_outputPayload_selValid_897) || _zz_s1_outputPayload_selValid_898);
  assign _zz_s1_outputPayload_sel_28_3 = (((((((((((((((_zz_s1_outputPayload_selValid_875 || _zz_s1_outputPayload_selValid_876) || _zz_s1_outputPayload_selValid_877) || _zz_s1_outputPayload_selValid_878) || _zz_s1_outputPayload_selValid_879) || _zz_s1_outputPayload_selValid_880) || _zz_s1_outputPayload_selValid_881) || _zz_s1_outputPayload_selValid_882) || _zz_s1_outputPayload_selValid_891) || _zz_s1_outputPayload_selValid_892) || _zz_s1_outputPayload_selValid_893) || _zz_s1_outputPayload_selValid_894) || _zz_s1_outputPayload_selValid_895) || _zz_s1_outputPayload_selValid_896) || _zz_s1_outputPayload_selValid_897) || _zz_s1_outputPayload_selValid_898);
  assign _zz_s1_outputPayload_sel_28_4 = (((((((((((((((_zz_s1_outputPayload_selValid_883 || _zz_s1_outputPayload_selValid_884) || _zz_s1_outputPayload_selValid_885) || _zz_s1_outputPayload_selValid_886) || _zz_s1_outputPayload_selValid_887) || _zz_s1_outputPayload_selValid_888) || _zz_s1_outputPayload_selValid_889) || _zz_s1_outputPayload_selValid_890) || _zz_s1_outputPayload_selValid_891) || _zz_s1_outputPayload_selValid_892) || _zz_s1_outputPayload_selValid_893) || _zz_s1_outputPayload_selValid_894) || _zz_s1_outputPayload_selValid_895) || _zz_s1_outputPayload_selValid_896) || _zz_s1_outputPayload_selValid_897) || _zz_s1_outputPayload_selValid_898);
  assign s1_outputPayload_sel_28 = {_zz_s1_outputPayload_sel_28_4,{_zz_s1_outputPayload_sel_28_3,{_zz_s1_outputPayload_sel_28_2,{_zz_s1_outputPayload_sel_28_1,_zz_s1_outputPayload_sel_28}}}};
  assign _zz_s1_outputPayload_selValid_899 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_900 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_901 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_902 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_903 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_904 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_905 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_906 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_907 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_908 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_909 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_910 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_911 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_912 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_913 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_914 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_915 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_916 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_917 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_918 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_919 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_920 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_921 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_922 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_923 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_924 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_925 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_926 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_927 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_928 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h1d));
  assign _zz_s1_outputPayload_selValid_929 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h1d));
  assign _zz_s1_outputPayload_sel_29 = (((((((((((((((_zz_s1_outputPayload_selValid_899 || _zz_s1_outputPayload_selValid_901) || _zz_s1_outputPayload_selValid_903) || _zz_s1_outputPayload_selValid_905) || _zz_s1_outputPayload_selValid_907) || _zz_s1_outputPayload_selValid_909) || _zz_s1_outputPayload_selValid_911) || _zz_s1_outputPayload_selValid_913) || _zz_s1_outputPayload_selValid_915) || _zz_s1_outputPayload_selValid_917) || _zz_s1_outputPayload_selValid_919) || _zz_s1_outputPayload_selValid_921) || _zz_s1_outputPayload_selValid_923) || _zz_s1_outputPayload_selValid_925) || _zz_s1_outputPayload_selValid_927) || _zz_s1_outputPayload_selValid_929);
  assign _zz_s1_outputPayload_sel_29_1 = (((((((((((((((_zz_s1_outputPayload_selValid_900 || _zz_s1_outputPayload_selValid_901) || _zz_s1_outputPayload_selValid_904) || _zz_s1_outputPayload_selValid_905) || _zz_s1_outputPayload_selValid_908) || _zz_s1_outputPayload_selValid_909) || _zz_s1_outputPayload_selValid_912) || _zz_s1_outputPayload_selValid_913) || _zz_s1_outputPayload_selValid_916) || _zz_s1_outputPayload_selValid_917) || _zz_s1_outputPayload_selValid_920) || _zz_s1_outputPayload_selValid_921) || _zz_s1_outputPayload_selValid_924) || _zz_s1_outputPayload_selValid_925) || _zz_s1_outputPayload_selValid_928) || _zz_s1_outputPayload_selValid_929);
  assign _zz_s1_outputPayload_sel_29_2 = (((((((((((((((_zz_s1_outputPayload_selValid_902 || _zz_s1_outputPayload_selValid_903) || _zz_s1_outputPayload_selValid_904) || _zz_s1_outputPayload_selValid_905) || _zz_s1_outputPayload_selValid_910) || _zz_s1_outputPayload_selValid_911) || _zz_s1_outputPayload_selValid_912) || _zz_s1_outputPayload_selValid_913) || _zz_s1_outputPayload_selValid_918) || _zz_s1_outputPayload_selValid_919) || _zz_s1_outputPayload_selValid_920) || _zz_s1_outputPayload_selValid_921) || _zz_s1_outputPayload_selValid_926) || _zz_s1_outputPayload_selValid_927) || _zz_s1_outputPayload_selValid_928) || _zz_s1_outputPayload_selValid_929);
  assign _zz_s1_outputPayload_sel_29_3 = (((((((((((((((_zz_s1_outputPayload_selValid_906 || _zz_s1_outputPayload_selValid_907) || _zz_s1_outputPayload_selValid_908) || _zz_s1_outputPayload_selValid_909) || _zz_s1_outputPayload_selValid_910) || _zz_s1_outputPayload_selValid_911) || _zz_s1_outputPayload_selValid_912) || _zz_s1_outputPayload_selValid_913) || _zz_s1_outputPayload_selValid_922) || _zz_s1_outputPayload_selValid_923) || _zz_s1_outputPayload_selValid_924) || _zz_s1_outputPayload_selValid_925) || _zz_s1_outputPayload_selValid_926) || _zz_s1_outputPayload_selValid_927) || _zz_s1_outputPayload_selValid_928) || _zz_s1_outputPayload_selValid_929);
  assign _zz_s1_outputPayload_sel_29_4 = (((((((((((((((_zz_s1_outputPayload_selValid_914 || _zz_s1_outputPayload_selValid_915) || _zz_s1_outputPayload_selValid_916) || _zz_s1_outputPayload_selValid_917) || _zz_s1_outputPayload_selValid_918) || _zz_s1_outputPayload_selValid_919) || _zz_s1_outputPayload_selValid_920) || _zz_s1_outputPayload_selValid_921) || _zz_s1_outputPayload_selValid_922) || _zz_s1_outputPayload_selValid_923) || _zz_s1_outputPayload_selValid_924) || _zz_s1_outputPayload_selValid_925) || _zz_s1_outputPayload_selValid_926) || _zz_s1_outputPayload_selValid_927) || _zz_s1_outputPayload_selValid_928) || _zz_s1_outputPayload_selValid_929);
  assign s1_outputPayload_sel_29 = {_zz_s1_outputPayload_sel_29_4,{_zz_s1_outputPayload_sel_29_3,{_zz_s1_outputPayload_sel_29_2,{_zz_s1_outputPayload_sel_29_1,_zz_s1_outputPayload_sel_29}}}};
  assign _zz_s1_outputPayload_selValid_930 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_931 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_932 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_933 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_934 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_935 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_936 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_937 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_938 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_939 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_940 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_941 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_942 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_943 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_944 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_945 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_946 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_947 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_948 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_949 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_950 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_951 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_952 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_953 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_954 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_955 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_956 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_957 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_958 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_959 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h1e));
  assign _zz_s1_outputPayload_selValid_960 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h1e));
  assign _zz_s1_outputPayload_sel_30 = (((((((((((((((_zz_s1_outputPayload_selValid_930 || _zz_s1_outputPayload_selValid_932) || _zz_s1_outputPayload_selValid_934) || _zz_s1_outputPayload_selValid_936) || _zz_s1_outputPayload_selValid_938) || _zz_s1_outputPayload_selValid_940) || _zz_s1_outputPayload_selValid_942) || _zz_s1_outputPayload_selValid_944) || _zz_s1_outputPayload_selValid_946) || _zz_s1_outputPayload_selValid_948) || _zz_s1_outputPayload_selValid_950) || _zz_s1_outputPayload_selValid_952) || _zz_s1_outputPayload_selValid_954) || _zz_s1_outputPayload_selValid_956) || _zz_s1_outputPayload_selValid_958) || _zz_s1_outputPayload_selValid_960);
  assign _zz_s1_outputPayload_sel_30_1 = (((((((((((((((_zz_s1_outputPayload_selValid_931 || _zz_s1_outputPayload_selValid_932) || _zz_s1_outputPayload_selValid_935) || _zz_s1_outputPayload_selValid_936) || _zz_s1_outputPayload_selValid_939) || _zz_s1_outputPayload_selValid_940) || _zz_s1_outputPayload_selValid_943) || _zz_s1_outputPayload_selValid_944) || _zz_s1_outputPayload_selValid_947) || _zz_s1_outputPayload_selValid_948) || _zz_s1_outputPayload_selValid_951) || _zz_s1_outputPayload_selValid_952) || _zz_s1_outputPayload_selValid_955) || _zz_s1_outputPayload_selValid_956) || _zz_s1_outputPayload_selValid_959) || _zz_s1_outputPayload_selValid_960);
  assign _zz_s1_outputPayload_sel_30_2 = (((((((((((((((_zz_s1_outputPayload_selValid_933 || _zz_s1_outputPayload_selValid_934) || _zz_s1_outputPayload_selValid_935) || _zz_s1_outputPayload_selValid_936) || _zz_s1_outputPayload_selValid_941) || _zz_s1_outputPayload_selValid_942) || _zz_s1_outputPayload_selValid_943) || _zz_s1_outputPayload_selValid_944) || _zz_s1_outputPayload_selValid_949) || _zz_s1_outputPayload_selValid_950) || _zz_s1_outputPayload_selValid_951) || _zz_s1_outputPayload_selValid_952) || _zz_s1_outputPayload_selValid_957) || _zz_s1_outputPayload_selValid_958) || _zz_s1_outputPayload_selValid_959) || _zz_s1_outputPayload_selValid_960);
  assign _zz_s1_outputPayload_sel_30_3 = (((((((((((((((_zz_s1_outputPayload_selValid_937 || _zz_s1_outputPayload_selValid_938) || _zz_s1_outputPayload_selValid_939) || _zz_s1_outputPayload_selValid_940) || _zz_s1_outputPayload_selValid_941) || _zz_s1_outputPayload_selValid_942) || _zz_s1_outputPayload_selValid_943) || _zz_s1_outputPayload_selValid_944) || _zz_s1_outputPayload_selValid_953) || _zz_s1_outputPayload_selValid_954) || _zz_s1_outputPayload_selValid_955) || _zz_s1_outputPayload_selValid_956) || _zz_s1_outputPayload_selValid_957) || _zz_s1_outputPayload_selValid_958) || _zz_s1_outputPayload_selValid_959) || _zz_s1_outputPayload_selValid_960);
  assign _zz_s1_outputPayload_sel_30_4 = (((((((((((((((_zz_s1_outputPayload_selValid_945 || _zz_s1_outputPayload_selValid_946) || _zz_s1_outputPayload_selValid_947) || _zz_s1_outputPayload_selValid_948) || _zz_s1_outputPayload_selValid_949) || _zz_s1_outputPayload_selValid_950) || _zz_s1_outputPayload_selValid_951) || _zz_s1_outputPayload_selValid_952) || _zz_s1_outputPayload_selValid_953) || _zz_s1_outputPayload_selValid_954) || _zz_s1_outputPayload_selValid_955) || _zz_s1_outputPayload_selValid_956) || _zz_s1_outputPayload_selValid_957) || _zz_s1_outputPayload_selValid_958) || _zz_s1_outputPayload_selValid_959) || _zz_s1_outputPayload_selValid_960);
  assign s1_outputPayload_sel_30 = {_zz_s1_outputPayload_sel_30_4,{_zz_s1_outputPayload_sel_30_3,{_zz_s1_outputPayload_sel_30_2,{_zz_s1_outputPayload_sel_30_1,_zz_s1_outputPayload_sel_30}}}};
  assign _zz_s1_outputPayload_selValid_961 = (s1_input_payload_cmd_mask[1] && (s1_inputIndexes_1 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_962 = (s1_input_payload_cmd_mask[2] && (s1_inputIndexes_2 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_963 = (s1_input_payload_cmd_mask[3] && (s1_inputIndexes_3 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_964 = (s1_input_payload_cmd_mask[4] && (s1_inputIndexes_4 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_965 = (s1_input_payload_cmd_mask[5] && (s1_inputIndexes_5 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_966 = (s1_input_payload_cmd_mask[6] && (s1_inputIndexes_6 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_967 = (s1_input_payload_cmd_mask[7] && (s1_inputIndexes_7 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_968 = (s1_input_payload_cmd_mask[8] && (s1_inputIndexes_8 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_969 = (s1_input_payload_cmd_mask[9] && (s1_inputIndexes_9 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_970 = (s1_input_payload_cmd_mask[10] && (s1_inputIndexes_10 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_971 = (s1_input_payload_cmd_mask[11] && (s1_inputIndexes_11 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_972 = (s1_input_payload_cmd_mask[12] && (s1_inputIndexes_12 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_973 = (s1_input_payload_cmd_mask[13] && (s1_inputIndexes_13 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_974 = (s1_input_payload_cmd_mask[14] && (s1_inputIndexes_14 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_975 = (s1_input_payload_cmd_mask[15] && (s1_inputIndexes_15 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_976 = (s1_input_payload_cmd_mask[16] && (s1_inputIndexes_16 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_977 = (s1_input_payload_cmd_mask[17] && (s1_inputIndexes_17 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_978 = (s1_input_payload_cmd_mask[18] && (s1_inputIndexes_18 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_979 = (s1_input_payload_cmd_mask[19] && (s1_inputIndexes_19 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_980 = (s1_input_payload_cmd_mask[20] && (s1_inputIndexes_20 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_981 = (s1_input_payload_cmd_mask[21] && (s1_inputIndexes_21 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_982 = (s1_input_payload_cmd_mask[22] && (s1_inputIndexes_22 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_983 = (s1_input_payload_cmd_mask[23] && (s1_inputIndexes_23 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_984 = (s1_input_payload_cmd_mask[24] && (s1_inputIndexes_24 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_985 = (s1_input_payload_cmd_mask[25] && (s1_inputIndexes_25 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_986 = (s1_input_payload_cmd_mask[26] && (s1_inputIndexes_26 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_987 = (s1_input_payload_cmd_mask[27] && (s1_inputIndexes_27 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_988 = (s1_input_payload_cmd_mask[28] && (s1_inputIndexes_28 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_989 = (s1_input_payload_cmd_mask[29] && (s1_inputIndexes_29 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_990 = (s1_input_payload_cmd_mask[30] && (s1_inputIndexes_30 == 5'h1f));
  assign _zz_s1_outputPayload_selValid_991 = (s1_input_payload_cmd_mask[31] && (s1_inputIndexes_31 == 5'h1f));
  assign _zz_s1_outputPayload_sel_31 = (((((((((((((((_zz_s1_outputPayload_selValid_961 || _zz_s1_outputPayload_selValid_963) || _zz_s1_outputPayload_selValid_965) || _zz_s1_outputPayload_selValid_967) || _zz_s1_outputPayload_selValid_969) || _zz_s1_outputPayload_selValid_971) || _zz_s1_outputPayload_selValid_973) || _zz_s1_outputPayload_selValid_975) || _zz_s1_outputPayload_selValid_977) || _zz_s1_outputPayload_selValid_979) || _zz_s1_outputPayload_selValid_981) || _zz_s1_outputPayload_selValid_983) || _zz_s1_outputPayload_selValid_985) || _zz_s1_outputPayload_selValid_987) || _zz_s1_outputPayload_selValid_989) || _zz_s1_outputPayload_selValid_991);
  assign _zz_s1_outputPayload_sel_31_1 = (((((((((((((((_zz_s1_outputPayload_selValid_962 || _zz_s1_outputPayload_selValid_963) || _zz_s1_outputPayload_selValid_966) || _zz_s1_outputPayload_selValid_967) || _zz_s1_outputPayload_selValid_970) || _zz_s1_outputPayload_selValid_971) || _zz_s1_outputPayload_selValid_974) || _zz_s1_outputPayload_selValid_975) || _zz_s1_outputPayload_selValid_978) || _zz_s1_outputPayload_selValid_979) || _zz_s1_outputPayload_selValid_982) || _zz_s1_outputPayload_selValid_983) || _zz_s1_outputPayload_selValid_986) || _zz_s1_outputPayload_selValid_987) || _zz_s1_outputPayload_selValid_990) || _zz_s1_outputPayload_selValid_991);
  assign _zz_s1_outputPayload_sel_31_2 = (((((((((((((((_zz_s1_outputPayload_selValid_964 || _zz_s1_outputPayload_selValid_965) || _zz_s1_outputPayload_selValid_966) || _zz_s1_outputPayload_selValid_967) || _zz_s1_outputPayload_selValid_972) || _zz_s1_outputPayload_selValid_973) || _zz_s1_outputPayload_selValid_974) || _zz_s1_outputPayload_selValid_975) || _zz_s1_outputPayload_selValid_980) || _zz_s1_outputPayload_selValid_981) || _zz_s1_outputPayload_selValid_982) || _zz_s1_outputPayload_selValid_983) || _zz_s1_outputPayload_selValid_988) || _zz_s1_outputPayload_selValid_989) || _zz_s1_outputPayload_selValid_990) || _zz_s1_outputPayload_selValid_991);
  assign _zz_s1_outputPayload_sel_31_3 = (((((((((((((((_zz_s1_outputPayload_selValid_968 || _zz_s1_outputPayload_selValid_969) || _zz_s1_outputPayload_selValid_970) || _zz_s1_outputPayload_selValid_971) || _zz_s1_outputPayload_selValid_972) || _zz_s1_outputPayload_selValid_973) || _zz_s1_outputPayload_selValid_974) || _zz_s1_outputPayload_selValid_975) || _zz_s1_outputPayload_selValid_984) || _zz_s1_outputPayload_selValid_985) || _zz_s1_outputPayload_selValid_986) || _zz_s1_outputPayload_selValid_987) || _zz_s1_outputPayload_selValid_988) || _zz_s1_outputPayload_selValid_989) || _zz_s1_outputPayload_selValid_990) || _zz_s1_outputPayload_selValid_991);
  assign _zz_s1_outputPayload_sel_31_4 = (((((((((((((((_zz_s1_outputPayload_selValid_976 || _zz_s1_outputPayload_selValid_977) || _zz_s1_outputPayload_selValid_978) || _zz_s1_outputPayload_selValid_979) || _zz_s1_outputPayload_selValid_980) || _zz_s1_outputPayload_selValid_981) || _zz_s1_outputPayload_selValid_982) || _zz_s1_outputPayload_selValid_983) || _zz_s1_outputPayload_selValid_984) || _zz_s1_outputPayload_selValid_985) || _zz_s1_outputPayload_selValid_986) || _zz_s1_outputPayload_selValid_987) || _zz_s1_outputPayload_selValid_988) || _zz_s1_outputPayload_selValid_989) || _zz_s1_outputPayload_selValid_990) || _zz_s1_outputPayload_selValid_991);
  assign s1_outputPayload_sel_31 = {_zz_s1_outputPayload_sel_31_4,{_zz_s1_outputPayload_sel_31_3,{_zz_s1_outputPayload_sel_31_2,{_zz_s1_outputPayload_sel_31_1,_zz_s1_outputPayload_sel_31}}}};
  assign s1_output_valid = s1_input_valid;
  assign s1_input_ready = s1_output_ready;
  assign s1_output_payload_cmd_data = s1_outputPayload_cmd_data;
  assign s1_output_payload_cmd_mask = s1_outputPayload_cmd_mask;
  assign s1_output_payload_index_0 = s1_outputPayload_index_0;
  assign s1_output_payload_index_1 = s1_outputPayload_index_1;
  assign s1_output_payload_index_2 = s1_outputPayload_index_2;
  assign s1_output_payload_index_3 = s1_outputPayload_index_3;
  assign s1_output_payload_index_4 = s1_outputPayload_index_4;
  assign s1_output_payload_index_5 = s1_outputPayload_index_5;
  assign s1_output_payload_index_6 = s1_outputPayload_index_6;
  assign s1_output_payload_index_7 = s1_outputPayload_index_7;
  assign s1_output_payload_index_8 = s1_outputPayload_index_8;
  assign s1_output_payload_index_9 = s1_outputPayload_index_9;
  assign s1_output_payload_index_10 = s1_outputPayload_index_10;
  assign s1_output_payload_index_11 = s1_outputPayload_index_11;
  assign s1_output_payload_index_12 = s1_outputPayload_index_12;
  assign s1_output_payload_index_13 = s1_outputPayload_index_13;
  assign s1_output_payload_index_14 = s1_outputPayload_index_14;
  assign s1_output_payload_index_15 = s1_outputPayload_index_15;
  assign s1_output_payload_index_16 = s1_outputPayload_index_16;
  assign s1_output_payload_index_17 = s1_outputPayload_index_17;
  assign s1_output_payload_index_18 = s1_outputPayload_index_18;
  assign s1_output_payload_index_19 = s1_outputPayload_index_19;
  assign s1_output_payload_index_20 = s1_outputPayload_index_20;
  assign s1_output_payload_index_21 = s1_outputPayload_index_21;
  assign s1_output_payload_index_22 = s1_outputPayload_index_22;
  assign s1_output_payload_index_23 = s1_outputPayload_index_23;
  assign s1_output_payload_index_24 = s1_outputPayload_index_24;
  assign s1_output_payload_index_25 = s1_outputPayload_index_25;
  assign s1_output_payload_index_26 = s1_outputPayload_index_26;
  assign s1_output_payload_index_27 = s1_outputPayload_index_27;
  assign s1_output_payload_index_28 = s1_outputPayload_index_28;
  assign s1_output_payload_index_29 = s1_outputPayload_index_29;
  assign s1_output_payload_index_30 = s1_outputPayload_index_30;
  assign s1_output_payload_index_31 = s1_outputPayload_index_31;
  assign s1_output_payload_last = s1_outputPayload_last;
  assign s1_output_payload_sel_0 = s1_outputPayload_sel_0;
  assign s1_output_payload_sel_1 = s1_outputPayload_sel_1;
  assign s1_output_payload_sel_2 = s1_outputPayload_sel_2;
  assign s1_output_payload_sel_3 = s1_outputPayload_sel_3;
  assign s1_output_payload_sel_4 = s1_outputPayload_sel_4;
  assign s1_output_payload_sel_5 = s1_outputPayload_sel_5;
  assign s1_output_payload_sel_6 = s1_outputPayload_sel_6;
  assign s1_output_payload_sel_7 = s1_outputPayload_sel_7;
  assign s1_output_payload_sel_8 = s1_outputPayload_sel_8;
  assign s1_output_payload_sel_9 = s1_outputPayload_sel_9;
  assign s1_output_payload_sel_10 = s1_outputPayload_sel_10;
  assign s1_output_payload_sel_11 = s1_outputPayload_sel_11;
  assign s1_output_payload_sel_12 = s1_outputPayload_sel_12;
  assign s1_output_payload_sel_13 = s1_outputPayload_sel_13;
  assign s1_output_payload_sel_14 = s1_outputPayload_sel_14;
  assign s1_output_payload_sel_15 = s1_outputPayload_sel_15;
  assign s1_output_payload_sel_16 = s1_outputPayload_sel_16;
  assign s1_output_payload_sel_17 = s1_outputPayload_sel_17;
  assign s1_output_payload_sel_18 = s1_outputPayload_sel_18;
  assign s1_output_payload_sel_19 = s1_outputPayload_sel_19;
  assign s1_output_payload_sel_20 = s1_outputPayload_sel_20;
  assign s1_output_payload_sel_21 = s1_outputPayload_sel_21;
  assign s1_output_payload_sel_22 = s1_outputPayload_sel_22;
  assign s1_output_payload_sel_23 = s1_outputPayload_sel_23;
  assign s1_output_payload_sel_24 = s1_outputPayload_sel_24;
  assign s1_output_payload_sel_25 = s1_outputPayload_sel_25;
  assign s1_output_payload_sel_26 = s1_outputPayload_sel_26;
  assign s1_output_payload_sel_27 = s1_outputPayload_sel_27;
  assign s1_output_payload_sel_28 = s1_outputPayload_sel_28;
  assign s1_output_payload_sel_29 = s1_outputPayload_sel_29;
  assign s1_output_payload_sel_30 = s1_outputPayload_sel_30;
  assign s1_output_payload_sel_31 = s1_outputPayload_sel_31;
  assign s1_output_payload_selValid = s1_outputPayload_selValid;
  always @(*) begin
    s1_output_ready = s2_input_ready;
    if(when_Stream_l375_2) begin
      s1_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_2 = (! s2_input_valid);
  assign s2_input_valid = s1_output_rValid;
  assign s2_input_payload_cmd_data = s1_output_rData_cmd_data;
  assign s2_input_payload_cmd_mask = s1_output_rData_cmd_mask;
  assign s2_input_payload_index_0 = s1_output_rData_index_0;
  assign s2_input_payload_index_1 = s1_output_rData_index_1;
  assign s2_input_payload_index_2 = s1_output_rData_index_2;
  assign s2_input_payload_index_3 = s1_output_rData_index_3;
  assign s2_input_payload_index_4 = s1_output_rData_index_4;
  assign s2_input_payload_index_5 = s1_output_rData_index_5;
  assign s2_input_payload_index_6 = s1_output_rData_index_6;
  assign s2_input_payload_index_7 = s1_output_rData_index_7;
  assign s2_input_payload_index_8 = s1_output_rData_index_8;
  assign s2_input_payload_index_9 = s1_output_rData_index_9;
  assign s2_input_payload_index_10 = s1_output_rData_index_10;
  assign s2_input_payload_index_11 = s1_output_rData_index_11;
  assign s2_input_payload_index_12 = s1_output_rData_index_12;
  assign s2_input_payload_index_13 = s1_output_rData_index_13;
  assign s2_input_payload_index_14 = s1_output_rData_index_14;
  assign s2_input_payload_index_15 = s1_output_rData_index_15;
  assign s2_input_payload_index_16 = s1_output_rData_index_16;
  assign s2_input_payload_index_17 = s1_output_rData_index_17;
  assign s2_input_payload_index_18 = s1_output_rData_index_18;
  assign s2_input_payload_index_19 = s1_output_rData_index_19;
  assign s2_input_payload_index_20 = s1_output_rData_index_20;
  assign s2_input_payload_index_21 = s1_output_rData_index_21;
  assign s2_input_payload_index_22 = s1_output_rData_index_22;
  assign s2_input_payload_index_23 = s1_output_rData_index_23;
  assign s2_input_payload_index_24 = s1_output_rData_index_24;
  assign s2_input_payload_index_25 = s1_output_rData_index_25;
  assign s2_input_payload_index_26 = s1_output_rData_index_26;
  assign s2_input_payload_index_27 = s1_output_rData_index_27;
  assign s2_input_payload_index_28 = s1_output_rData_index_28;
  assign s2_input_payload_index_29 = s1_output_rData_index_29;
  assign s2_input_payload_index_30 = s1_output_rData_index_30;
  assign s2_input_payload_index_31 = s1_output_rData_index_31;
  assign s2_input_payload_last = s1_output_rData_last;
  assign s2_input_payload_sel_0 = s1_output_rData_sel_0;
  assign s2_input_payload_sel_1 = s1_output_rData_sel_1;
  assign s2_input_payload_sel_2 = s1_output_rData_sel_2;
  assign s2_input_payload_sel_3 = s1_output_rData_sel_3;
  assign s2_input_payload_sel_4 = s1_output_rData_sel_4;
  assign s2_input_payload_sel_5 = s1_output_rData_sel_5;
  assign s2_input_payload_sel_6 = s1_output_rData_sel_6;
  assign s2_input_payload_sel_7 = s1_output_rData_sel_7;
  assign s2_input_payload_sel_8 = s1_output_rData_sel_8;
  assign s2_input_payload_sel_9 = s1_output_rData_sel_9;
  assign s2_input_payload_sel_10 = s1_output_rData_sel_10;
  assign s2_input_payload_sel_11 = s1_output_rData_sel_11;
  assign s2_input_payload_sel_12 = s1_output_rData_sel_12;
  assign s2_input_payload_sel_13 = s1_output_rData_sel_13;
  assign s2_input_payload_sel_14 = s1_output_rData_sel_14;
  assign s2_input_payload_sel_15 = s1_output_rData_sel_15;
  assign s2_input_payload_sel_16 = s1_output_rData_sel_16;
  assign s2_input_payload_sel_17 = s1_output_rData_sel_17;
  assign s2_input_payload_sel_18 = s1_output_rData_sel_18;
  assign s2_input_payload_sel_19 = s1_output_rData_sel_19;
  assign s2_input_payload_sel_20 = s1_output_rData_sel_20;
  assign s2_input_payload_sel_21 = s1_output_rData_sel_21;
  assign s2_input_payload_sel_22 = s1_output_rData_sel_22;
  assign s2_input_payload_sel_23 = s1_output_rData_sel_23;
  assign s2_input_payload_sel_24 = s1_output_rData_sel_24;
  assign s2_input_payload_sel_25 = s1_output_rData_sel_25;
  assign s2_input_payload_sel_26 = s1_output_rData_sel_26;
  assign s2_input_payload_sel_27 = s1_output_rData_sel_27;
  assign s2_input_payload_sel_28 = s1_output_rData_sel_28;
  assign s2_input_payload_sel_29 = s1_output_rData_sel_29;
  assign s2_input_payload_sel_30 = s1_output_rData_sel_30;
  assign s2_input_payload_sel_31 = s1_output_rData_sel_31;
  assign s2_input_payload_selValid = s1_output_rData_selValid;
  always @(*) begin
    s2_input_ready = ((! io_output_enough) || io_output_consume);
    if(when_DmaSg_l1464) begin
      s2_input_ready = 1'b0;
    end
  end

  assign when_DmaSg_l1464 = (_zz_when_DmaSg_l1464 < s1_byteCounter);
  assign s2_input_fire = (s2_input_valid && s2_input_ready);
  assign io_output_consumed = s2_input_fire;
  assign s2_inputDataBytes_0 = s2_input_payload_cmd_data[7 : 0];
  assign s2_inputDataBytes_1 = s2_input_payload_cmd_data[15 : 8];
  assign s2_inputDataBytes_2 = s2_input_payload_cmd_data[23 : 16];
  assign s2_inputDataBytes_3 = s2_input_payload_cmd_data[31 : 24];
  assign s2_inputDataBytes_4 = s2_input_payload_cmd_data[39 : 32];
  assign s2_inputDataBytes_5 = s2_input_payload_cmd_data[47 : 40];
  assign s2_inputDataBytes_6 = s2_input_payload_cmd_data[55 : 48];
  assign s2_inputDataBytes_7 = s2_input_payload_cmd_data[63 : 56];
  assign s2_inputDataBytes_8 = s2_input_payload_cmd_data[71 : 64];
  assign s2_inputDataBytes_9 = s2_input_payload_cmd_data[79 : 72];
  assign s2_inputDataBytes_10 = s2_input_payload_cmd_data[87 : 80];
  assign s2_inputDataBytes_11 = s2_input_payload_cmd_data[95 : 88];
  assign s2_inputDataBytes_12 = s2_input_payload_cmd_data[103 : 96];
  assign s2_inputDataBytes_13 = s2_input_payload_cmd_data[111 : 104];
  assign s2_inputDataBytes_14 = s2_input_payload_cmd_data[119 : 112];
  assign s2_inputDataBytes_15 = s2_input_payload_cmd_data[127 : 120];
  assign s2_inputDataBytes_16 = s2_input_payload_cmd_data[135 : 128];
  assign s2_inputDataBytes_17 = s2_input_payload_cmd_data[143 : 136];
  assign s2_inputDataBytes_18 = s2_input_payload_cmd_data[151 : 144];
  assign s2_inputDataBytes_19 = s2_input_payload_cmd_data[159 : 152];
  assign s2_inputDataBytes_20 = s2_input_payload_cmd_data[167 : 160];
  assign s2_inputDataBytes_21 = s2_input_payload_cmd_data[175 : 168];
  assign s2_inputDataBytes_22 = s2_input_payload_cmd_data[183 : 176];
  assign s2_inputDataBytes_23 = s2_input_payload_cmd_data[191 : 184];
  assign s2_inputDataBytes_24 = s2_input_payload_cmd_data[199 : 192];
  assign s2_inputDataBytes_25 = s2_input_payload_cmd_data[207 : 200];
  assign s2_inputDataBytes_26 = s2_input_payload_cmd_data[215 : 208];
  assign s2_inputDataBytes_27 = s2_input_payload_cmd_data[223 : 216];
  assign s2_inputDataBytes_28 = s2_input_payload_cmd_data[231 : 224];
  assign s2_inputDataBytes_29 = s2_input_payload_cmd_data[239 : 232];
  assign s2_inputDataBytes_30 = s2_input_payload_cmd_data[247 : 240];
  assign s2_inputDataBytes_31 = s2_input_payload_cmd_data[255 : 248];
  assign s2_byteLogic_0_lastUsed = (5'h0 == io_output_lastByteUsed);
  assign s2_byteLogic_0_inputMask = s2_input_payload_selValid[0];
  assign s2_byteLogic_0_inputData = _zz_s2_byteLogic_0_inputData;
  assign s2_byteLogic_0_outputMask = (s2_byteLogic_0_buffer_valid || (s2_input_valid && s2_byteLogic_0_inputMask));
  assign s2_byteLogic_0_outputData = (s2_byteLogic_0_buffer_valid ? s2_byteLogic_0_buffer_data : s2_byteLogic_0_inputData);
  always @(*) begin
    io_output_mask[0] = s2_byteLogic_0_outputMask;
    io_output_mask[1] = s2_byteLogic_1_outputMask;
    io_output_mask[2] = s2_byteLogic_2_outputMask;
    io_output_mask[3] = s2_byteLogic_3_outputMask;
    io_output_mask[4] = s2_byteLogic_4_outputMask;
    io_output_mask[5] = s2_byteLogic_5_outputMask;
    io_output_mask[6] = s2_byteLogic_6_outputMask;
    io_output_mask[7] = s2_byteLogic_7_outputMask;
    io_output_mask[8] = s2_byteLogic_8_outputMask;
    io_output_mask[9] = s2_byteLogic_9_outputMask;
    io_output_mask[10] = s2_byteLogic_10_outputMask;
    io_output_mask[11] = s2_byteLogic_11_outputMask;
    io_output_mask[12] = s2_byteLogic_12_outputMask;
    io_output_mask[13] = s2_byteLogic_13_outputMask;
    io_output_mask[14] = s2_byteLogic_14_outputMask;
    io_output_mask[15] = s2_byteLogic_15_outputMask;
    io_output_mask[16] = s2_byteLogic_16_outputMask;
    io_output_mask[17] = s2_byteLogic_17_outputMask;
    io_output_mask[18] = s2_byteLogic_18_outputMask;
    io_output_mask[19] = s2_byteLogic_19_outputMask;
    io_output_mask[20] = s2_byteLogic_20_outputMask;
    io_output_mask[21] = s2_byteLogic_21_outputMask;
    io_output_mask[22] = s2_byteLogic_22_outputMask;
    io_output_mask[23] = s2_byteLogic_23_outputMask;
    io_output_mask[24] = s2_byteLogic_24_outputMask;
    io_output_mask[25] = s2_byteLogic_25_outputMask;
    io_output_mask[26] = s2_byteLogic_26_outputMask;
    io_output_mask[27] = s2_byteLogic_27_outputMask;
    io_output_mask[28] = s2_byteLogic_28_outputMask;
    io_output_mask[29] = s2_byteLogic_29_outputMask;
    io_output_mask[30] = s2_byteLogic_30_outputMask;
    io_output_mask[31] = s2_byteLogic_31_outputMask;
  end

  always @(*) begin
    io_output_data[7 : 0] = s2_byteLogic_0_outputData;
    io_output_data[15 : 8] = s2_byteLogic_1_outputData;
    io_output_data[23 : 16] = s2_byteLogic_2_outputData;
    io_output_data[31 : 24] = s2_byteLogic_3_outputData;
    io_output_data[39 : 32] = s2_byteLogic_4_outputData;
    io_output_data[47 : 40] = s2_byteLogic_5_outputData;
    io_output_data[55 : 48] = s2_byteLogic_6_outputData;
    io_output_data[63 : 56] = s2_byteLogic_7_outputData;
    io_output_data[71 : 64] = s2_byteLogic_8_outputData;
    io_output_data[79 : 72] = s2_byteLogic_9_outputData;
    io_output_data[87 : 80] = s2_byteLogic_10_outputData;
    io_output_data[95 : 88] = s2_byteLogic_11_outputData;
    io_output_data[103 : 96] = s2_byteLogic_12_outputData;
    io_output_data[111 : 104] = s2_byteLogic_13_outputData;
    io_output_data[119 : 112] = s2_byteLogic_14_outputData;
    io_output_data[127 : 120] = s2_byteLogic_15_outputData;
    io_output_data[135 : 128] = s2_byteLogic_16_outputData;
    io_output_data[143 : 136] = s2_byteLogic_17_outputData;
    io_output_data[151 : 144] = s2_byteLogic_18_outputData;
    io_output_data[159 : 152] = s2_byteLogic_19_outputData;
    io_output_data[167 : 160] = s2_byteLogic_20_outputData;
    io_output_data[175 : 168] = s2_byteLogic_21_outputData;
    io_output_data[183 : 176] = s2_byteLogic_22_outputData;
    io_output_data[191 : 184] = s2_byteLogic_23_outputData;
    io_output_data[199 : 192] = s2_byteLogic_24_outputData;
    io_output_data[207 : 200] = s2_byteLogic_25_outputData;
    io_output_data[215 : 208] = s2_byteLogic_26_outputData;
    io_output_data[223 : 216] = s2_byteLogic_27_outputData;
    io_output_data[231 : 224] = s2_byteLogic_28_outputData;
    io_output_data[239 : 232] = s2_byteLogic_29_outputData;
    io_output_data[247 : 240] = s2_byteLogic_30_outputData;
    io_output_data[255 : 248] = s2_byteLogic_31_outputData;
  end

  assign when_DmaSg_l1493 = (s2_byteLogic_0_inputMask && ((! io_output_consume) || s2_byteLogic_0_buffer_valid));
  assign s2_byteLogic_1_lastUsed = (5'h01 == io_output_lastByteUsed);
  assign s2_byteLogic_1_inputMask = s2_input_payload_selValid[1];
  assign s2_byteLogic_1_inputData = _zz_s2_byteLogic_1_inputData;
  assign s2_byteLogic_1_outputMask = (s2_byteLogic_1_buffer_valid || (s2_input_valid && s2_byteLogic_1_inputMask));
  assign s2_byteLogic_1_outputData = (s2_byteLogic_1_buffer_valid ? s2_byteLogic_1_buffer_data : s2_byteLogic_1_inputData);
  assign when_DmaSg_l1493_1 = (s2_byteLogic_1_inputMask && ((! io_output_consume) || s2_byteLogic_1_buffer_valid));
  assign s2_byteLogic_2_lastUsed = (5'h02 == io_output_lastByteUsed);
  assign s2_byteLogic_2_inputMask = s2_input_payload_selValid[2];
  assign s2_byteLogic_2_inputData = _zz_s2_byteLogic_2_inputData;
  assign s2_byteLogic_2_outputMask = (s2_byteLogic_2_buffer_valid || (s2_input_valid && s2_byteLogic_2_inputMask));
  assign s2_byteLogic_2_outputData = (s2_byteLogic_2_buffer_valid ? s2_byteLogic_2_buffer_data : s2_byteLogic_2_inputData);
  assign when_DmaSg_l1493_2 = (s2_byteLogic_2_inputMask && ((! io_output_consume) || s2_byteLogic_2_buffer_valid));
  assign s2_byteLogic_3_lastUsed = (5'h03 == io_output_lastByteUsed);
  assign s2_byteLogic_3_inputMask = s2_input_payload_selValid[3];
  assign s2_byteLogic_3_inputData = _zz_s2_byteLogic_3_inputData;
  assign s2_byteLogic_3_outputMask = (s2_byteLogic_3_buffer_valid || (s2_input_valid && s2_byteLogic_3_inputMask));
  assign s2_byteLogic_3_outputData = (s2_byteLogic_3_buffer_valid ? s2_byteLogic_3_buffer_data : s2_byteLogic_3_inputData);
  assign when_DmaSg_l1493_3 = (s2_byteLogic_3_inputMask && ((! io_output_consume) || s2_byteLogic_3_buffer_valid));
  assign s2_byteLogic_4_lastUsed = (5'h04 == io_output_lastByteUsed);
  assign s2_byteLogic_4_inputMask = s2_input_payload_selValid[4];
  assign s2_byteLogic_4_inputData = _zz_s2_byteLogic_4_inputData;
  assign s2_byteLogic_4_outputMask = (s2_byteLogic_4_buffer_valid || (s2_input_valid && s2_byteLogic_4_inputMask));
  assign s2_byteLogic_4_outputData = (s2_byteLogic_4_buffer_valid ? s2_byteLogic_4_buffer_data : s2_byteLogic_4_inputData);
  assign when_DmaSg_l1493_4 = (s2_byteLogic_4_inputMask && ((! io_output_consume) || s2_byteLogic_4_buffer_valid));
  assign s2_byteLogic_5_lastUsed = (5'h05 == io_output_lastByteUsed);
  assign s2_byteLogic_5_inputMask = s2_input_payload_selValid[5];
  assign s2_byteLogic_5_inputData = _zz_s2_byteLogic_5_inputData;
  assign s2_byteLogic_5_outputMask = (s2_byteLogic_5_buffer_valid || (s2_input_valid && s2_byteLogic_5_inputMask));
  assign s2_byteLogic_5_outputData = (s2_byteLogic_5_buffer_valid ? s2_byteLogic_5_buffer_data : s2_byteLogic_5_inputData);
  assign when_DmaSg_l1493_5 = (s2_byteLogic_5_inputMask && ((! io_output_consume) || s2_byteLogic_5_buffer_valid));
  assign s2_byteLogic_6_lastUsed = (5'h06 == io_output_lastByteUsed);
  assign s2_byteLogic_6_inputMask = s2_input_payload_selValid[6];
  assign s2_byteLogic_6_inputData = _zz_s2_byteLogic_6_inputData;
  assign s2_byteLogic_6_outputMask = (s2_byteLogic_6_buffer_valid || (s2_input_valid && s2_byteLogic_6_inputMask));
  assign s2_byteLogic_6_outputData = (s2_byteLogic_6_buffer_valid ? s2_byteLogic_6_buffer_data : s2_byteLogic_6_inputData);
  assign when_DmaSg_l1493_6 = (s2_byteLogic_6_inputMask && ((! io_output_consume) || s2_byteLogic_6_buffer_valid));
  assign s2_byteLogic_7_lastUsed = (5'h07 == io_output_lastByteUsed);
  assign s2_byteLogic_7_inputMask = s2_input_payload_selValid[7];
  assign s2_byteLogic_7_inputData = _zz_s2_byteLogic_7_inputData;
  assign s2_byteLogic_7_outputMask = (s2_byteLogic_7_buffer_valid || (s2_input_valid && s2_byteLogic_7_inputMask));
  assign s2_byteLogic_7_outputData = (s2_byteLogic_7_buffer_valid ? s2_byteLogic_7_buffer_data : s2_byteLogic_7_inputData);
  assign when_DmaSg_l1493_7 = (s2_byteLogic_7_inputMask && ((! io_output_consume) || s2_byteLogic_7_buffer_valid));
  assign s2_byteLogic_8_lastUsed = (5'h08 == io_output_lastByteUsed);
  assign s2_byteLogic_8_inputMask = s2_input_payload_selValid[8];
  assign s2_byteLogic_8_inputData = _zz_s2_byteLogic_8_inputData;
  assign s2_byteLogic_8_outputMask = (s2_byteLogic_8_buffer_valid || (s2_input_valid && s2_byteLogic_8_inputMask));
  assign s2_byteLogic_8_outputData = (s2_byteLogic_8_buffer_valid ? s2_byteLogic_8_buffer_data : s2_byteLogic_8_inputData);
  assign when_DmaSg_l1493_8 = (s2_byteLogic_8_inputMask && ((! io_output_consume) || s2_byteLogic_8_buffer_valid));
  assign s2_byteLogic_9_lastUsed = (5'h09 == io_output_lastByteUsed);
  assign s2_byteLogic_9_inputMask = s2_input_payload_selValid[9];
  assign s2_byteLogic_9_inputData = _zz_s2_byteLogic_9_inputData;
  assign s2_byteLogic_9_outputMask = (s2_byteLogic_9_buffer_valid || (s2_input_valid && s2_byteLogic_9_inputMask));
  assign s2_byteLogic_9_outputData = (s2_byteLogic_9_buffer_valid ? s2_byteLogic_9_buffer_data : s2_byteLogic_9_inputData);
  assign when_DmaSg_l1493_9 = (s2_byteLogic_9_inputMask && ((! io_output_consume) || s2_byteLogic_9_buffer_valid));
  assign s2_byteLogic_10_lastUsed = (5'h0a == io_output_lastByteUsed);
  assign s2_byteLogic_10_inputMask = s2_input_payload_selValid[10];
  assign s2_byteLogic_10_inputData = _zz_s2_byteLogic_10_inputData;
  assign s2_byteLogic_10_outputMask = (s2_byteLogic_10_buffer_valid || (s2_input_valid && s2_byteLogic_10_inputMask));
  assign s2_byteLogic_10_outputData = (s2_byteLogic_10_buffer_valid ? s2_byteLogic_10_buffer_data : s2_byteLogic_10_inputData);
  assign when_DmaSg_l1493_10 = (s2_byteLogic_10_inputMask && ((! io_output_consume) || s2_byteLogic_10_buffer_valid));
  assign s2_byteLogic_11_lastUsed = (5'h0b == io_output_lastByteUsed);
  assign s2_byteLogic_11_inputMask = s2_input_payload_selValid[11];
  assign s2_byteLogic_11_inputData = _zz_s2_byteLogic_11_inputData;
  assign s2_byteLogic_11_outputMask = (s2_byteLogic_11_buffer_valid || (s2_input_valid && s2_byteLogic_11_inputMask));
  assign s2_byteLogic_11_outputData = (s2_byteLogic_11_buffer_valid ? s2_byteLogic_11_buffer_data : s2_byteLogic_11_inputData);
  assign when_DmaSg_l1493_11 = (s2_byteLogic_11_inputMask && ((! io_output_consume) || s2_byteLogic_11_buffer_valid));
  assign s2_byteLogic_12_lastUsed = (5'h0c == io_output_lastByteUsed);
  assign s2_byteLogic_12_inputMask = s2_input_payload_selValid[12];
  assign s2_byteLogic_12_inputData = _zz_s2_byteLogic_12_inputData;
  assign s2_byteLogic_12_outputMask = (s2_byteLogic_12_buffer_valid || (s2_input_valid && s2_byteLogic_12_inputMask));
  assign s2_byteLogic_12_outputData = (s2_byteLogic_12_buffer_valid ? s2_byteLogic_12_buffer_data : s2_byteLogic_12_inputData);
  assign when_DmaSg_l1493_12 = (s2_byteLogic_12_inputMask && ((! io_output_consume) || s2_byteLogic_12_buffer_valid));
  assign s2_byteLogic_13_lastUsed = (5'h0d == io_output_lastByteUsed);
  assign s2_byteLogic_13_inputMask = s2_input_payload_selValid[13];
  assign s2_byteLogic_13_inputData = _zz_s2_byteLogic_13_inputData;
  assign s2_byteLogic_13_outputMask = (s2_byteLogic_13_buffer_valid || (s2_input_valid && s2_byteLogic_13_inputMask));
  assign s2_byteLogic_13_outputData = (s2_byteLogic_13_buffer_valid ? s2_byteLogic_13_buffer_data : s2_byteLogic_13_inputData);
  assign when_DmaSg_l1493_13 = (s2_byteLogic_13_inputMask && ((! io_output_consume) || s2_byteLogic_13_buffer_valid));
  assign s2_byteLogic_14_lastUsed = (5'h0e == io_output_lastByteUsed);
  assign s2_byteLogic_14_inputMask = s2_input_payload_selValid[14];
  assign s2_byteLogic_14_inputData = _zz_s2_byteLogic_14_inputData;
  assign s2_byteLogic_14_outputMask = (s2_byteLogic_14_buffer_valid || (s2_input_valid && s2_byteLogic_14_inputMask));
  assign s2_byteLogic_14_outputData = (s2_byteLogic_14_buffer_valid ? s2_byteLogic_14_buffer_data : s2_byteLogic_14_inputData);
  assign when_DmaSg_l1493_14 = (s2_byteLogic_14_inputMask && ((! io_output_consume) || s2_byteLogic_14_buffer_valid));
  assign s2_byteLogic_15_lastUsed = (5'h0f == io_output_lastByteUsed);
  assign s2_byteLogic_15_inputMask = s2_input_payload_selValid[15];
  assign s2_byteLogic_15_inputData = _zz_s2_byteLogic_15_inputData;
  assign s2_byteLogic_15_outputMask = (s2_byteLogic_15_buffer_valid || (s2_input_valid && s2_byteLogic_15_inputMask));
  assign s2_byteLogic_15_outputData = (s2_byteLogic_15_buffer_valid ? s2_byteLogic_15_buffer_data : s2_byteLogic_15_inputData);
  assign when_DmaSg_l1493_15 = (s2_byteLogic_15_inputMask && ((! io_output_consume) || s2_byteLogic_15_buffer_valid));
  assign s2_byteLogic_16_lastUsed = (5'h10 == io_output_lastByteUsed);
  assign s2_byteLogic_16_inputMask = s2_input_payload_selValid[16];
  assign s2_byteLogic_16_inputData = _zz_s2_byteLogic_16_inputData;
  assign s2_byteLogic_16_outputMask = (s2_byteLogic_16_buffer_valid || (s2_input_valid && s2_byteLogic_16_inputMask));
  assign s2_byteLogic_16_outputData = (s2_byteLogic_16_buffer_valid ? s2_byteLogic_16_buffer_data : s2_byteLogic_16_inputData);
  assign when_DmaSg_l1493_16 = (s2_byteLogic_16_inputMask && ((! io_output_consume) || s2_byteLogic_16_buffer_valid));
  assign s2_byteLogic_17_lastUsed = (5'h11 == io_output_lastByteUsed);
  assign s2_byteLogic_17_inputMask = s2_input_payload_selValid[17];
  assign s2_byteLogic_17_inputData = _zz_s2_byteLogic_17_inputData;
  assign s2_byteLogic_17_outputMask = (s2_byteLogic_17_buffer_valid || (s2_input_valid && s2_byteLogic_17_inputMask));
  assign s2_byteLogic_17_outputData = (s2_byteLogic_17_buffer_valid ? s2_byteLogic_17_buffer_data : s2_byteLogic_17_inputData);
  assign when_DmaSg_l1493_17 = (s2_byteLogic_17_inputMask && ((! io_output_consume) || s2_byteLogic_17_buffer_valid));
  assign s2_byteLogic_18_lastUsed = (5'h12 == io_output_lastByteUsed);
  assign s2_byteLogic_18_inputMask = s2_input_payload_selValid[18];
  assign s2_byteLogic_18_inputData = _zz_s2_byteLogic_18_inputData;
  assign s2_byteLogic_18_outputMask = (s2_byteLogic_18_buffer_valid || (s2_input_valid && s2_byteLogic_18_inputMask));
  assign s2_byteLogic_18_outputData = (s2_byteLogic_18_buffer_valid ? s2_byteLogic_18_buffer_data : s2_byteLogic_18_inputData);
  assign when_DmaSg_l1493_18 = (s2_byteLogic_18_inputMask && ((! io_output_consume) || s2_byteLogic_18_buffer_valid));
  assign s2_byteLogic_19_lastUsed = (5'h13 == io_output_lastByteUsed);
  assign s2_byteLogic_19_inputMask = s2_input_payload_selValid[19];
  assign s2_byteLogic_19_inputData = _zz_s2_byteLogic_19_inputData;
  assign s2_byteLogic_19_outputMask = (s2_byteLogic_19_buffer_valid || (s2_input_valid && s2_byteLogic_19_inputMask));
  assign s2_byteLogic_19_outputData = (s2_byteLogic_19_buffer_valid ? s2_byteLogic_19_buffer_data : s2_byteLogic_19_inputData);
  assign when_DmaSg_l1493_19 = (s2_byteLogic_19_inputMask && ((! io_output_consume) || s2_byteLogic_19_buffer_valid));
  assign s2_byteLogic_20_lastUsed = (5'h14 == io_output_lastByteUsed);
  assign s2_byteLogic_20_inputMask = s2_input_payload_selValid[20];
  assign s2_byteLogic_20_inputData = _zz_s2_byteLogic_20_inputData;
  assign s2_byteLogic_20_outputMask = (s2_byteLogic_20_buffer_valid || (s2_input_valid && s2_byteLogic_20_inputMask));
  assign s2_byteLogic_20_outputData = (s2_byteLogic_20_buffer_valid ? s2_byteLogic_20_buffer_data : s2_byteLogic_20_inputData);
  assign when_DmaSg_l1493_20 = (s2_byteLogic_20_inputMask && ((! io_output_consume) || s2_byteLogic_20_buffer_valid));
  assign s2_byteLogic_21_lastUsed = (5'h15 == io_output_lastByteUsed);
  assign s2_byteLogic_21_inputMask = s2_input_payload_selValid[21];
  assign s2_byteLogic_21_inputData = _zz_s2_byteLogic_21_inputData;
  assign s2_byteLogic_21_outputMask = (s2_byteLogic_21_buffer_valid || (s2_input_valid && s2_byteLogic_21_inputMask));
  assign s2_byteLogic_21_outputData = (s2_byteLogic_21_buffer_valid ? s2_byteLogic_21_buffer_data : s2_byteLogic_21_inputData);
  assign when_DmaSg_l1493_21 = (s2_byteLogic_21_inputMask && ((! io_output_consume) || s2_byteLogic_21_buffer_valid));
  assign s2_byteLogic_22_lastUsed = (5'h16 == io_output_lastByteUsed);
  assign s2_byteLogic_22_inputMask = s2_input_payload_selValid[22];
  assign s2_byteLogic_22_inputData = _zz_s2_byteLogic_22_inputData;
  assign s2_byteLogic_22_outputMask = (s2_byteLogic_22_buffer_valid || (s2_input_valid && s2_byteLogic_22_inputMask));
  assign s2_byteLogic_22_outputData = (s2_byteLogic_22_buffer_valid ? s2_byteLogic_22_buffer_data : s2_byteLogic_22_inputData);
  assign when_DmaSg_l1493_22 = (s2_byteLogic_22_inputMask && ((! io_output_consume) || s2_byteLogic_22_buffer_valid));
  assign s2_byteLogic_23_lastUsed = (5'h17 == io_output_lastByteUsed);
  assign s2_byteLogic_23_inputMask = s2_input_payload_selValid[23];
  assign s2_byteLogic_23_inputData = _zz_s2_byteLogic_23_inputData;
  assign s2_byteLogic_23_outputMask = (s2_byteLogic_23_buffer_valid || (s2_input_valid && s2_byteLogic_23_inputMask));
  assign s2_byteLogic_23_outputData = (s2_byteLogic_23_buffer_valid ? s2_byteLogic_23_buffer_data : s2_byteLogic_23_inputData);
  assign when_DmaSg_l1493_23 = (s2_byteLogic_23_inputMask && ((! io_output_consume) || s2_byteLogic_23_buffer_valid));
  assign s2_byteLogic_24_lastUsed = (5'h18 == io_output_lastByteUsed);
  assign s2_byteLogic_24_inputMask = s2_input_payload_selValid[24];
  assign s2_byteLogic_24_inputData = _zz_s2_byteLogic_24_inputData;
  assign s2_byteLogic_24_outputMask = (s2_byteLogic_24_buffer_valid || (s2_input_valid && s2_byteLogic_24_inputMask));
  assign s2_byteLogic_24_outputData = (s2_byteLogic_24_buffer_valid ? s2_byteLogic_24_buffer_data : s2_byteLogic_24_inputData);
  assign when_DmaSg_l1493_24 = (s2_byteLogic_24_inputMask && ((! io_output_consume) || s2_byteLogic_24_buffer_valid));
  assign s2_byteLogic_25_lastUsed = (5'h19 == io_output_lastByteUsed);
  assign s2_byteLogic_25_inputMask = s2_input_payload_selValid[25];
  assign s2_byteLogic_25_inputData = _zz_s2_byteLogic_25_inputData;
  assign s2_byteLogic_25_outputMask = (s2_byteLogic_25_buffer_valid || (s2_input_valid && s2_byteLogic_25_inputMask));
  assign s2_byteLogic_25_outputData = (s2_byteLogic_25_buffer_valid ? s2_byteLogic_25_buffer_data : s2_byteLogic_25_inputData);
  assign when_DmaSg_l1493_25 = (s2_byteLogic_25_inputMask && ((! io_output_consume) || s2_byteLogic_25_buffer_valid));
  assign s2_byteLogic_26_lastUsed = (5'h1a == io_output_lastByteUsed);
  assign s2_byteLogic_26_inputMask = s2_input_payload_selValid[26];
  assign s2_byteLogic_26_inputData = _zz_s2_byteLogic_26_inputData;
  assign s2_byteLogic_26_outputMask = (s2_byteLogic_26_buffer_valid || (s2_input_valid && s2_byteLogic_26_inputMask));
  assign s2_byteLogic_26_outputData = (s2_byteLogic_26_buffer_valid ? s2_byteLogic_26_buffer_data : s2_byteLogic_26_inputData);
  assign when_DmaSg_l1493_26 = (s2_byteLogic_26_inputMask && ((! io_output_consume) || s2_byteLogic_26_buffer_valid));
  assign s2_byteLogic_27_lastUsed = (5'h1b == io_output_lastByteUsed);
  assign s2_byteLogic_27_inputMask = s2_input_payload_selValid[27];
  assign s2_byteLogic_27_inputData = _zz_s2_byteLogic_27_inputData;
  assign s2_byteLogic_27_outputMask = (s2_byteLogic_27_buffer_valid || (s2_input_valid && s2_byteLogic_27_inputMask));
  assign s2_byteLogic_27_outputData = (s2_byteLogic_27_buffer_valid ? s2_byteLogic_27_buffer_data : s2_byteLogic_27_inputData);
  assign when_DmaSg_l1493_27 = (s2_byteLogic_27_inputMask && ((! io_output_consume) || s2_byteLogic_27_buffer_valid));
  assign s2_byteLogic_28_lastUsed = (5'h1c == io_output_lastByteUsed);
  assign s2_byteLogic_28_inputMask = s2_input_payload_selValid[28];
  assign s2_byteLogic_28_inputData = _zz_s2_byteLogic_28_inputData;
  assign s2_byteLogic_28_outputMask = (s2_byteLogic_28_buffer_valid || (s2_input_valid && s2_byteLogic_28_inputMask));
  assign s2_byteLogic_28_outputData = (s2_byteLogic_28_buffer_valid ? s2_byteLogic_28_buffer_data : s2_byteLogic_28_inputData);
  assign when_DmaSg_l1493_28 = (s2_byteLogic_28_inputMask && ((! io_output_consume) || s2_byteLogic_28_buffer_valid));
  assign s2_byteLogic_29_lastUsed = (5'h1d == io_output_lastByteUsed);
  assign s2_byteLogic_29_inputMask = s2_input_payload_selValid[29];
  assign s2_byteLogic_29_inputData = _zz_s2_byteLogic_29_inputData;
  assign s2_byteLogic_29_outputMask = (s2_byteLogic_29_buffer_valid || (s2_input_valid && s2_byteLogic_29_inputMask));
  assign s2_byteLogic_29_outputData = (s2_byteLogic_29_buffer_valid ? s2_byteLogic_29_buffer_data : s2_byteLogic_29_inputData);
  assign when_DmaSg_l1493_29 = (s2_byteLogic_29_inputMask && ((! io_output_consume) || s2_byteLogic_29_buffer_valid));
  assign s2_byteLogic_30_lastUsed = (5'h1e == io_output_lastByteUsed);
  assign s2_byteLogic_30_inputMask = s2_input_payload_selValid[30];
  assign s2_byteLogic_30_inputData = _zz_s2_byteLogic_30_inputData;
  assign s2_byteLogic_30_outputMask = (s2_byteLogic_30_buffer_valid || (s2_input_valid && s2_byteLogic_30_inputMask));
  assign s2_byteLogic_30_outputData = (s2_byteLogic_30_buffer_valid ? s2_byteLogic_30_buffer_data : s2_byteLogic_30_inputData);
  assign when_DmaSg_l1493_30 = (s2_byteLogic_30_inputMask && ((! io_output_consume) || s2_byteLogic_30_buffer_valid));
  assign s2_byteLogic_31_lastUsed = (5'h1f == io_output_lastByteUsed);
  assign s2_byteLogic_31_inputMask = s2_input_payload_selValid[31];
  assign s2_byteLogic_31_inputData = _zz_s2_byteLogic_31_inputData;
  assign s2_byteLogic_31_outputMask = (s2_byteLogic_31_buffer_valid || (s2_input_valid && s2_byteLogic_31_inputMask));
  assign s2_byteLogic_31_outputData = (s2_byteLogic_31_buffer_valid ? s2_byteLogic_31_buffer_data : s2_byteLogic_31_inputData);
  assign when_DmaSg_l1493_31 = (s2_byteLogic_31_inputMask && ((! io_output_consume) || s2_byteLogic_31_buffer_valid));
  assign _zz_io_output_usedUntil = (((((((((((((((s2_byteLogic_1_lastUsed || s2_byteLogic_3_lastUsed) || s2_byteLogic_5_lastUsed) || s2_byteLogic_7_lastUsed) || s2_byteLogic_9_lastUsed) || s2_byteLogic_11_lastUsed) || s2_byteLogic_13_lastUsed) || s2_byteLogic_15_lastUsed) || s2_byteLogic_17_lastUsed) || s2_byteLogic_19_lastUsed) || s2_byteLogic_21_lastUsed) || s2_byteLogic_23_lastUsed) || s2_byteLogic_25_lastUsed) || s2_byteLogic_27_lastUsed) || s2_byteLogic_29_lastUsed) || s2_byteLogic_31_lastUsed);
  assign _zz_io_output_usedUntil_1 = (((((((((((((((s2_byteLogic_2_lastUsed || s2_byteLogic_3_lastUsed) || s2_byteLogic_6_lastUsed) || s2_byteLogic_7_lastUsed) || s2_byteLogic_10_lastUsed) || s2_byteLogic_11_lastUsed) || s2_byteLogic_14_lastUsed) || s2_byteLogic_15_lastUsed) || s2_byteLogic_18_lastUsed) || s2_byteLogic_19_lastUsed) || s2_byteLogic_22_lastUsed) || s2_byteLogic_23_lastUsed) || s2_byteLogic_26_lastUsed) || s2_byteLogic_27_lastUsed) || s2_byteLogic_30_lastUsed) || s2_byteLogic_31_lastUsed);
  assign _zz_io_output_usedUntil_2 = (((((((((((((((s2_byteLogic_4_lastUsed || s2_byteLogic_5_lastUsed) || s2_byteLogic_6_lastUsed) || s2_byteLogic_7_lastUsed) || s2_byteLogic_12_lastUsed) || s2_byteLogic_13_lastUsed) || s2_byteLogic_14_lastUsed) || s2_byteLogic_15_lastUsed) || s2_byteLogic_20_lastUsed) || s2_byteLogic_21_lastUsed) || s2_byteLogic_22_lastUsed) || s2_byteLogic_23_lastUsed) || s2_byteLogic_28_lastUsed) || s2_byteLogic_29_lastUsed) || s2_byteLogic_30_lastUsed) || s2_byteLogic_31_lastUsed);
  assign _zz_io_output_usedUntil_3 = (((((((((((((((s2_byteLogic_8_lastUsed || s2_byteLogic_9_lastUsed) || s2_byteLogic_10_lastUsed) || s2_byteLogic_11_lastUsed) || s2_byteLogic_12_lastUsed) || s2_byteLogic_13_lastUsed) || s2_byteLogic_14_lastUsed) || s2_byteLogic_15_lastUsed) || s2_byteLogic_24_lastUsed) || s2_byteLogic_25_lastUsed) || s2_byteLogic_26_lastUsed) || s2_byteLogic_27_lastUsed) || s2_byteLogic_28_lastUsed) || s2_byteLogic_29_lastUsed) || s2_byteLogic_30_lastUsed) || s2_byteLogic_31_lastUsed);
  assign _zz_io_output_usedUntil_4 = (((((((((((((((s2_byteLogic_16_lastUsed || s2_byteLogic_17_lastUsed) || s2_byteLogic_18_lastUsed) || s2_byteLogic_19_lastUsed) || s2_byteLogic_20_lastUsed) || s2_byteLogic_21_lastUsed) || s2_byteLogic_22_lastUsed) || s2_byteLogic_23_lastUsed) || s2_byteLogic_24_lastUsed) || s2_byteLogic_25_lastUsed) || s2_byteLogic_26_lastUsed) || s2_byteLogic_27_lastUsed) || s2_byteLogic_28_lastUsed) || s2_byteLogic_29_lastUsed) || s2_byteLogic_30_lastUsed) || s2_byteLogic_31_lastUsed);
  assign io_output_usedUntil = _zz_io_output_usedUntil_5;
  always @(posedge clk) begin
    if(reset) begin
      io_input_rValid <= 1'b0;
      s0_output_rValid <= 1'b0;
      s1_output_rValid <= 1'b0;
    end else begin
      if(io_input_ready) begin
        io_input_rValid <= io_input_valid;
      end
      if(io_flush) begin
        io_input_rValid <= 1'b0;
      end
      if(s0_output_ready) begin
        s0_output_rValid <= s0_output_valid;
      end
      if(io_flush) begin
        s0_output_rValid <= 1'b0;
      end
      if(s1_output_ready) begin
        s1_output_rValid <= s1_output_valid;
      end
      if(io_flush) begin
        s1_output_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_input_ready) begin
      io_input_rData_data <= io_input_payload_data;
      io_input_rData_mask <= io_input_payload_mask;
    end
    if(s0_output_ready) begin
      s0_output_rData_cmd_data <= s0_output_payload_cmd_data;
      s0_output_rData_cmd_mask <= s0_output_payload_cmd_mask;
      s0_output_rData_countOnes_0 <= s0_output_payload_countOnes_0;
      s0_output_rData_countOnes_1 <= s0_output_payload_countOnes_1;
      s0_output_rData_countOnes_2 <= s0_output_payload_countOnes_2;
      s0_output_rData_countOnes_3 <= s0_output_payload_countOnes_3;
      s0_output_rData_countOnes_4 <= s0_output_payload_countOnes_4;
      s0_output_rData_countOnes_5 <= s0_output_payload_countOnes_5;
      s0_output_rData_countOnes_6 <= s0_output_payload_countOnes_6;
      s0_output_rData_countOnes_7 <= s0_output_payload_countOnes_7;
      s0_output_rData_countOnes_8 <= s0_output_payload_countOnes_8;
      s0_output_rData_countOnes_9 <= s0_output_payload_countOnes_9;
      s0_output_rData_countOnes_10 <= s0_output_payload_countOnes_10;
      s0_output_rData_countOnes_11 <= s0_output_payload_countOnes_11;
      s0_output_rData_countOnes_12 <= s0_output_payload_countOnes_12;
      s0_output_rData_countOnes_13 <= s0_output_payload_countOnes_13;
      s0_output_rData_countOnes_14 <= s0_output_payload_countOnes_14;
      s0_output_rData_countOnes_15 <= s0_output_payload_countOnes_15;
      s0_output_rData_countOnes_16 <= s0_output_payload_countOnes_16;
      s0_output_rData_countOnes_17 <= s0_output_payload_countOnes_17;
      s0_output_rData_countOnes_18 <= s0_output_payload_countOnes_18;
      s0_output_rData_countOnes_19 <= s0_output_payload_countOnes_19;
      s0_output_rData_countOnes_20 <= s0_output_payload_countOnes_20;
      s0_output_rData_countOnes_21 <= s0_output_payload_countOnes_21;
      s0_output_rData_countOnes_22 <= s0_output_payload_countOnes_22;
      s0_output_rData_countOnes_23 <= s0_output_payload_countOnes_23;
      s0_output_rData_countOnes_24 <= s0_output_payload_countOnes_24;
      s0_output_rData_countOnes_25 <= s0_output_payload_countOnes_25;
      s0_output_rData_countOnes_26 <= s0_output_payload_countOnes_26;
      s0_output_rData_countOnes_27 <= s0_output_payload_countOnes_27;
      s0_output_rData_countOnes_28 <= s0_output_payload_countOnes_28;
      s0_output_rData_countOnes_29 <= s0_output_payload_countOnes_29;
      s0_output_rData_countOnes_30 <= s0_output_payload_countOnes_30;
      s0_output_rData_countOnes_31 <= s0_output_payload_countOnes_31;
    end
    if(s1_input_fire) begin
      s1_offset <= s1_offsetNext[4:0];
    end
    if(io_flush) begin
      s1_offset <= io_offset;
    end
    if(s1_input_fire) begin
      s1_byteCounter <= (s1_byteCounter + _zz_s1_byteCounter);
    end
    if(io_flush) begin
      s1_byteCounter <= 14'h0;
    end
    if(s1_output_ready) begin
      s1_output_rData_cmd_data <= s1_output_payload_cmd_data;
      s1_output_rData_cmd_mask <= s1_output_payload_cmd_mask;
      s1_output_rData_index_0 <= s1_output_payload_index_0;
      s1_output_rData_index_1 <= s1_output_payload_index_1;
      s1_output_rData_index_2 <= s1_output_payload_index_2;
      s1_output_rData_index_3 <= s1_output_payload_index_3;
      s1_output_rData_index_4 <= s1_output_payload_index_4;
      s1_output_rData_index_5 <= s1_output_payload_index_5;
      s1_output_rData_index_6 <= s1_output_payload_index_6;
      s1_output_rData_index_7 <= s1_output_payload_index_7;
      s1_output_rData_index_8 <= s1_output_payload_index_8;
      s1_output_rData_index_9 <= s1_output_payload_index_9;
      s1_output_rData_index_10 <= s1_output_payload_index_10;
      s1_output_rData_index_11 <= s1_output_payload_index_11;
      s1_output_rData_index_12 <= s1_output_payload_index_12;
      s1_output_rData_index_13 <= s1_output_payload_index_13;
      s1_output_rData_index_14 <= s1_output_payload_index_14;
      s1_output_rData_index_15 <= s1_output_payload_index_15;
      s1_output_rData_index_16 <= s1_output_payload_index_16;
      s1_output_rData_index_17 <= s1_output_payload_index_17;
      s1_output_rData_index_18 <= s1_output_payload_index_18;
      s1_output_rData_index_19 <= s1_output_payload_index_19;
      s1_output_rData_index_20 <= s1_output_payload_index_20;
      s1_output_rData_index_21 <= s1_output_payload_index_21;
      s1_output_rData_index_22 <= s1_output_payload_index_22;
      s1_output_rData_index_23 <= s1_output_payload_index_23;
      s1_output_rData_index_24 <= s1_output_payload_index_24;
      s1_output_rData_index_25 <= s1_output_payload_index_25;
      s1_output_rData_index_26 <= s1_output_payload_index_26;
      s1_output_rData_index_27 <= s1_output_payload_index_27;
      s1_output_rData_index_28 <= s1_output_payload_index_28;
      s1_output_rData_index_29 <= s1_output_payload_index_29;
      s1_output_rData_index_30 <= s1_output_payload_index_30;
      s1_output_rData_index_31 <= s1_output_payload_index_31;
      s1_output_rData_last <= s1_output_payload_last;
      s1_output_rData_sel_0 <= s1_output_payload_sel_0;
      s1_output_rData_sel_1 <= s1_output_payload_sel_1;
      s1_output_rData_sel_2 <= s1_output_payload_sel_2;
      s1_output_rData_sel_3 <= s1_output_payload_sel_3;
      s1_output_rData_sel_4 <= s1_output_payload_sel_4;
      s1_output_rData_sel_5 <= s1_output_payload_sel_5;
      s1_output_rData_sel_6 <= s1_output_payload_sel_6;
      s1_output_rData_sel_7 <= s1_output_payload_sel_7;
      s1_output_rData_sel_8 <= s1_output_payload_sel_8;
      s1_output_rData_sel_9 <= s1_output_payload_sel_9;
      s1_output_rData_sel_10 <= s1_output_payload_sel_10;
      s1_output_rData_sel_11 <= s1_output_payload_sel_11;
      s1_output_rData_sel_12 <= s1_output_payload_sel_12;
      s1_output_rData_sel_13 <= s1_output_payload_sel_13;
      s1_output_rData_sel_14 <= s1_output_payload_sel_14;
      s1_output_rData_sel_15 <= s1_output_payload_sel_15;
      s1_output_rData_sel_16 <= s1_output_payload_sel_16;
      s1_output_rData_sel_17 <= s1_output_payload_sel_17;
      s1_output_rData_sel_18 <= s1_output_payload_sel_18;
      s1_output_rData_sel_19 <= s1_output_payload_sel_19;
      s1_output_rData_sel_20 <= s1_output_payload_sel_20;
      s1_output_rData_sel_21 <= s1_output_payload_sel_21;
      s1_output_rData_sel_22 <= s1_output_payload_sel_22;
      s1_output_rData_sel_23 <= s1_output_payload_sel_23;
      s1_output_rData_sel_24 <= s1_output_payload_sel_24;
      s1_output_rData_sel_25 <= s1_output_payload_sel_25;
      s1_output_rData_sel_26 <= s1_output_payload_sel_26;
      s1_output_rData_sel_27 <= s1_output_payload_sel_27;
      s1_output_rData_sel_28 <= s1_output_payload_sel_28;
      s1_output_rData_sel_29 <= s1_output_payload_sel_29;
      s1_output_rData_sel_30 <= s1_output_payload_sel_30;
      s1_output_rData_sel_31 <= s1_output_payload_sel_31;
      s1_output_rData_selValid <= s1_output_payload_selValid;
    end
    if(io_output_consume) begin
      s2_byteLogic_0_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_0_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493) begin
        s2_byteLogic_0_buffer_valid <= 1'b1;
        s2_byteLogic_0_buffer_data <= s2_byteLogic_0_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_0_buffer_valid <= (5'h0 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_1_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_1_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_1) begin
        s2_byteLogic_1_buffer_valid <= 1'b1;
        s2_byteLogic_1_buffer_data <= s2_byteLogic_1_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_1_buffer_valid <= (5'h01 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_2_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_2_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_2) begin
        s2_byteLogic_2_buffer_valid <= 1'b1;
        s2_byteLogic_2_buffer_data <= s2_byteLogic_2_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_2_buffer_valid <= (5'h02 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_3_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_3_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_3) begin
        s2_byteLogic_3_buffer_valid <= 1'b1;
        s2_byteLogic_3_buffer_data <= s2_byteLogic_3_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_3_buffer_valid <= (5'h03 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_4_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_4_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_4) begin
        s2_byteLogic_4_buffer_valid <= 1'b1;
        s2_byteLogic_4_buffer_data <= s2_byteLogic_4_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_4_buffer_valid <= (5'h04 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_5_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_5_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_5) begin
        s2_byteLogic_5_buffer_valid <= 1'b1;
        s2_byteLogic_5_buffer_data <= s2_byteLogic_5_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_5_buffer_valid <= (5'h05 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_6_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_6_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_6) begin
        s2_byteLogic_6_buffer_valid <= 1'b1;
        s2_byteLogic_6_buffer_data <= s2_byteLogic_6_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_6_buffer_valid <= (5'h06 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_7_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_7_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_7) begin
        s2_byteLogic_7_buffer_valid <= 1'b1;
        s2_byteLogic_7_buffer_data <= s2_byteLogic_7_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_7_buffer_valid <= (5'h07 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_8_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_8_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_8) begin
        s2_byteLogic_8_buffer_valid <= 1'b1;
        s2_byteLogic_8_buffer_data <= s2_byteLogic_8_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_8_buffer_valid <= (5'h08 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_9_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_9_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_9) begin
        s2_byteLogic_9_buffer_valid <= 1'b1;
        s2_byteLogic_9_buffer_data <= s2_byteLogic_9_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_9_buffer_valid <= (5'h09 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_10_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_10_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_10) begin
        s2_byteLogic_10_buffer_valid <= 1'b1;
        s2_byteLogic_10_buffer_data <= s2_byteLogic_10_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_10_buffer_valid <= (5'h0a < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_11_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_11_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_11) begin
        s2_byteLogic_11_buffer_valid <= 1'b1;
        s2_byteLogic_11_buffer_data <= s2_byteLogic_11_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_11_buffer_valid <= (5'h0b < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_12_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_12_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_12) begin
        s2_byteLogic_12_buffer_valid <= 1'b1;
        s2_byteLogic_12_buffer_data <= s2_byteLogic_12_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_12_buffer_valid <= (5'h0c < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_13_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_13_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_13) begin
        s2_byteLogic_13_buffer_valid <= 1'b1;
        s2_byteLogic_13_buffer_data <= s2_byteLogic_13_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_13_buffer_valid <= (5'h0d < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_14_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_14_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_14) begin
        s2_byteLogic_14_buffer_valid <= 1'b1;
        s2_byteLogic_14_buffer_data <= s2_byteLogic_14_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_14_buffer_valid <= (5'h0e < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_15_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_15_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_15) begin
        s2_byteLogic_15_buffer_valid <= 1'b1;
        s2_byteLogic_15_buffer_data <= s2_byteLogic_15_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_15_buffer_valid <= (5'h0f < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_16_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_16_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_16) begin
        s2_byteLogic_16_buffer_valid <= 1'b1;
        s2_byteLogic_16_buffer_data <= s2_byteLogic_16_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_16_buffer_valid <= (5'h10 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_17_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_17_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_17) begin
        s2_byteLogic_17_buffer_valid <= 1'b1;
        s2_byteLogic_17_buffer_data <= s2_byteLogic_17_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_17_buffer_valid <= (5'h11 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_18_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_18_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_18) begin
        s2_byteLogic_18_buffer_valid <= 1'b1;
        s2_byteLogic_18_buffer_data <= s2_byteLogic_18_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_18_buffer_valid <= (5'h12 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_19_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_19_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_19) begin
        s2_byteLogic_19_buffer_valid <= 1'b1;
        s2_byteLogic_19_buffer_data <= s2_byteLogic_19_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_19_buffer_valid <= (5'h13 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_20_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_20_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_20) begin
        s2_byteLogic_20_buffer_valid <= 1'b1;
        s2_byteLogic_20_buffer_data <= s2_byteLogic_20_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_20_buffer_valid <= (5'h14 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_21_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_21_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_21) begin
        s2_byteLogic_21_buffer_valid <= 1'b1;
        s2_byteLogic_21_buffer_data <= s2_byteLogic_21_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_21_buffer_valid <= (5'h15 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_22_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_22_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_22) begin
        s2_byteLogic_22_buffer_valid <= 1'b1;
        s2_byteLogic_22_buffer_data <= s2_byteLogic_22_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_22_buffer_valid <= (5'h16 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_23_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_23_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_23) begin
        s2_byteLogic_23_buffer_valid <= 1'b1;
        s2_byteLogic_23_buffer_data <= s2_byteLogic_23_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_23_buffer_valid <= (5'h17 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_24_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_24_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_24) begin
        s2_byteLogic_24_buffer_valid <= 1'b1;
        s2_byteLogic_24_buffer_data <= s2_byteLogic_24_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_24_buffer_valid <= (5'h18 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_25_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_25_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_25) begin
        s2_byteLogic_25_buffer_valid <= 1'b1;
        s2_byteLogic_25_buffer_data <= s2_byteLogic_25_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_25_buffer_valid <= (5'h19 < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_26_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_26_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_26) begin
        s2_byteLogic_26_buffer_valid <= 1'b1;
        s2_byteLogic_26_buffer_data <= s2_byteLogic_26_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_26_buffer_valid <= (5'h1a < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_27_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_27_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_27) begin
        s2_byteLogic_27_buffer_valid <= 1'b1;
        s2_byteLogic_27_buffer_data <= s2_byteLogic_27_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_27_buffer_valid <= (5'h1b < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_28_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_28_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_28) begin
        s2_byteLogic_28_buffer_valid <= 1'b1;
        s2_byteLogic_28_buffer_data <= s2_byteLogic_28_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_28_buffer_valid <= (5'h1c < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_29_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_29_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_29) begin
        s2_byteLogic_29_buffer_valid <= 1'b1;
        s2_byteLogic_29_buffer_data <= s2_byteLogic_29_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_29_buffer_valid <= (5'h1d < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_30_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_30_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_30) begin
        s2_byteLogic_30_buffer_valid <= 1'b1;
        s2_byteLogic_30_buffer_data <= s2_byteLogic_30_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_30_buffer_valid <= (5'h1e < io_offset);
    end
    if(io_output_consume) begin
      s2_byteLogic_31_buffer_valid <= 1'b0;
    end
    if(s2_input_fire) begin
      if(s2_input_payload_last) begin
        s2_byteLogic_31_buffer_valid <= 1'b0;
      end
      if(when_DmaSg_l1493_31) begin
        s2_byteLogic_31_buffer_valid <= 1'b1;
        s2_byteLogic_31_buffer_data <= s2_byteLogic_31_inputData;
      end
    end
    if(io_flush) begin
      s2_byteLogic_31_buffer_valid <= (5'h1f < io_offset);
    end
  end


endmodule

module EfxDMA_DmaMemoryCore (
  input  wire          io_writes_0_cmd_valid,
  output wire          io_writes_0_cmd_ready,
  input  wire [12:0]   io_writes_0_cmd_payload_address,
  input  wire [127:0]  io_writes_0_cmd_payload_data,
  input  wire [15:0]   io_writes_0_cmd_payload_mask,
  input  wire [1:0]    io_writes_0_cmd_payload_priority,
  input  wire [7:0]    io_writes_0_cmd_payload_context,
  output wire          io_writes_0_rsp_valid,
  output wire [7:0]    io_writes_0_rsp_payload_context,
  input  wire          io_writes_1_cmd_valid,
  output wire          io_writes_1_cmd_ready,
  input  wire [12:0]   io_writes_1_cmd_payload_address,
  input  wire [127:0]  io_writes_1_cmd_payload_data,
  input  wire [15:0]   io_writes_1_cmd_payload_mask,
  input  wire [1:0]    io_writes_1_cmd_payload_priority,
  input  wire [7:0]    io_writes_1_cmd_payload_context,
  output wire          io_writes_1_rsp_valid,
  output wire [7:0]    io_writes_1_rsp_payload_context,
  input  wire          io_writes_2_cmd_valid,
  output wire          io_writes_2_cmd_ready,
  input  wire [12:0]   io_writes_2_cmd_payload_address,
  input  wire [255:0]  io_writes_2_cmd_payload_data,
  input  wire [31:0]   io_writes_2_cmd_payload_mask,
  input  wire [8:0]    io_writes_2_cmd_payload_context,
  output wire          io_writes_2_rsp_valid,
  output wire [8:0]    io_writes_2_rsp_payload_context,
  input  wire          io_reads_0_cmd_valid,
  output wire          io_reads_0_cmd_ready,
  input  wire [12:0]   io_reads_0_cmd_payload_address,
  input  wire [1:0]    io_reads_0_cmd_payload_priority,
  input  wire [2:0]    io_reads_0_cmd_payload_context,
  output wire          io_reads_0_rsp_valid,
  input  wire          io_reads_0_rsp_ready,
  output wire [127:0]  io_reads_0_rsp_payload_data,
  output wire [15:0]   io_reads_0_rsp_payload_mask,
  output wire [2:0]    io_reads_0_rsp_payload_context,
  input  wire          io_reads_1_cmd_valid,
  output wire          io_reads_1_cmd_ready,
  input  wire [12:0]   io_reads_1_cmd_payload_address,
  input  wire [1:0]    io_reads_1_cmd_payload_priority,
  input  wire [2:0]    io_reads_1_cmd_payload_context,
  output wire          io_reads_1_rsp_valid,
  input  wire          io_reads_1_rsp_ready,
  output wire [127:0]  io_reads_1_rsp_payload_data,
  output wire [15:0]   io_reads_1_rsp_payload_mask,
  output wire [2:0]    io_reads_1_rsp_payload_context,
  input  wire          io_reads_2_cmd_valid,
  output wire          io_reads_2_cmd_ready,
  input  wire [12:0]   io_reads_2_cmd_payload_address,
  input  wire [14:0]   io_reads_2_cmd_payload_context,
  output wire          io_reads_2_rsp_valid,
  input  wire          io_reads_2_rsp_ready,
  output wire [255:0]  io_reads_2_rsp_payload_data,
  output wire [31:0]   io_reads_2_rsp_payload_mask,
  output wire [14:0]   io_reads_2_rsp_payload_context,
  input  wire          clk,
  input  wire          reset
);

  reg        [143:0]  banks_0_ram_spinal_port1;
  reg        [143:0]  banks_1_ram_spinal_port1;
  wire       [143:0]  _zz_banks_0_ram_port;
  wire       [143:0]  _zz_banks_1_ram_port;
  wire       [7:0]    _zz_write_ports_0_priority_value;
  wire       [7:0]    _zz_write_ports_1_priority_value;
  wire       [12:0]   _zz_when_MemoryCore_l136;
  wire       [12:0]   _zz_when_MemoryCore_l136_1;
  wire       [12:0]   _zz_when_MemoryCore_l136_2;
  wire       [12:0]   _zz_when_MemoryCore_l136_3;
  reg        [127:0]  _zz_read_ports_0_buffer_bufferIn_payload_data;
  reg        [15:0]   _zz_read_ports_0_buffer_bufferIn_payload_mask;
  wire       [7:0]    _zz_read_ports_0_priority_value;
  reg        [127:0]  _zz_read_ports_1_buffer_bufferIn_payload_data;
  reg        [15:0]   _zz_read_ports_1_buffer_bufferIn_payload_mask;
  wire       [7:0]    _zz_read_ports_1_priority_value;
  wire       [12:0]   _zz_when_MemoryCore_l221;
  wire       [12:0]   _zz_when_MemoryCore_l221_1;
  wire       [12:0]   _zz_when_MemoryCore_l221_2;
  wire       [12:0]   _zz_when_MemoryCore_l221_3;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 banks_0_write_valid;
  reg        [11:0]   banks_0_write_payload_address;
  reg        [127:0]  banks_0_write_payload_data_data;
  reg        [15:0]   banks_0_write_payload_data_mask;
  wire                banks_0_read_cmd_valid;
  wire       [11:0]   banks_0_read_cmd_payload;
  wire       [127:0]  banks_0_read_rsp_data;
  wire       [15:0]   banks_0_read_rsp_mask;
  wire       [143:0]  _zz_banks_0_read_rsp_data;
  wire                banks_0_writeOr_value_valid;
  wire       [11:0]   banks_0_writeOr_value_payload_address;
  wire       [127:0]  banks_0_writeOr_value_payload_data_data;
  wire       [15:0]   banks_0_writeOr_value_payload_data_mask;
  wire                banks_0_readOr_value_valid;
  wire       [11:0]   banks_0_readOr_value_payload;
  reg                 banks_1_write_valid;
  reg        [11:0]   banks_1_write_payload_address;
  reg        [127:0]  banks_1_write_payload_data_data;
  reg        [15:0]   banks_1_write_payload_data_mask;
  wire                banks_1_read_cmd_valid;
  wire       [11:0]   banks_1_read_cmd_payload;
  wire       [127:0]  banks_1_read_rsp_data;
  wire       [15:0]   banks_1_read_rsp_mask;
  wire       [143:0]  _zz_banks_1_read_rsp_data;
  wire                banks_1_writeOr_value_valid;
  wire       [11:0]   banks_1_writeOr_value_payload_address;
  wire       [127:0]  banks_1_writeOr_value_payload_data_data;
  wire       [15:0]   banks_1_writeOr_value_payload_data_mask;
  wire                banks_1_readOr_value_valid;
  wire       [11:0]   banks_1_readOr_value_payload;
  reg        [7:0]    write_ports_0_priority_value;
  reg        [7:0]    write_ports_1_priority_value;
  wire                write_nodes_0_0_priority;
  wire                write_nodes_0_0_conflict;
  wire                write_nodes_0_1_priority;
  wire                write_nodes_0_1_conflict;
  wire                write_nodes_0_2_priority;
  wire                write_nodes_0_2_conflict;
  wire                write_nodes_1_0_priority;
  wire                write_nodes_1_0_conflict;
  wire                write_nodes_1_1_priority;
  wire                write_nodes_1_1_conflict;
  wire                write_nodes_1_2_priority;
  wire                write_nodes_1_2_conflict;
  wire                write_nodes_2_0_priority;
  wire                write_nodes_2_0_conflict;
  wire                write_nodes_2_1_priority;
  wire                write_nodes_2_1_conflict;
  wire                write_nodes_2_2_priority;
  wire                write_nodes_2_2_conflict;
  wire       [1:0]    write_arbiter_0_losedAgainst;
  reg                 write_arbiter_0_doIt;
  reg                 _zz_banks_0_writeOr_value_valid;
  reg        [11:0]   _zz_banks_0_writeOr_value_valid_1;
  reg        [127:0]  _zz_banks_0_writeOr_value_valid_2;
  reg        [15:0]   _zz_banks_0_writeOr_value_valid_3;
  wire                when_MemoryCore_l136;
  reg                 _zz_banks_1_writeOr_value_valid;
  reg        [11:0]   _zz_banks_1_writeOr_value_valid_1;
  reg        [127:0]  _zz_banks_1_writeOr_value_valid_2;
  reg        [15:0]   _zz_banks_1_writeOr_value_valid_3;
  wire                when_MemoryCore_l136_1;
  reg                 write_arbiter_0_doIt_regNext;
  reg        [7:0]    io_writes_0_cmd_payload_context_regNext;
  wire       [1:0]    write_arbiter_1_losedAgainst;
  reg                 write_arbiter_1_doIt;
  reg                 _zz_banks_0_writeOr_value_valid_4;
  reg        [11:0]   _zz_banks_0_writeOr_value_valid_5;
  reg        [127:0]  _zz_banks_0_writeOr_value_valid_6;
  reg        [15:0]   _zz_banks_0_writeOr_value_valid_7;
  wire                when_MemoryCore_l136_2;
  reg                 _zz_banks_1_writeOr_value_valid_4;
  reg        [11:0]   _zz_banks_1_writeOr_value_valid_5;
  reg        [127:0]  _zz_banks_1_writeOr_value_valid_6;
  reg        [15:0]   _zz_banks_1_writeOr_value_valid_7;
  wire                when_MemoryCore_l136_3;
  reg                 write_arbiter_1_doIt_regNext;
  reg        [7:0]    io_writes_1_cmd_payload_context_regNext;
  wire       [1:0]    write_arbiter_2_losedAgainst;
  reg                 write_arbiter_2_doIt;
  reg                 _zz_banks_0_writeOr_value_valid_8;
  reg        [11:0]   _zz_banks_0_writeOr_value_valid_9;
  reg        [127:0]  _zz_banks_0_writeOr_value_valid_10;
  reg        [15:0]   _zz_banks_0_writeOr_value_valid_11;
  wire                when_MemoryCore_l136_4;
  reg                 _zz_banks_1_writeOr_value_valid_8;
  reg        [11:0]   _zz_banks_1_writeOr_value_valid_9;
  reg        [127:0]  _zz_banks_1_writeOr_value_valid_10;
  reg        [15:0]   _zz_banks_1_writeOr_value_valid_11;
  wire                when_MemoryCore_l136_5;
  reg                 write_arbiter_2_doIt_regNext;
  reg        [8:0]    io_writes_2_cmd_payload_context_regNext;
  wire                read_ports_0_buffer_s0_valid;
  wire       [2:0]    read_ports_0_buffer_s0_payload_context;
  wire       [12:0]   read_ports_0_buffer_s0_payload_address;
  reg                 read_ports_0_buffer_s1_valid;
  reg        [2:0]    read_ports_0_buffer_s1_payload_context;
  reg        [12:0]   read_ports_0_buffer_s1_payload_address;
  wire       [0:0]    read_ports_0_buffer_groupSel;
  wire                read_ports_0_buffer_bufferIn_valid;
  wire                read_ports_0_buffer_bufferIn_ready;
  wire       [127:0]  read_ports_0_buffer_bufferIn_payload_data;
  wire       [15:0]   read_ports_0_buffer_bufferIn_payload_mask;
  wire       [2:0]    read_ports_0_buffer_bufferIn_payload_context;
  wire                read_ports_0_buffer_bufferOut_valid;
  wire                read_ports_0_buffer_bufferOut_ready;
  wire       [127:0]  read_ports_0_buffer_bufferOut_payload_data;
  wire       [15:0]   read_ports_0_buffer_bufferOut_payload_mask;
  wire       [2:0]    read_ports_0_buffer_bufferOut_payload_context;
  reg                 read_ports_0_buffer_bufferIn_rValidN;
  reg        [127:0]  read_ports_0_buffer_bufferIn_rData_data;
  reg        [15:0]   read_ports_0_buffer_bufferIn_rData_mask;
  reg        [2:0]    read_ports_0_buffer_bufferIn_rData_context;
  wire                read_ports_0_buffer_full;
  wire                _zz_io_reads_0_cmd_ready;
  wire                read_ports_0_cmd_valid;
  wire                read_ports_0_cmd_ready;
  wire       [12:0]   read_ports_0_cmd_payload_address;
  wire       [1:0]    read_ports_0_cmd_payload_priority;
  wire       [2:0]    read_ports_0_cmd_payload_context;
  reg        [7:0]    read_ports_0_priority_value;
  wire                read_ports_1_buffer_s0_valid;
  wire       [2:0]    read_ports_1_buffer_s0_payload_context;
  wire       [12:0]   read_ports_1_buffer_s0_payload_address;
  reg                 read_ports_1_buffer_s1_valid;
  reg        [2:0]    read_ports_1_buffer_s1_payload_context;
  reg        [12:0]   read_ports_1_buffer_s1_payload_address;
  wire       [0:0]    read_ports_1_buffer_groupSel;
  wire                read_ports_1_buffer_bufferIn_valid;
  wire                read_ports_1_buffer_bufferIn_ready;
  wire       [127:0]  read_ports_1_buffer_bufferIn_payload_data;
  wire       [15:0]   read_ports_1_buffer_bufferIn_payload_mask;
  wire       [2:0]    read_ports_1_buffer_bufferIn_payload_context;
  wire                read_ports_1_buffer_bufferOut_valid;
  wire                read_ports_1_buffer_bufferOut_ready;
  wire       [127:0]  read_ports_1_buffer_bufferOut_payload_data;
  wire       [15:0]   read_ports_1_buffer_bufferOut_payload_mask;
  wire       [2:0]    read_ports_1_buffer_bufferOut_payload_context;
  reg                 read_ports_1_buffer_bufferIn_rValidN;
  reg        [127:0]  read_ports_1_buffer_bufferIn_rData_data;
  reg        [15:0]   read_ports_1_buffer_bufferIn_rData_mask;
  reg        [2:0]    read_ports_1_buffer_bufferIn_rData_context;
  wire                read_ports_1_buffer_full;
  wire                _zz_io_reads_1_cmd_ready;
  wire                read_ports_1_cmd_valid;
  wire                read_ports_1_cmd_ready;
  wire       [12:0]   read_ports_1_cmd_payload_address;
  wire       [1:0]    read_ports_1_cmd_payload_priority;
  wire       [2:0]    read_ports_1_cmd_payload_context;
  reg        [7:0]    read_ports_1_priority_value;
  wire                read_ports_2_buffer_s0_valid;
  wire       [14:0]   read_ports_2_buffer_s0_payload_context;
  wire       [12:0]   read_ports_2_buffer_s0_payload_address;
  reg                 read_ports_2_buffer_s1_valid;
  reg        [14:0]   read_ports_2_buffer_s1_payload_context;
  reg        [12:0]   read_ports_2_buffer_s1_payload_address;
  wire                read_ports_2_buffer_bufferIn_valid;
  wire                read_ports_2_buffer_bufferIn_ready;
  wire       [255:0]  read_ports_2_buffer_bufferIn_payload_data;
  wire       [31:0]   read_ports_2_buffer_bufferIn_payload_mask;
  wire       [14:0]   read_ports_2_buffer_bufferIn_payload_context;
  wire                read_ports_2_buffer_bufferOut_valid;
  wire                read_ports_2_buffer_bufferOut_ready;
  wire       [255:0]  read_ports_2_buffer_bufferOut_payload_data;
  wire       [31:0]   read_ports_2_buffer_bufferOut_payload_mask;
  wire       [14:0]   read_ports_2_buffer_bufferOut_payload_context;
  reg                 read_ports_2_buffer_bufferIn_rValidN;
  reg        [255:0]  read_ports_2_buffer_bufferIn_rData_data;
  reg        [31:0]   read_ports_2_buffer_bufferIn_rData_mask;
  reg        [14:0]   read_ports_2_buffer_bufferIn_rData_context;
  wire                read_ports_2_buffer_full;
  wire                _zz_io_reads_2_cmd_ready;
  wire                read_ports_2_cmd_valid;
  wire                read_ports_2_cmd_ready;
  wire       [12:0]   read_ports_2_cmd_payload_address;
  wire       [14:0]   read_ports_2_cmd_payload_context;
  wire                read_nodes_0_0_priority;
  wire                read_nodes_0_0_conflict;
  wire                read_nodes_0_1_priority;
  wire                read_nodes_0_1_conflict;
  wire                read_nodes_0_2_priority;
  wire                read_nodes_0_2_conflict;
  wire                read_nodes_1_0_priority;
  wire                read_nodes_1_0_conflict;
  wire                read_nodes_1_1_priority;
  wire                read_nodes_1_1_conflict;
  wire                read_nodes_1_2_priority;
  wire                read_nodes_1_2_conflict;
  wire                read_nodes_2_0_priority;
  wire                read_nodes_2_0_conflict;
  wire                read_nodes_2_1_priority;
  wire                read_nodes_2_1_conflict;
  wire                read_nodes_2_2_priority;
  wire                read_nodes_2_2_conflict;
  wire       [1:0]    read_arbiter_0_losedAgainst;
  wire                read_arbiter_0_doIt;
  reg                 _zz_banks_0_readOr_value_valid;
  reg        [11:0]   _zz_banks_0_readOr_value_valid_1;
  wire                when_MemoryCore_l221;
  reg                 _zz_banks_1_readOr_value_valid;
  reg        [11:0]   _zz_banks_1_readOr_value_valid_1;
  wire                when_MemoryCore_l221_1;
  wire       [1:0]    read_arbiter_1_losedAgainst;
  wire                read_arbiter_1_doIt;
  reg                 _zz_banks_0_readOr_value_valid_2;
  reg        [11:0]   _zz_banks_0_readOr_value_valid_3;
  wire                when_MemoryCore_l221_2;
  reg                 _zz_banks_1_readOr_value_valid_2;
  reg        [11:0]   _zz_banks_1_readOr_value_valid_3;
  wire                when_MemoryCore_l221_3;
  wire       [1:0]    read_arbiter_2_losedAgainst;
  wire                read_arbiter_2_doIt;
  reg                 _zz_banks_0_readOr_value_valid_4;
  reg        [11:0]   _zz_banks_0_readOr_value_valid_5;
  wire                when_MemoryCore_l221_4;
  reg                 _zz_banks_1_readOr_value_valid_4;
  reg        [11:0]   _zz_banks_1_readOr_value_valid_5;
  wire                when_MemoryCore_l221_5;
  reg        [12:0]   initialiser_counter;
  wire                initialiser_done;
  wire                when_MemoryCore_l239;
  wire       [143:0]  _zz_banks_0_write_payload_data_data;
  wire       [143:0]  _zz_banks_1_write_payload_data_data;
  wire       [156:0]  _zz_banks_0_writeOr_value_valid_12;
  wire       [155:0]  _zz_banks_0_writeOr_value_payload_address;
  wire       [143:0]  _zz_banks_0_writeOr_value_payload_data_data;
  wire       [12:0]   _zz_banks_0_readOr_value_valid_6;
  wire       [156:0]  _zz_banks_1_writeOr_value_valid_12;
  wire       [155:0]  _zz_banks_1_writeOr_value_payload_address;
  wire       [143:0]  _zz_banks_1_writeOr_value_payload_data_data;
  wire       [12:0]   _zz_banks_1_readOr_value_valid_6;
  (* ram_style = "block" *) reg [143:0] banks_0_ram [0:4095];
  (* ram_style = "block" *) reg [143:0] banks_1_ram [0:4095];

  assign _zz_write_ports_0_priority_value = {6'd0, io_writes_0_cmd_payload_priority};
  assign _zz_write_ports_1_priority_value = {6'd0, io_writes_1_cmd_payload_priority};
  assign _zz_when_MemoryCore_l136 = (io_writes_0_cmd_payload_address ^ 13'h0);
  assign _zz_when_MemoryCore_l136_1 = (io_writes_0_cmd_payload_address ^ 13'h0001);
  assign _zz_when_MemoryCore_l136_2 = (io_writes_1_cmd_payload_address ^ 13'h0);
  assign _zz_when_MemoryCore_l136_3 = (io_writes_1_cmd_payload_address ^ 13'h0001);
  assign _zz_read_ports_0_priority_value = {6'd0, read_ports_0_cmd_payload_priority};
  assign _zz_read_ports_1_priority_value = {6'd0, read_ports_1_cmd_payload_priority};
  assign _zz_when_MemoryCore_l221 = (read_ports_0_cmd_payload_address ^ 13'h0);
  assign _zz_when_MemoryCore_l221_1 = (read_ports_0_cmd_payload_address ^ 13'h0001);
  assign _zz_when_MemoryCore_l221_2 = (read_ports_1_cmd_payload_address ^ 13'h0);
  assign _zz_when_MemoryCore_l221_3 = (read_ports_1_cmd_payload_address ^ 13'h0001);
  assign _zz_banks_0_ram_port = {banks_0_write_payload_data_mask,banks_0_write_payload_data_data};
  assign _zz_banks_1_ram_port = {banks_1_write_payload_data_mask,banks_1_write_payload_data_data};
  always @(posedge clk) begin
    if(_zz_2) begin
      banks_0_ram[banks_0_write_payload_address] <= _zz_banks_0_ram_port;
    end
  end

  always @(posedge clk) begin
    if(banks_0_read_cmd_valid) begin
      banks_0_ram_spinal_port1 <= banks_0_ram[banks_0_read_cmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      banks_1_ram[banks_1_write_payload_address] <= _zz_banks_1_ram_port;
    end
  end

  always @(posedge clk) begin
    if(banks_1_read_cmd_valid) begin
      banks_1_ram_spinal_port1 <= banks_1_ram[banks_1_read_cmd_payload];
    end
  end

  initial begin
  `ifndef SYNTHESIS
    write_ports_0_priority_value = {$urandom};
    write_ports_1_priority_value = {$urandom};
    read_ports_0_priority_value = {$urandom};
    read_ports_1_priority_value = {$urandom};
  `endif
  end

  always @(*) begin
    case(read_ports_0_buffer_groupSel)
      1'b0 : begin
        _zz_read_ports_0_buffer_bufferIn_payload_data = banks_0_read_rsp_data;
        _zz_read_ports_0_buffer_bufferIn_payload_mask = banks_0_read_rsp_mask;
      end
      default : begin
        _zz_read_ports_0_buffer_bufferIn_payload_data = banks_1_read_rsp_data;
        _zz_read_ports_0_buffer_bufferIn_payload_mask = banks_1_read_rsp_mask;
      end
    endcase
  end

  always @(*) begin
    case(read_ports_1_buffer_groupSel)
      1'b0 : begin
        _zz_read_ports_1_buffer_bufferIn_payload_data = banks_0_read_rsp_data;
        _zz_read_ports_1_buffer_bufferIn_payload_mask = banks_0_read_rsp_mask;
      end
      default : begin
        _zz_read_ports_1_buffer_bufferIn_payload_data = banks_1_read_rsp_data;
        _zz_read_ports_1_buffer_bufferIn_payload_mask = banks_1_read_rsp_mask;
      end
    endcase
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(banks_1_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(banks_0_write_valid) begin
      _zz_2 = 1'b1;
    end
  end

  assign _zz_banks_0_read_rsp_data = banks_0_ram_spinal_port1;
  assign banks_0_read_rsp_data = _zz_banks_0_read_rsp_data[127 : 0];
  assign banks_0_read_rsp_mask = _zz_banks_0_read_rsp_data[143 : 128];
  always @(*) begin
    banks_0_write_valid = banks_0_writeOr_value_valid;
    if(when_MemoryCore_l239) begin
      banks_0_write_valid = 1'b1;
    end
  end

  always @(*) begin
    banks_0_write_payload_address = banks_0_writeOr_value_payload_address;
    if(when_MemoryCore_l239) begin
      banks_0_write_payload_address = initialiser_counter[11:0];
    end
  end

  always @(*) begin
    banks_0_write_payload_data_data = banks_0_writeOr_value_payload_data_data;
    if(when_MemoryCore_l239) begin
      banks_0_write_payload_data_data = _zz_banks_0_write_payload_data_data[127 : 0];
    end
  end

  always @(*) begin
    banks_0_write_payload_data_mask = banks_0_writeOr_value_payload_data_mask;
    if(when_MemoryCore_l239) begin
      banks_0_write_payload_data_mask = _zz_banks_0_write_payload_data_data[143 : 128];
    end
  end

  assign banks_0_read_cmd_valid = banks_0_readOr_value_valid;
  assign banks_0_read_cmd_payload = banks_0_readOr_value_payload;
  assign _zz_banks_1_read_rsp_data = banks_1_ram_spinal_port1;
  assign banks_1_read_rsp_data = _zz_banks_1_read_rsp_data[127 : 0];
  assign banks_1_read_rsp_mask = _zz_banks_1_read_rsp_data[143 : 128];
  always @(*) begin
    banks_1_write_valid = banks_1_writeOr_value_valid;
    if(when_MemoryCore_l239) begin
      banks_1_write_valid = 1'b1;
    end
  end

  always @(*) begin
    banks_1_write_payload_address = banks_1_writeOr_value_payload_address;
    if(when_MemoryCore_l239) begin
      banks_1_write_payload_address = initialiser_counter[11:0];
    end
  end

  always @(*) begin
    banks_1_write_payload_data_data = banks_1_writeOr_value_payload_data_data;
    if(when_MemoryCore_l239) begin
      banks_1_write_payload_data_data = _zz_banks_1_write_payload_data_data[127 : 0];
    end
  end

  always @(*) begin
    banks_1_write_payload_data_mask = banks_1_writeOr_value_payload_data_mask;
    if(when_MemoryCore_l239) begin
      banks_1_write_payload_data_mask = _zz_banks_1_write_payload_data_data[143 : 128];
    end
  end

  assign banks_1_read_cmd_valid = banks_1_readOr_value_valid;
  assign banks_1_read_cmd_payload = banks_1_readOr_value_payload;
  assign write_nodes_0_1_priority = (write_ports_1_priority_value < write_ports_0_priority_value);
  assign write_nodes_1_0_priority = (! write_nodes_0_1_priority);
  assign write_nodes_0_1_conflict = ((io_writes_0_cmd_valid && io_writes_1_cmd_valid) && (((io_writes_0_cmd_payload_address ^ io_writes_1_cmd_payload_address) & 13'h0001) == 13'h0));
  assign write_nodes_1_0_conflict = write_nodes_0_1_conflict;
  assign write_nodes_0_2_priority = 1'b0;
  assign write_nodes_2_0_priority = 1'b1;
  assign write_nodes_0_2_conflict = ((io_writes_0_cmd_valid && io_writes_2_cmd_valid) && (((io_writes_0_cmd_payload_address ^ io_writes_2_cmd_payload_address) & 13'h0) == 13'h0));
  assign write_nodes_2_0_conflict = write_nodes_0_2_conflict;
  assign write_nodes_1_2_priority = 1'b0;
  assign write_nodes_2_1_priority = 1'b1;
  assign write_nodes_1_2_conflict = ((io_writes_1_cmd_valid && io_writes_2_cmd_valid) && (((io_writes_1_cmd_payload_address ^ io_writes_2_cmd_payload_address) & 13'h0) == 13'h0));
  assign write_nodes_2_1_conflict = write_nodes_1_2_conflict;
  assign write_arbiter_0_losedAgainst = {(write_nodes_0_2_conflict && (! write_nodes_0_2_priority)),(write_nodes_0_1_conflict && (! write_nodes_0_1_priority))};
  always @(*) begin
    write_arbiter_0_doIt = (io_writes_0_cmd_valid && (write_arbiter_0_losedAgainst == 2'b00));
    if(when_MemoryCore_l239) begin
      write_arbiter_0_doIt = 1'b0;
    end
  end

  assign when_MemoryCore_l136 = (write_arbiter_0_doIt && (_zz_when_MemoryCore_l136[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l136) begin
      _zz_banks_0_writeOr_value_valid = 1'b1;
    end else begin
      _zz_banks_0_writeOr_value_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136) begin
      _zz_banks_0_writeOr_value_valid_1 = (io_writes_0_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_0_writeOr_value_valid_1 = 12'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136) begin
      _zz_banks_0_writeOr_value_valid_2 = io_writes_0_cmd_payload_data[127 : 0];
    end else begin
      _zz_banks_0_writeOr_value_valid_2 = 128'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136) begin
      _zz_banks_0_writeOr_value_valid_3 = io_writes_0_cmd_payload_mask[15 : 0];
    end else begin
      _zz_banks_0_writeOr_value_valid_3 = 16'h0;
    end
  end

  assign when_MemoryCore_l136_1 = (write_arbiter_0_doIt && (_zz_when_MemoryCore_l136_1[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l136_1) begin
      _zz_banks_1_writeOr_value_valid = 1'b1;
    end else begin
      _zz_banks_1_writeOr_value_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_1) begin
      _zz_banks_1_writeOr_value_valid_1 = (io_writes_0_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_1_writeOr_value_valid_1 = 12'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_1) begin
      _zz_banks_1_writeOr_value_valid_2 = io_writes_0_cmd_payload_data[127 : 0];
    end else begin
      _zz_banks_1_writeOr_value_valid_2 = 128'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_1) begin
      _zz_banks_1_writeOr_value_valid_3 = io_writes_0_cmd_payload_mask[15 : 0];
    end else begin
      _zz_banks_1_writeOr_value_valid_3 = 16'h0;
    end
  end

  assign io_writes_0_cmd_ready = write_arbiter_0_doIt;
  assign io_writes_0_rsp_valid = write_arbiter_0_doIt_regNext;
  assign io_writes_0_rsp_payload_context = io_writes_0_cmd_payload_context_regNext;
  assign write_arbiter_1_losedAgainst = {(write_nodes_1_2_conflict && (! write_nodes_1_2_priority)),(write_nodes_1_0_conflict && (! write_nodes_1_0_priority))};
  always @(*) begin
    write_arbiter_1_doIt = (io_writes_1_cmd_valid && (write_arbiter_1_losedAgainst == 2'b00));
    if(when_MemoryCore_l239) begin
      write_arbiter_1_doIt = 1'b0;
    end
  end

  assign when_MemoryCore_l136_2 = (write_arbiter_1_doIt && (_zz_when_MemoryCore_l136_2[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l136_2) begin
      _zz_banks_0_writeOr_value_valid_4 = 1'b1;
    end else begin
      _zz_banks_0_writeOr_value_valid_4 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_2) begin
      _zz_banks_0_writeOr_value_valid_5 = (io_writes_1_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_0_writeOr_value_valid_5 = 12'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_2) begin
      _zz_banks_0_writeOr_value_valid_6 = io_writes_1_cmd_payload_data[127 : 0];
    end else begin
      _zz_banks_0_writeOr_value_valid_6 = 128'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_2) begin
      _zz_banks_0_writeOr_value_valid_7 = io_writes_1_cmd_payload_mask[15 : 0];
    end else begin
      _zz_banks_0_writeOr_value_valid_7 = 16'h0;
    end
  end

  assign when_MemoryCore_l136_3 = (write_arbiter_1_doIt && (_zz_when_MemoryCore_l136_3[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l136_3) begin
      _zz_banks_1_writeOr_value_valid_4 = 1'b1;
    end else begin
      _zz_banks_1_writeOr_value_valid_4 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_3) begin
      _zz_banks_1_writeOr_value_valid_5 = (io_writes_1_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_1_writeOr_value_valid_5 = 12'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_3) begin
      _zz_banks_1_writeOr_value_valid_6 = io_writes_1_cmd_payload_data[127 : 0];
    end else begin
      _zz_banks_1_writeOr_value_valid_6 = 128'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_3) begin
      _zz_banks_1_writeOr_value_valid_7 = io_writes_1_cmd_payload_mask[15 : 0];
    end else begin
      _zz_banks_1_writeOr_value_valid_7 = 16'h0;
    end
  end

  assign io_writes_1_cmd_ready = write_arbiter_1_doIt;
  assign io_writes_1_rsp_valid = write_arbiter_1_doIt_regNext;
  assign io_writes_1_rsp_payload_context = io_writes_1_cmd_payload_context_regNext;
  assign write_arbiter_2_losedAgainst = {(write_nodes_2_1_conflict && (! write_nodes_2_1_priority)),(write_nodes_2_0_conflict && (! write_nodes_2_0_priority))};
  always @(*) begin
    write_arbiter_2_doIt = (io_writes_2_cmd_valid && (write_arbiter_2_losedAgainst == 2'b00));
    if(when_MemoryCore_l239) begin
      write_arbiter_2_doIt = 1'b0;
    end
  end

  assign when_MemoryCore_l136_4 = (write_arbiter_2_doIt && 1'b1);
  always @(*) begin
    if(when_MemoryCore_l136_4) begin
      _zz_banks_0_writeOr_value_valid_8 = 1'b1;
    end else begin
      _zz_banks_0_writeOr_value_valid_8 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_4) begin
      _zz_banks_0_writeOr_value_valid_9 = (io_writes_2_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_0_writeOr_value_valid_9 = 12'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_4) begin
      _zz_banks_0_writeOr_value_valid_10 = io_writes_2_cmd_payload_data[127 : 0];
    end else begin
      _zz_banks_0_writeOr_value_valid_10 = 128'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_4) begin
      _zz_banks_0_writeOr_value_valid_11 = io_writes_2_cmd_payload_mask[15 : 0];
    end else begin
      _zz_banks_0_writeOr_value_valid_11 = 16'h0;
    end
  end

  assign when_MemoryCore_l136_5 = (write_arbiter_2_doIt && 1'b1);
  always @(*) begin
    if(when_MemoryCore_l136_5) begin
      _zz_banks_1_writeOr_value_valid_8 = 1'b1;
    end else begin
      _zz_banks_1_writeOr_value_valid_8 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_5) begin
      _zz_banks_1_writeOr_value_valid_9 = (io_writes_2_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_1_writeOr_value_valid_9 = 12'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_5) begin
      _zz_banks_1_writeOr_value_valid_10 = io_writes_2_cmd_payload_data[255 : 128];
    end else begin
      _zz_banks_1_writeOr_value_valid_10 = 128'h0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l136_5) begin
      _zz_banks_1_writeOr_value_valid_11 = io_writes_2_cmd_payload_mask[31 : 16];
    end else begin
      _zz_banks_1_writeOr_value_valid_11 = 16'h0;
    end
  end

  assign io_writes_2_cmd_ready = write_arbiter_2_doIt;
  assign io_writes_2_rsp_valid = write_arbiter_2_doIt_regNext;
  assign io_writes_2_rsp_payload_context = io_writes_2_cmd_payload_context_regNext;
  assign read_ports_0_buffer_groupSel = read_ports_0_buffer_s1_payload_address[0 : 0];
  assign read_ports_0_buffer_bufferIn_valid = read_ports_0_buffer_s1_valid;
  assign read_ports_0_buffer_bufferIn_payload_context = read_ports_0_buffer_s1_payload_context;
  assign read_ports_0_buffer_bufferIn_payload_data = _zz_read_ports_0_buffer_bufferIn_payload_data;
  assign read_ports_0_buffer_bufferIn_payload_mask = _zz_read_ports_0_buffer_bufferIn_payload_mask;
  assign read_ports_0_buffer_bufferIn_ready = read_ports_0_buffer_bufferIn_rValidN;
  assign read_ports_0_buffer_bufferOut_valid = (read_ports_0_buffer_bufferIn_valid || (! read_ports_0_buffer_bufferIn_rValidN));
  assign read_ports_0_buffer_bufferOut_payload_data = (read_ports_0_buffer_bufferIn_rValidN ? read_ports_0_buffer_bufferIn_payload_data : read_ports_0_buffer_bufferIn_rData_data);
  assign read_ports_0_buffer_bufferOut_payload_mask = (read_ports_0_buffer_bufferIn_rValidN ? read_ports_0_buffer_bufferIn_payload_mask : read_ports_0_buffer_bufferIn_rData_mask);
  assign read_ports_0_buffer_bufferOut_payload_context = (read_ports_0_buffer_bufferIn_rValidN ? read_ports_0_buffer_bufferIn_payload_context : read_ports_0_buffer_bufferIn_rData_context);
  assign io_reads_0_rsp_valid = read_ports_0_buffer_bufferOut_valid;
  assign read_ports_0_buffer_bufferOut_ready = io_reads_0_rsp_ready;
  assign io_reads_0_rsp_payload_data = read_ports_0_buffer_bufferOut_payload_data;
  assign io_reads_0_rsp_payload_mask = read_ports_0_buffer_bufferOut_payload_mask;
  assign io_reads_0_rsp_payload_context = read_ports_0_buffer_bufferOut_payload_context;
  assign read_ports_0_buffer_full = (read_ports_0_buffer_bufferOut_valid && (! read_ports_0_buffer_bufferOut_ready));
  assign _zz_io_reads_0_cmd_ready = (! read_ports_0_buffer_full);
  assign read_ports_0_cmd_valid = (io_reads_0_cmd_valid && _zz_io_reads_0_cmd_ready);
  assign io_reads_0_cmd_ready = (read_ports_0_cmd_ready && _zz_io_reads_0_cmd_ready);
  assign read_ports_0_cmd_payload_address = io_reads_0_cmd_payload_address;
  assign read_ports_0_cmd_payload_priority = io_reads_0_cmd_payload_priority;
  assign read_ports_0_cmd_payload_context = io_reads_0_cmd_payload_context;
  assign read_ports_1_buffer_groupSel = read_ports_1_buffer_s1_payload_address[0 : 0];
  assign read_ports_1_buffer_bufferIn_valid = read_ports_1_buffer_s1_valid;
  assign read_ports_1_buffer_bufferIn_payload_context = read_ports_1_buffer_s1_payload_context;
  assign read_ports_1_buffer_bufferIn_payload_data = _zz_read_ports_1_buffer_bufferIn_payload_data;
  assign read_ports_1_buffer_bufferIn_payload_mask = _zz_read_ports_1_buffer_bufferIn_payload_mask;
  assign read_ports_1_buffer_bufferIn_ready = read_ports_1_buffer_bufferIn_rValidN;
  assign read_ports_1_buffer_bufferOut_valid = (read_ports_1_buffer_bufferIn_valid || (! read_ports_1_buffer_bufferIn_rValidN));
  assign read_ports_1_buffer_bufferOut_payload_data = (read_ports_1_buffer_bufferIn_rValidN ? read_ports_1_buffer_bufferIn_payload_data : read_ports_1_buffer_bufferIn_rData_data);
  assign read_ports_1_buffer_bufferOut_payload_mask = (read_ports_1_buffer_bufferIn_rValidN ? read_ports_1_buffer_bufferIn_payload_mask : read_ports_1_buffer_bufferIn_rData_mask);
  assign read_ports_1_buffer_bufferOut_payload_context = (read_ports_1_buffer_bufferIn_rValidN ? read_ports_1_buffer_bufferIn_payload_context : read_ports_1_buffer_bufferIn_rData_context);
  assign io_reads_1_rsp_valid = read_ports_1_buffer_bufferOut_valid;
  assign read_ports_1_buffer_bufferOut_ready = io_reads_1_rsp_ready;
  assign io_reads_1_rsp_payload_data = read_ports_1_buffer_bufferOut_payload_data;
  assign io_reads_1_rsp_payload_mask = read_ports_1_buffer_bufferOut_payload_mask;
  assign io_reads_1_rsp_payload_context = read_ports_1_buffer_bufferOut_payload_context;
  assign read_ports_1_buffer_full = (read_ports_1_buffer_bufferOut_valid && (! read_ports_1_buffer_bufferOut_ready));
  assign _zz_io_reads_1_cmd_ready = (! read_ports_1_buffer_full);
  assign read_ports_1_cmd_valid = (io_reads_1_cmd_valid && _zz_io_reads_1_cmd_ready);
  assign io_reads_1_cmd_ready = (read_ports_1_cmd_ready && _zz_io_reads_1_cmd_ready);
  assign read_ports_1_cmd_payload_address = io_reads_1_cmd_payload_address;
  assign read_ports_1_cmd_payload_priority = io_reads_1_cmd_payload_priority;
  assign read_ports_1_cmd_payload_context = io_reads_1_cmd_payload_context;
  assign read_ports_2_buffer_bufferIn_valid = read_ports_2_buffer_s1_valid;
  assign read_ports_2_buffer_bufferIn_payload_context = read_ports_2_buffer_s1_payload_context;
  assign read_ports_2_buffer_bufferIn_payload_data = {banks_1_read_rsp_data,banks_0_read_rsp_data};
  assign read_ports_2_buffer_bufferIn_payload_mask = {banks_1_read_rsp_mask,banks_0_read_rsp_mask};
  assign read_ports_2_buffer_bufferIn_ready = read_ports_2_buffer_bufferIn_rValidN;
  assign read_ports_2_buffer_bufferOut_valid = (read_ports_2_buffer_bufferIn_valid || (! read_ports_2_buffer_bufferIn_rValidN));
  assign read_ports_2_buffer_bufferOut_payload_data = (read_ports_2_buffer_bufferIn_rValidN ? read_ports_2_buffer_bufferIn_payload_data : read_ports_2_buffer_bufferIn_rData_data);
  assign read_ports_2_buffer_bufferOut_payload_mask = (read_ports_2_buffer_bufferIn_rValidN ? read_ports_2_buffer_bufferIn_payload_mask : read_ports_2_buffer_bufferIn_rData_mask);
  assign read_ports_2_buffer_bufferOut_payload_context = (read_ports_2_buffer_bufferIn_rValidN ? read_ports_2_buffer_bufferIn_payload_context : read_ports_2_buffer_bufferIn_rData_context);
  assign io_reads_2_rsp_valid = read_ports_2_buffer_bufferOut_valid;
  assign read_ports_2_buffer_bufferOut_ready = io_reads_2_rsp_ready;
  assign io_reads_2_rsp_payload_data = read_ports_2_buffer_bufferOut_payload_data;
  assign io_reads_2_rsp_payload_mask = read_ports_2_buffer_bufferOut_payload_mask;
  assign io_reads_2_rsp_payload_context = read_ports_2_buffer_bufferOut_payload_context;
  assign read_ports_2_buffer_full = (read_ports_2_buffer_bufferOut_valid && (! read_ports_2_buffer_bufferOut_ready));
  assign _zz_io_reads_2_cmd_ready = (! read_ports_2_buffer_full);
  assign read_ports_2_cmd_valid = (io_reads_2_cmd_valid && _zz_io_reads_2_cmd_ready);
  assign io_reads_2_cmd_ready = (read_ports_2_cmd_ready && _zz_io_reads_2_cmd_ready);
  assign read_ports_2_cmd_payload_address = io_reads_2_cmd_payload_address;
  assign read_ports_2_cmd_payload_context = io_reads_2_cmd_payload_context;
  assign read_nodes_0_1_priority = (read_ports_1_priority_value < read_ports_0_priority_value);
  assign read_nodes_1_0_priority = (! read_nodes_0_1_priority);
  assign read_nodes_0_1_conflict = ((read_ports_0_cmd_valid && read_ports_1_cmd_valid) && (((read_ports_0_cmd_payload_address ^ io_reads_1_cmd_payload_address) & 13'h0001) == 13'h0));
  assign read_nodes_1_0_conflict = read_nodes_0_1_conflict;
  assign read_nodes_0_2_priority = 1'b0;
  assign read_nodes_2_0_priority = 1'b1;
  assign read_nodes_0_2_conflict = ((read_ports_0_cmd_valid && read_ports_2_cmd_valid) && (((read_ports_0_cmd_payload_address ^ io_reads_2_cmd_payload_address) & 13'h0) == 13'h0));
  assign read_nodes_2_0_conflict = read_nodes_0_2_conflict;
  assign read_nodes_1_2_priority = 1'b0;
  assign read_nodes_2_1_priority = 1'b1;
  assign read_nodes_1_2_conflict = ((read_ports_1_cmd_valid && read_ports_2_cmd_valid) && (((read_ports_1_cmd_payload_address ^ io_reads_2_cmd_payload_address) & 13'h0) == 13'h0));
  assign read_nodes_2_1_conflict = read_nodes_1_2_conflict;
  assign read_arbiter_0_losedAgainst = {(read_nodes_0_2_conflict && (! read_nodes_0_2_priority)),(read_nodes_0_1_conflict && (! read_nodes_0_1_priority))};
  assign read_arbiter_0_doIt = (read_ports_0_cmd_valid && (read_arbiter_0_losedAgainst == 2'b00));
  assign when_MemoryCore_l221 = (read_arbiter_0_doIt && (_zz_when_MemoryCore_l221[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l221) begin
      _zz_banks_0_readOr_value_valid = 1'b1;
    end else begin
      _zz_banks_0_readOr_value_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l221) begin
      _zz_banks_0_readOr_value_valid_1 = (read_ports_0_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_0_readOr_value_valid_1 = 12'h0;
    end
  end

  assign when_MemoryCore_l221_1 = (read_arbiter_0_doIt && (_zz_when_MemoryCore_l221_1[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l221_1) begin
      _zz_banks_1_readOr_value_valid = 1'b1;
    end else begin
      _zz_banks_1_readOr_value_valid = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l221_1) begin
      _zz_banks_1_readOr_value_valid_1 = (read_ports_0_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_1_readOr_value_valid_1 = 12'h0;
    end
  end

  assign read_ports_0_cmd_ready = read_arbiter_0_doIt;
  assign read_ports_0_buffer_s0_valid = read_arbiter_0_doIt;
  assign read_ports_0_buffer_s0_payload_context = read_ports_0_cmd_payload_context;
  assign read_ports_0_buffer_s0_payload_address = read_ports_0_cmd_payload_address;
  assign read_arbiter_1_losedAgainst = {(read_nodes_1_2_conflict && (! read_nodes_1_2_priority)),(read_nodes_1_0_conflict && (! read_nodes_1_0_priority))};
  assign read_arbiter_1_doIt = (read_ports_1_cmd_valid && (read_arbiter_1_losedAgainst == 2'b00));
  assign when_MemoryCore_l221_2 = (read_arbiter_1_doIt && (_zz_when_MemoryCore_l221_2[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l221_2) begin
      _zz_banks_0_readOr_value_valid_2 = 1'b1;
    end else begin
      _zz_banks_0_readOr_value_valid_2 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l221_2) begin
      _zz_banks_0_readOr_value_valid_3 = (read_ports_1_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_0_readOr_value_valid_3 = 12'h0;
    end
  end

  assign when_MemoryCore_l221_3 = (read_arbiter_1_doIt && (_zz_when_MemoryCore_l221_3[0 : 0] == 1'b0));
  always @(*) begin
    if(when_MemoryCore_l221_3) begin
      _zz_banks_1_readOr_value_valid_2 = 1'b1;
    end else begin
      _zz_banks_1_readOr_value_valid_2 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l221_3) begin
      _zz_banks_1_readOr_value_valid_3 = (read_ports_1_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_1_readOr_value_valid_3 = 12'h0;
    end
  end

  assign read_ports_1_cmd_ready = read_arbiter_1_doIt;
  assign read_ports_1_buffer_s0_valid = read_arbiter_1_doIt;
  assign read_ports_1_buffer_s0_payload_context = read_ports_1_cmd_payload_context;
  assign read_ports_1_buffer_s0_payload_address = read_ports_1_cmd_payload_address;
  assign read_arbiter_2_losedAgainst = {(read_nodes_2_1_conflict && (! read_nodes_2_1_priority)),(read_nodes_2_0_conflict && (! read_nodes_2_0_priority))};
  assign read_arbiter_2_doIt = (read_ports_2_cmd_valid && (read_arbiter_2_losedAgainst == 2'b00));
  assign when_MemoryCore_l221_4 = (read_arbiter_2_doIt && 1'b1);
  always @(*) begin
    if(when_MemoryCore_l221_4) begin
      _zz_banks_0_readOr_value_valid_4 = 1'b1;
    end else begin
      _zz_banks_0_readOr_value_valid_4 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l221_4) begin
      _zz_banks_0_readOr_value_valid_5 = (read_ports_2_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_0_readOr_value_valid_5 = 12'h0;
    end
  end

  assign when_MemoryCore_l221_5 = (read_arbiter_2_doIt && 1'b1);
  always @(*) begin
    if(when_MemoryCore_l221_5) begin
      _zz_banks_1_readOr_value_valid_4 = 1'b1;
    end else begin
      _zz_banks_1_readOr_value_valid_4 = 1'b0;
    end
  end

  always @(*) begin
    if(when_MemoryCore_l221_5) begin
      _zz_banks_1_readOr_value_valid_5 = (read_ports_2_cmd_payload_address >>> 1'd1);
    end else begin
      _zz_banks_1_readOr_value_valid_5 = 12'h0;
    end
  end

  assign read_ports_2_cmd_ready = read_arbiter_2_doIt;
  assign read_ports_2_buffer_s0_valid = read_arbiter_2_doIt;
  assign read_ports_2_buffer_s0_payload_context = read_ports_2_cmd_payload_context;
  assign read_ports_2_buffer_s0_payload_address = read_ports_2_cmd_payload_address;
  assign initialiser_done = initialiser_counter[12];
  assign when_MemoryCore_l239 = (! initialiser_done);
  assign _zz_banks_0_write_payload_data_data = 144'h0;
  assign _zz_banks_1_write_payload_data_data = 144'h0;
  assign _zz_banks_0_writeOr_value_valid_12 = (({{{_zz_banks_0_writeOr_value_valid_3,_zz_banks_0_writeOr_value_valid_2},_zz_banks_0_writeOr_value_valid_1},_zz_banks_0_writeOr_value_valid} | {{{_zz_banks_0_writeOr_value_valid_7,_zz_banks_0_writeOr_value_valid_6},_zz_banks_0_writeOr_value_valid_5},_zz_banks_0_writeOr_value_valid_4}) | {{{_zz_banks_0_writeOr_value_valid_11,_zz_banks_0_writeOr_value_valid_10},_zz_banks_0_writeOr_value_valid_9},_zz_banks_0_writeOr_value_valid_8});
  assign banks_0_writeOr_value_valid = _zz_banks_0_writeOr_value_valid_12[0];
  assign _zz_banks_0_writeOr_value_payload_address = _zz_banks_0_writeOr_value_valid_12[156 : 1];
  assign banks_0_writeOr_value_payload_address = _zz_banks_0_writeOr_value_payload_address[11 : 0];
  assign _zz_banks_0_writeOr_value_payload_data_data = _zz_banks_0_writeOr_value_payload_address[155 : 12];
  assign banks_0_writeOr_value_payload_data_data = _zz_banks_0_writeOr_value_payload_data_data[127 : 0];
  assign banks_0_writeOr_value_payload_data_mask = _zz_banks_0_writeOr_value_payload_data_data[143 : 128];
  assign _zz_banks_0_readOr_value_valid_6 = (({_zz_banks_0_readOr_value_valid_1,_zz_banks_0_readOr_value_valid} | {_zz_banks_0_readOr_value_valid_3,_zz_banks_0_readOr_value_valid_2}) | {_zz_banks_0_readOr_value_valid_5,_zz_banks_0_readOr_value_valid_4});
  assign banks_0_readOr_value_valid = _zz_banks_0_readOr_value_valid_6[0];
  assign banks_0_readOr_value_payload = _zz_banks_0_readOr_value_valid_6[12 : 1];
  assign _zz_banks_1_writeOr_value_valid_12 = (({{{_zz_banks_1_writeOr_value_valid_3,_zz_banks_1_writeOr_value_valid_2},_zz_banks_1_writeOr_value_valid_1},_zz_banks_1_writeOr_value_valid} | {{{_zz_banks_1_writeOr_value_valid_7,_zz_banks_1_writeOr_value_valid_6},_zz_banks_1_writeOr_value_valid_5},_zz_banks_1_writeOr_value_valid_4}) | {{{_zz_banks_1_writeOr_value_valid_11,_zz_banks_1_writeOr_value_valid_10},_zz_banks_1_writeOr_value_valid_9},_zz_banks_1_writeOr_value_valid_8});
  assign banks_1_writeOr_value_valid = _zz_banks_1_writeOr_value_valid_12[0];
  assign _zz_banks_1_writeOr_value_payload_address = _zz_banks_1_writeOr_value_valid_12[156 : 1];
  assign banks_1_writeOr_value_payload_address = _zz_banks_1_writeOr_value_payload_address[11 : 0];
  assign _zz_banks_1_writeOr_value_payload_data_data = _zz_banks_1_writeOr_value_payload_address[155 : 12];
  assign banks_1_writeOr_value_payload_data_data = _zz_banks_1_writeOr_value_payload_data_data[127 : 0];
  assign banks_1_writeOr_value_payload_data_mask = _zz_banks_1_writeOr_value_payload_data_data[143 : 128];
  assign _zz_banks_1_readOr_value_valid_6 = (({_zz_banks_1_readOr_value_valid_1,_zz_banks_1_readOr_value_valid} | {_zz_banks_1_readOr_value_valid_3,_zz_banks_1_readOr_value_valid_2}) | {_zz_banks_1_readOr_value_valid_5,_zz_banks_1_readOr_value_valid_4});
  assign banks_1_readOr_value_valid = _zz_banks_1_readOr_value_valid_6[0];
  assign banks_1_readOr_value_payload = _zz_banks_1_readOr_value_valid_6[12 : 1];
  always @(posedge clk) begin
    if(io_writes_0_cmd_valid) begin
      write_ports_0_priority_value <= (write_ports_0_priority_value + _zz_write_ports_0_priority_value);
      if(io_writes_0_cmd_ready) begin
        write_ports_0_priority_value <= 8'h0;
      end
    end
    if(io_writes_1_cmd_valid) begin
      write_ports_1_priority_value <= (write_ports_1_priority_value + _zz_write_ports_1_priority_value);
      if(io_writes_1_cmd_ready) begin
        write_ports_1_priority_value <= 8'h0;
      end
    end
    io_writes_0_cmd_payload_context_regNext <= io_writes_0_cmd_payload_context;
    io_writes_1_cmd_payload_context_regNext <= io_writes_1_cmd_payload_context;
    io_writes_2_cmd_payload_context_regNext <= io_writes_2_cmd_payload_context;
    read_ports_0_buffer_s1_payload_context <= read_ports_0_buffer_s0_payload_context;
    read_ports_0_buffer_s1_payload_address <= read_ports_0_buffer_s0_payload_address;
    if(read_ports_0_buffer_bufferIn_ready) begin
      read_ports_0_buffer_bufferIn_rData_data <= read_ports_0_buffer_bufferIn_payload_data;
      read_ports_0_buffer_bufferIn_rData_mask <= read_ports_0_buffer_bufferIn_payload_mask;
      read_ports_0_buffer_bufferIn_rData_context <= read_ports_0_buffer_bufferIn_payload_context;
    end
    if(read_ports_0_cmd_valid) begin
      read_ports_0_priority_value <= (read_ports_0_priority_value + _zz_read_ports_0_priority_value);
      if(read_ports_0_cmd_ready) begin
        read_ports_0_priority_value <= 8'h0;
      end
    end
    read_ports_1_buffer_s1_payload_context <= read_ports_1_buffer_s0_payload_context;
    read_ports_1_buffer_s1_payload_address <= read_ports_1_buffer_s0_payload_address;
    if(read_ports_1_buffer_bufferIn_ready) begin
      read_ports_1_buffer_bufferIn_rData_data <= read_ports_1_buffer_bufferIn_payload_data;
      read_ports_1_buffer_bufferIn_rData_mask <= read_ports_1_buffer_bufferIn_payload_mask;
      read_ports_1_buffer_bufferIn_rData_context <= read_ports_1_buffer_bufferIn_payload_context;
    end
    if(read_ports_1_cmd_valid) begin
      read_ports_1_priority_value <= (read_ports_1_priority_value + _zz_read_ports_1_priority_value);
      if(read_ports_1_cmd_ready) begin
        read_ports_1_priority_value <= 8'h0;
      end
    end
    read_ports_2_buffer_s1_payload_context <= read_ports_2_buffer_s0_payload_context;
    read_ports_2_buffer_s1_payload_address <= read_ports_2_buffer_s0_payload_address;
    if(read_ports_2_buffer_bufferIn_ready) begin
      read_ports_2_buffer_bufferIn_rData_data <= read_ports_2_buffer_bufferIn_payload_data;
      read_ports_2_buffer_bufferIn_rData_mask <= read_ports_2_buffer_bufferIn_payload_mask;
      read_ports_2_buffer_bufferIn_rData_context <= read_ports_2_buffer_bufferIn_payload_context;
    end
  end

  always @(posedge clk) begin
    if(reset) begin
      write_arbiter_0_doIt_regNext <= 1'b0;
      write_arbiter_1_doIt_regNext <= 1'b0;
      write_arbiter_2_doIt_regNext <= 1'b0;
      read_ports_0_buffer_s1_valid <= 1'b0;
      read_ports_0_buffer_bufferIn_rValidN <= 1'b1;
      read_ports_1_buffer_s1_valid <= 1'b0;
      read_ports_1_buffer_bufferIn_rValidN <= 1'b1;
      read_ports_2_buffer_s1_valid <= 1'b0;
      read_ports_2_buffer_bufferIn_rValidN <= 1'b1;
      initialiser_counter <= 13'h0;
    end else begin
      write_arbiter_0_doIt_regNext <= write_arbiter_0_doIt;
      write_arbiter_1_doIt_regNext <= write_arbiter_1_doIt;
      write_arbiter_2_doIt_regNext <= write_arbiter_2_doIt;
      read_ports_0_buffer_s1_valid <= read_ports_0_buffer_s0_valid;
      if(read_ports_0_buffer_bufferIn_valid) begin
        read_ports_0_buffer_bufferIn_rValidN <= 1'b0;
      end
      if(read_ports_0_buffer_bufferOut_ready) begin
        read_ports_0_buffer_bufferIn_rValidN <= 1'b1;
      end
      read_ports_1_buffer_s1_valid <= read_ports_1_buffer_s0_valid;
      if(read_ports_1_buffer_bufferIn_valid) begin
        read_ports_1_buffer_bufferIn_rValidN <= 1'b0;
      end
      if(read_ports_1_buffer_bufferOut_ready) begin
        read_ports_1_buffer_bufferIn_rValidN <= 1'b1;
      end
      read_ports_2_buffer_s1_valid <= read_ports_2_buffer_s0_valid;
      if(read_ports_2_buffer_bufferIn_valid) begin
        read_ports_2_buffer_bufferIn_rValidN <= 1'b0;
      end
      if(read_ports_2_buffer_bufferOut_ready) begin
        read_ports_2_buffer_bufferIn_rValidN <= 1'b1;
      end
      if(when_MemoryCore_l239) begin
        initialiser_counter <= (initialiser_counter + 13'h0001);
      end
    end
  end


endmodule

module EfxDMA_StreamFifo_1 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [15:0]   io_push_payload_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [15:0]   io_pop_payload_context,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [15:0]   logic_ram_spinal_port1;
  wire       [2:0]    _zz_logic_ptr_notPow2_counter;
  wire       [2:0]    _zz_logic_ptr_notPow2_counter_1;
  wire       [0:0]    _zz_logic_ptr_notPow2_counter_2;
  wire       [2:0]    _zz_logic_ptr_notPow2_counter_3;
  wire       [0:0]    _zz_logic_ptr_notPow2_counter_4;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                when_Stream_l1283;
  wire                when_Stream_l1287;
  reg        [2:0]    logic_ptr_notPow2_counter;
  wire                io_push_fire;
  wire                io_pop_fire;
  wire                logic_push_onRam_write_valid;
  wire       [2:0]    logic_push_onRam_write_payload_address;
  wire       [15:0]   logic_push_onRam_write_payload_data_context;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [2:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [2:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [2:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [2:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [15:0]   logic_pop_sync_readPort_rsp_context;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [15:0]   logic_pop_sync_readArbitation_translated_payload_context;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [2:0]    logic_pop_sync_popReg;
  reg [15:0] logic_ram [0:6];

  assign _zz_logic_ptr_notPow2_counter = (logic_ptr_notPow2_counter + _zz_logic_ptr_notPow2_counter_1);
  assign _zz_logic_ptr_notPow2_counter_2 = io_push_fire;
  assign _zz_logic_ptr_notPow2_counter_1 = {2'd0, _zz_logic_ptr_notPow2_counter_2};
  assign _zz_logic_ptr_notPow2_counter_4 = io_pop_fire;
  assign _zz_logic_ptr_notPow2_counter_3 = {2'd0, _zz_logic_ptr_notPow2_counter_4};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= logic_push_onRam_write_payload_data_context;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = ((logic_ptr_push == logic_ptr_popOnIo) && logic_ptr_wentUp);
  assign logic_ptr_empty = ((logic_ptr_push == logic_ptr_pop) && (! logic_ptr_wentUp));
  assign when_Stream_l1283 = (logic_ptr_push == 3'b110);
  assign when_Stream_l1287 = (logic_ptr_pop == 3'b110);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign io_pop_fire = (io_pop_valid && io_pop_ready);
  assign logic_ptr_occupancy = logic_ptr_notPow2_counter;
  assign io_push_ready = (! logic_ptr_full);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push;
  assign logic_push_onRam_write_payload_data_context = io_push_payload_context;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop;
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign logic_pop_sync_readPort_rsp_context = logic_ram_spinal_port1[15 : 0];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_context = logic_pop_sync_readPort_rsp_context;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_context = logic_pop_sync_readArbitation_translated_payload_context;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b111 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
      logic_ptr_notPow2_counter <= 3'b000;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 3'b000;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
        if(when_Stream_l1283) begin
          logic_ptr_push <= 3'b000;
        end
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
        if(when_Stream_l1287) begin
          logic_ptr_pop <= 3'b000;
        end
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
      logic_ptr_notPow2_counter <= (_zz_logic_ptr_notPow2_counter - _zz_logic_ptr_notPow2_counter_3);
      if(io_flush) begin
        logic_ptr_notPow2_counter <= 3'b000;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 3'b000;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module EfxDMA_StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [25:0]   io_push_payload_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [25:0]   io_pop_payload_context,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [25:0]   logic_ram_spinal_port1;
  wire       [2:0]    _zz_logic_ptr_notPow2_counter;
  wire       [2:0]    _zz_logic_ptr_notPow2_counter_1;
  wire       [0:0]    _zz_logic_ptr_notPow2_counter_2;
  wire       [2:0]    _zz_logic_ptr_notPow2_counter_3;
  wire       [0:0]    _zz_logic_ptr_notPow2_counter_4;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                when_Stream_l1283;
  wire                when_Stream_l1287;
  reg        [2:0]    logic_ptr_notPow2_counter;
  wire                io_push_fire;
  wire                io_pop_fire;
  wire                logic_push_onRam_write_valid;
  wire       [2:0]    logic_push_onRam_write_payload_address;
  wire       [25:0]   logic_push_onRam_write_payload_data_context;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [2:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [2:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [2:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [2:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [25:0]   logic_pop_sync_readPort_rsp_context;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [25:0]   logic_pop_sync_readArbitation_translated_payload_context;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [2:0]    logic_pop_sync_popReg;
  reg [25:0] logic_ram [0:6];

  assign _zz_logic_ptr_notPow2_counter = (logic_ptr_notPow2_counter + _zz_logic_ptr_notPow2_counter_1);
  assign _zz_logic_ptr_notPow2_counter_2 = io_push_fire;
  assign _zz_logic_ptr_notPow2_counter_1 = {2'd0, _zz_logic_ptr_notPow2_counter_2};
  assign _zz_logic_ptr_notPow2_counter_4 = io_pop_fire;
  assign _zz_logic_ptr_notPow2_counter_3 = {2'd0, _zz_logic_ptr_notPow2_counter_4};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= logic_push_onRam_write_payload_data_context;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = ((logic_ptr_push == logic_ptr_popOnIo) && logic_ptr_wentUp);
  assign logic_ptr_empty = ((logic_ptr_push == logic_ptr_pop) && (! logic_ptr_wentUp));
  assign when_Stream_l1283 = (logic_ptr_push == 3'b110);
  assign when_Stream_l1287 = (logic_ptr_pop == 3'b110);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign io_pop_fire = (io_pop_valid && io_pop_ready);
  assign logic_ptr_occupancy = logic_ptr_notPow2_counter;
  assign io_push_ready = (! logic_ptr_full);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push;
  assign logic_push_onRam_write_payload_data_context = io_push_payload_context;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop;
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign logic_pop_sync_readPort_rsp_context = logic_ram_spinal_port1[25 : 0];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_context = logic_pop_sync_readPort_rsp_context;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_context = logic_pop_sync_readArbitation_translated_payload_context;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b111 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
      logic_ptr_notPow2_counter <= 3'b000;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 3'b000;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
        if(when_Stream_l1283) begin
          logic_ptr_push <= 3'b000;
        end
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
        if(when_Stream_l1287) begin
          logic_ptr_pop <= 3'b000;
        end
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
      logic_ptr_notPow2_counter <= (_zz_logic_ptr_notPow2_counter - _zz_logic_ptr_notPow2_counter_3);
      if(io_flush) begin
        logic_ptr_notPow2_counter <= 3'b000;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 3'b000;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module EfxDMA_BufferCC_1 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          ctrl_clk,
  input  wire          ctrl_reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge ctrl_clk) begin
    if(ctrl_reset) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module EfxDMA_BufferCC (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          clk,
  input  wire          reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge clk) begin
    if(reset) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule
