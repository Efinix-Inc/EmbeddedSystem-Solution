// Generator : SpinalHDL dev    git head : 81793df2c4f55a20f7eff1130c4bb74a4b11319f
// Component : EfxSapphireSoc
// Git hash  : 7746860cebf18cb019aaaa50cd9888a3b705694d

`timescale 1ns/1ps

module EfxSapphireSoc (
  input  wire          io_systemClk,
  input  wire          io_asyncReset,
  input  wire          io_memoryClk,
  input  wire          io_peripheralClk,
  input  wire          jtagCtrl_tck,
  input  wire          userInterruptA,
  input  wire          userInterruptD,
  input  wire          userInterruptC,
  input  wire          userInterruptB,
  output reg           io_memoryReset,
  output reg           io_peripheralReset,
  output reg           io_systemReset,
  output wire          cpu0_customInstruction_cmd_valid,
  input  wire          cpu0_customInstruction_cmd_ready,
  output wire [9:0]    cpu0_customInstruction_function_id,
  output wire [31:0]   cpu0_customInstruction_inputs_0,
  output wire [31:0]   cpu0_customInstruction_inputs_1,
  input  wire          cpu0_customInstruction_rsp_valid,
  output wire          cpu0_customInstruction_rsp_ready,
  input  wire [31:0]   cpu0_customInstruction_outputs_0,
  output wire          cpu1_customInstruction_cmd_valid,
  input  wire          cpu1_customInstruction_cmd_ready,
  output wire [9:0]    cpu1_customInstruction_function_id,
  output wire [31:0]   cpu1_customInstruction_inputs_0,
  output wire [31:0]   cpu1_customInstruction_inputs_1,
  input  wire          cpu1_customInstruction_rsp_valid,
  output wire          cpu1_customInstruction_rsp_ready,
  input  wire [31:0]   cpu1_customInstruction_outputs_0,
  output wire          io_ddrA_aw_valid,
  input  wire          io_ddrA_aw_ready,
  output wire [31:0]   io_ddrA_aw_payload_addr,
  output wire [7:0]    io_ddrA_aw_payload_id,
  output wire [3:0]    io_ddrA_aw_payload_region,
  output wire [7:0]    io_ddrA_aw_payload_len,
  output wire [2:0]    io_ddrA_aw_payload_size,
  output wire [1:0]    io_ddrA_aw_payload_burst,
  output wire [0:0]    io_ddrA_aw_payload_lock,
  output wire [3:0]    io_ddrA_aw_payload_cache,
  output wire [3:0]    io_ddrA_aw_payload_qos,
  output wire [2:0]    io_ddrA_aw_payload_prot,
  output wire          io_ddrA_w_valid,
  input  wire          io_ddrA_w_ready,
  output wire [127:0]  io_ddrA_w_payload_data,
  output wire [15:0]   io_ddrA_w_payload_strb,
  output wire          io_ddrA_w_payload_last,
  input  wire          io_ddrA_b_valid,
  output reg           io_ddrA_b_ready,
  input  wire [7:0]    io_ddrA_b_payload_id,
  input  wire [1:0]    io_ddrA_b_payload_resp,
  output wire          io_ddrA_ar_valid,
  input  wire          io_ddrA_ar_ready,
  output wire [31:0]   io_ddrA_ar_payload_addr,
  output wire [7:0]    io_ddrA_ar_payload_id,
  output wire [3:0]    io_ddrA_ar_payload_region,
  output wire [7:0]    io_ddrA_ar_payload_len,
  output wire [2:0]    io_ddrA_ar_payload_size,
  output wire [1:0]    io_ddrA_ar_payload_burst,
  output wire [0:0]    io_ddrA_ar_payload_lock,
  output wire [3:0]    io_ddrA_ar_payload_cache,
  output wire [3:0]    io_ddrA_ar_payload_qos,
  output wire [2:0]    io_ddrA_ar_payload_prot,
  input  wire          io_ddrA_r_valid,
  output reg           io_ddrA_r_ready,
  input  wire [127:0]  io_ddrA_r_payload_data,
  input  wire [7:0]    io_ddrA_r_payload_id,
  input  wire [1:0]    io_ddrA_r_payload_resp,
  input  wire          io_ddrA_r_payload_last,
  input  wire          io_ddrMasters_1_aw_valid,
  output wire          io_ddrMasters_1_aw_ready,
  input  wire [31:0]   io_ddrMasters_1_aw_payload_addr,
  input  wire [3:0]    io_ddrMasters_1_aw_payload_id,
  input  wire [3:0]    io_ddrMasters_1_aw_payload_region,
  input  wire [7:0]    io_ddrMasters_1_aw_payload_len,
  input  wire [2:0]    io_ddrMasters_1_aw_payload_size,
  input  wire [1:0]    io_ddrMasters_1_aw_payload_burst,
  input  wire [0:0]    io_ddrMasters_1_aw_payload_lock,
  input  wire [3:0]    io_ddrMasters_1_aw_payload_cache,
  input  wire [3:0]    io_ddrMasters_1_aw_payload_qos,
  input  wire [2:0]    io_ddrMasters_1_aw_payload_prot,
  input  wire          io_ddrMasters_1_w_valid,
  output wire          io_ddrMasters_1_w_ready,
  input  wire [31:0]   io_ddrMasters_1_w_payload_data,
  input  wire [3:0]    io_ddrMasters_1_w_payload_strb,
  input  wire          io_ddrMasters_1_w_payload_last,
  output wire          io_ddrMasters_1_b_valid,
  input  wire          io_ddrMasters_1_b_ready,
  output wire [3:0]    io_ddrMasters_1_b_payload_id,
  output wire [1:0]    io_ddrMasters_1_b_payload_resp,
  input  wire          io_ddrMasters_1_ar_valid,
  output wire          io_ddrMasters_1_ar_ready,
  input  wire [31:0]   io_ddrMasters_1_ar_payload_addr,
  input  wire [3:0]    io_ddrMasters_1_ar_payload_id,
  input  wire [3:0]    io_ddrMasters_1_ar_payload_region,
  input  wire [7:0]    io_ddrMasters_1_ar_payload_len,
  input  wire [2:0]    io_ddrMasters_1_ar_payload_size,
  input  wire [1:0]    io_ddrMasters_1_ar_payload_burst,
  input  wire [0:0]    io_ddrMasters_1_ar_payload_lock,
  input  wire [3:0]    io_ddrMasters_1_ar_payload_cache,
  input  wire [3:0]    io_ddrMasters_1_ar_payload_qos,
  input  wire [2:0]    io_ddrMasters_1_ar_payload_prot,
  output wire          io_ddrMasters_1_r_valid,
  input  wire          io_ddrMasters_1_r_ready,
  output wire [31:0]   io_ddrMasters_1_r_payload_data,
  output wire [3:0]    io_ddrMasters_1_r_payload_id,
  output wire [1:0]    io_ddrMasters_1_r_payload_resp,
  output wire          io_ddrMasters_1_r_payload_last,
  input  wire          io_ddrMasters_1_clk,
  output wire          io_ddrMasters_1_reset,
  input  wire          io_ddrMasters_0_aw_valid,
  output wire          io_ddrMasters_0_aw_ready,
  input  wire [31:0]   io_ddrMasters_0_aw_payload_addr,
  input  wire [3:0]    io_ddrMasters_0_aw_payload_id,
  input  wire [3:0]    io_ddrMasters_0_aw_payload_region,
  input  wire [7:0]    io_ddrMasters_0_aw_payload_len,
  input  wire [2:0]    io_ddrMasters_0_aw_payload_size,
  input  wire [1:0]    io_ddrMasters_0_aw_payload_burst,
  input  wire [0:0]    io_ddrMasters_0_aw_payload_lock,
  input  wire [3:0]    io_ddrMasters_0_aw_payload_cache,
  input  wire [3:0]    io_ddrMasters_0_aw_payload_qos,
  input  wire [2:0]    io_ddrMasters_0_aw_payload_prot,
  input  wire          io_ddrMasters_0_w_valid,
  output wire          io_ddrMasters_0_w_ready,
  input  wire [63:0]   io_ddrMasters_0_w_payload_data,
  input  wire [7:0]    io_ddrMasters_0_w_payload_strb,
  input  wire          io_ddrMasters_0_w_payload_last,
  output wire          io_ddrMasters_0_b_valid,
  input  wire          io_ddrMasters_0_b_ready,
  output wire [3:0]    io_ddrMasters_0_b_payload_id,
  output wire [1:0]    io_ddrMasters_0_b_payload_resp,
  input  wire          io_ddrMasters_0_ar_valid,
  output wire          io_ddrMasters_0_ar_ready,
  input  wire [31:0]   io_ddrMasters_0_ar_payload_addr,
  input  wire [3:0]    io_ddrMasters_0_ar_payload_id,
  input  wire [3:0]    io_ddrMasters_0_ar_payload_region,
  input  wire [7:0]    io_ddrMasters_0_ar_payload_len,
  input  wire [2:0]    io_ddrMasters_0_ar_payload_size,
  input  wire [1:0]    io_ddrMasters_0_ar_payload_burst,
  input  wire [0:0]    io_ddrMasters_0_ar_payload_lock,
  input  wire [3:0]    io_ddrMasters_0_ar_payload_cache,
  input  wire [3:0]    io_ddrMasters_0_ar_payload_qos,
  input  wire [2:0]    io_ddrMasters_0_ar_payload_prot,
  output wire          io_ddrMasters_0_r_valid,
  input  wire          io_ddrMasters_0_r_ready,
  output wire [63:0]   io_ddrMasters_0_r_payload_data,
  output wire [3:0]    io_ddrMasters_0_r_payload_id,
  output wire [1:0]    io_ddrMasters_0_r_payload_resp,
  output wire          io_ddrMasters_0_r_payload_last,
  input  wire          io_ddrMasters_0_clk,
  output wire          io_ddrMasters_0_reset,
  output wire          axiA_awvalid,
  input  wire          axiA_awready,
  output wire [31:0]   axiA_awaddr,
  output wire [7:0]    axiA_awid,
  output wire [3:0]    axiA_awregion,
  output wire [7:0]    axiA_awlen,
  output wire [2:0]    axiA_awsize,
  output wire [1:0]    axiA_awburst,
  output wire [0:0]    axiA_awlock,
  output wire [3:0]    axiA_awcache,
  output wire [3:0]    axiA_awqos,
  output wire [2:0]    axiA_awprot,
  output wire          axiA_wvalid,
  input  wire          axiA_wready,
  output wire [31:0]   axiA_wdata,
  output wire [3:0]    axiA_wstrb,
  output wire          axiA_wlast,
  input  wire          axiA_bvalid,
  output wire          axiA_bready,
  input  wire [7:0]    axiA_bid,
  input  wire [1:0]    axiA_bresp,
  output wire          axiA_arvalid,
  input  wire          axiA_arready,
  output wire [31:0]   axiA_araddr,
  output wire [7:0]    axiA_arid,
  output wire [3:0]    axiA_arregion,
  output wire [7:0]    axiA_arlen,
  output wire [2:0]    axiA_arsize,
  output wire [1:0]    axiA_arburst,
  output wire [0:0]    axiA_arlock,
  output wire [3:0]    axiA_arcache,
  output wire [3:0]    axiA_arqos,
  output wire [2:0]    axiA_arprot,
  input  wire          axiA_rvalid,
  output reg           axiA_rready,
  input  wire [31:0]   axiA_rdata,
  input  wire [7:0]    axiA_rid,
  input  wire [1:0]    axiA_rresp,
  input  wire          axiA_rlast,
  input  wire          axiAInterrupt,
  output wire          system_uart_0_io_txd,
  input  wire          system_uart_0_io_rxd,
  output wire          system_i2c_0_io_sda_write,
  input  wire          system_i2c_0_io_sda_read,
  output wire          system_i2c_0_io_scl_write,
  input  wire          system_i2c_0_io_scl_read,
  output wire          system_i2c_2_io_sda_write,
  input  wire          system_i2c_2_io_sda_read,
  output wire          system_i2c_2_io_scl_write,
  input  wire          system_i2c_2_io_scl_read,
  output wire          system_i2c_1_io_sda_write,
  input  wire          system_i2c_1_io_sda_read,
  output wire          system_i2c_1_io_scl_write,
  input  wire          system_i2c_1_io_scl_read,
  input  wire [3:0]    system_gpio_0_io_read,
  output wire [3:0]    system_gpio_0_io_write,
  output wire [3:0]    system_gpio_0_io_writeEnable,
  output wire [15:0]   io_apbSlave_2_PADDR,
  output wire [0:0]    io_apbSlave_2_PSEL,
  output wire          io_apbSlave_2_PENABLE,
  input  wire          io_apbSlave_2_PREADY,
  output wire          io_apbSlave_2_PWRITE,
  output wire [31:0]   io_apbSlave_2_PWDATA,
  input  wire [31:0]   io_apbSlave_2_PRDATA,
  input  wire          io_apbSlave_2_PSLVERROR,
  output wire [15:0]   io_apbSlave_1_PADDR,
  output wire [0:0]    io_apbSlave_1_PSEL,
  output wire          io_apbSlave_1_PENABLE,
  input  wire          io_apbSlave_1_PREADY,
  output wire          io_apbSlave_1_PWRITE,
  output wire [31:0]   io_apbSlave_1_PWDATA,
  input  wire [31:0]   io_apbSlave_1_PRDATA,
  input  wire          io_apbSlave_1_PSLVERROR,
  output wire [15:0]   io_apbSlave_4_PADDR,
  output wire [0:0]    io_apbSlave_4_PSEL,
  output wire          io_apbSlave_4_PENABLE,
  input  wire          io_apbSlave_4_PREADY,
  output wire          io_apbSlave_4_PWRITE,
  output wire [31:0]   io_apbSlave_4_PWDATA,
  input  wire [31:0]   io_apbSlave_4_PRDATA,
  input  wire          io_apbSlave_4_PSLVERROR,
  output wire [15:0]   io_apbSlave_0_PADDR,
  output wire [0:0]    io_apbSlave_0_PSEL,
  output wire          io_apbSlave_0_PENABLE,
  input  wire          io_apbSlave_0_PREADY,
  output wire          io_apbSlave_0_PWRITE,
  output wire [31:0]   io_apbSlave_0_PWDATA,
  input  wire [31:0]   io_apbSlave_0_PRDATA,
  input  wire          io_apbSlave_0_PSLVERROR,
  output wire [15:0]   io_apbSlave_3_PADDR,
  output wire [0:0]    io_apbSlave_3_PSEL,
  output wire          io_apbSlave_3_PENABLE,
  input  wire          io_apbSlave_3_PREADY,
  output wire          io_apbSlave_3_PWRITE,
  output wire [31:0]   io_apbSlave_3_PWDATA,
  input  wire [31:0]   io_apbSlave_3_PRDATA,
  input  wire          io_apbSlave_3_PSLVERROR,
  output wire [0:0]    system_spi_0_io_sclk_write,
  output wire          system_spi_0_io_data_0_writeEnable,
  input  wire [0:0]    system_spi_0_io_data_0_read,
  output wire [0:0]    system_spi_0_io_data_0_write,
  output wire          system_spi_0_io_data_1_writeEnable,
  input  wire [0:0]    system_spi_0_io_data_1_read,
  output wire [0:0]    system_spi_0_io_data_1_write,
  output wire          system_spi_0_io_data_2_writeEnable,
  input  wire [0:0]    system_spi_0_io_data_2_read,
  output wire [0:0]    system_spi_0_io_data_2_write,
  output wire          system_spi_0_io_data_3_writeEnable,
  input  wire [0:0]    system_spi_0_io_data_3_read,
  output wire [0:0]    system_spi_0_io_data_3_write,
  output wire [0:0]    system_spi_0_io_ss,
  output wire [0:0]    system_spi_1_io_sclk_write,
  output wire          system_spi_1_io_data_0_writeEnable,
  input  wire [0:0]    system_spi_1_io_data_0_read,
  output wire [0:0]    system_spi_1_io_data_0_write,
  output wire          system_spi_1_io_data_1_writeEnable,
  input  wire [0:0]    system_spi_1_io_data_1_read,
  output wire [0:0]    system_spi_1_io_data_1_write,
  output wire          system_spi_1_io_data_2_writeEnable,
  input  wire [0:0]    system_spi_1_io_data_2_read,
  output wire [0:0]    system_spi_1_io_data_2_write,
  output wire          system_spi_1_io_data_3_writeEnable,
  input  wire [0:0]    system_spi_1_io_data_3_read,
  output wire [0:0]    system_spi_1_io_data_3_write,
  output wire [0:0]    system_spi_1_io_ss,
  output wire          system_watchdog_hardPanic,
  input  wire          jtagCtrl_tdi,
  input  wire          jtagCtrl_enable,
  input  wire          jtagCtrl_capture,
  input  wire          jtagCtrl_shift,
  input  wire          jtagCtrl_update,
  input  wire          jtagCtrl_reset,
  output wire          jtagCtrl_tdo
);
  localparam DebugDmToHartOp_DATA = 2'd0;
  localparam DebugDmToHartOp_EXECUTE = 2'd1;
  localparam DebugDmToHartOp_REG_WRITE = 2'd2;
  localparam DebugDmToHartOp_REG_READ = 2'd3;
  localparam FpuOpcode_LOAD = 4'd0;
  localparam FpuOpcode_STORE = 4'd1;
  localparam FpuOpcode_MUL = 4'd2;
  localparam FpuOpcode_ADD = 4'd3;
  localparam FpuOpcode_FMA = 4'd4;
  localparam FpuOpcode_I2F = 4'd5;
  localparam FpuOpcode_F2I = 4'd6;
  localparam FpuOpcode_CMP = 4'd7;
  localparam FpuOpcode_DIV = 4'd8;
  localparam FpuOpcode_SQRT = 4'd9;
  localparam FpuOpcode_MIN_MAX = 4'd10;
  localparam FpuOpcode_SGNJ = 4'd11;
  localparam FpuOpcode_FMV_X_W = 4'd12;
  localparam FpuOpcode_FMV_W_X = 4'd13;
  localparam FpuOpcode_FCLASS = 4'd14;
  localparam FpuOpcode_FCVT_X_X = 4'd15;
  localparam FpuFormat_FLOAT = 1'd0;
  localparam FpuFormat_DOUBLE = 1'd1;
  localparam FpuRoundMode_RNE = 3'd0;
  localparam FpuRoundMode_RTZ = 3'd1;
  localparam FpuRoundMode_RDN = 3'd2;
  localparam FpuRoundMode_RUP = 3'd3;
  localparam FpuRoundMode_RMM = 3'd4;

  wire                system_cores_0_logic_cpu_dBus_rsp_payload_error;
  wire                system_cores_0_logic_cpu_dBus_inv_payload_last;
  wire       [31:0]   system_cores_0_logic_cpu_dBus_inv_payload_fragment_address;
  reg                 system_cores_0_logic_cpu_dBus_ack_ready;
  reg                 system_cores_0_logic_cpu_FpuPlugin_port_commit_ready;
  wire                system_cores_0_logic_cpu_iBus_rsp_payload_error;
  wire                system_cores_1_logic_cpu_dBus_rsp_payload_error;
  wire                system_cores_1_logic_cpu_dBus_inv_payload_last;
  wire       [31:0]   system_cores_1_logic_cpu_dBus_inv_payload_fragment_address;
  reg                 system_cores_1_logic_cpu_dBus_ack_ready;
  reg                 system_cores_1_logic_cpu_FpuPlugin_port_commit_ready;
  wire                system_cores_1_logic_cpu_iBus_rsp_payload_error;
  reg                 system_ddr_ddrLogic_cc_fifo_io_output_cmd_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_ar_valid;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_ar_payload_id;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_ar_payload_id;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_aw_valid;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_aw_payload_id;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_aw_payload_id;
  reg                 system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_ready;
  reg                 system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_ready;
  reg                 system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_ready;
  wire                system_axiA_logic_bmbToAxiBridge_io_output_arw_ready;
  wire                bufferCC_74_io_dataIn;
  wire                bufferCC_75_io_dataIn;
  wire                bufferCC_76_io_dataIn;
  wire                bufferCC_77_io_dataIn;
  wire                io_ddrMasters_1_reset_read_buffer;
  wire                io_ddrMasters_0_reset_read_buffer;
  wire                system_cores_0_logic_cpu_dBus_cmd_valid;
  wire                system_cores_0_logic_cpu_dBus_cmd_payload_wr;
  wire                system_cores_0_logic_cpu_dBus_cmd_payload_uncached;
  wire       [31:0]   system_cores_0_logic_cpu_dBus_cmd_payload_address;
  wire       [63:0]   system_cores_0_logic_cpu_dBus_cmd_payload_data;
  wire       [7:0]    system_cores_0_logic_cpu_dBus_cmd_payload_mask;
  wire       [2:0]    system_cores_0_logic_cpu_dBus_cmd_payload_size;
  wire                system_cores_0_logic_cpu_dBus_cmd_payload_exclusive;
  wire                system_cores_0_logic_cpu_dBus_cmd_payload_last;
  wire                system_cores_0_logic_cpu_dBus_inv_ready;
  wire                system_cores_0_logic_cpu_dBus_ack_valid;
  wire                system_cores_0_logic_cpu_dBus_ack_payload_last;
  wire                system_cores_0_logic_cpu_dBus_ack_payload_fragment_hit;
  wire                system_cores_0_logic_cpu_dBus_sync_ready;
  wire                system_cores_0_logic_cpu_debugBus_halted;
  wire                system_cores_0_logic_cpu_debugBus_running;
  wire                system_cores_0_logic_cpu_debugBus_unavailable;
  wire                system_cores_0_logic_cpu_debugBus_haveReset;
  wire                system_cores_0_logic_cpu_debugBus_exception;
  wire                system_cores_0_logic_cpu_debugBus_commit;
  wire                system_cores_0_logic_cpu_debugBus_ebreak;
  wire                system_cores_0_logic_cpu_debugBus_redo;
  wire                system_cores_0_logic_cpu_debugBus_regSuccess;
  wire                system_cores_0_logic_cpu_debugBus_resume_rsp_valid;
  wire                system_cores_0_logic_cpu_debugBus_hartToDm_valid;
  wire       [3:0]    system_cores_0_logic_cpu_debugBus_hartToDm_payload_address;
  wire       [31:0]   system_cores_0_logic_cpu_debugBus_hartToDm_payload_data;
  wire                system_cores_0_logic_cpu_FpuPlugin_port_cmd_valid;
  wire       [3:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_opcode;
  wire       [1:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_arg;
  wire       [4:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs1;
  wire       [4:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs2;
  wire       [4:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs3;
  wire       [4:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rd;
  wire       [0:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_format;
  wire       [2:0]    system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_roundMode;
  wire                system_cores_0_logic_cpu_FpuPlugin_port_commit_valid;
  wire       [3:0]    system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_opcode;
  wire       [4:0]    system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_rd;
  wire                system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_write;
  wire       [63:0]   system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_value;
  wire                system_cores_0_logic_cpu_FpuPlugin_port_rsp_ready;
  wire                system_cores_0_logic_cpu_CfuPlugin_bus_cmd_valid;
  wire       [9:0]    system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_function_id;
  wire       [31:0]   system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_0;
  wire       [31:0]   system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_1;
  wire                system_cores_0_logic_cpu_CfuPlugin_bus_rsp_ready;
  wire                system_cores_0_logic_cpu_iBus_cmd_valid;
  wire       [31:0]   system_cores_0_logic_cpu_iBus_cmd_payload_address;
  wire       [2:0]    system_cores_0_logic_cpu_iBus_cmd_payload_size;
  wire                system_cores_0_logic_cpu_stoptime;
  wire                system_cores_1_logic_cpu_dBus_cmd_valid;
  wire                system_cores_1_logic_cpu_dBus_cmd_payload_wr;
  wire                system_cores_1_logic_cpu_dBus_cmd_payload_uncached;
  wire       [31:0]   system_cores_1_logic_cpu_dBus_cmd_payload_address;
  wire       [63:0]   system_cores_1_logic_cpu_dBus_cmd_payload_data;
  wire       [7:0]    system_cores_1_logic_cpu_dBus_cmd_payload_mask;
  wire       [2:0]    system_cores_1_logic_cpu_dBus_cmd_payload_size;
  wire                system_cores_1_logic_cpu_dBus_cmd_payload_exclusive;
  wire                system_cores_1_logic_cpu_dBus_cmd_payload_last;
  wire                system_cores_1_logic_cpu_dBus_inv_ready;
  wire                system_cores_1_logic_cpu_dBus_ack_valid;
  wire                system_cores_1_logic_cpu_dBus_ack_payload_last;
  wire                system_cores_1_logic_cpu_dBus_ack_payload_fragment_hit;
  wire                system_cores_1_logic_cpu_dBus_sync_ready;
  wire                system_cores_1_logic_cpu_debugBus_halted;
  wire                system_cores_1_logic_cpu_debugBus_running;
  wire                system_cores_1_logic_cpu_debugBus_unavailable;
  wire                system_cores_1_logic_cpu_debugBus_haveReset;
  wire                system_cores_1_logic_cpu_debugBus_exception;
  wire                system_cores_1_logic_cpu_debugBus_commit;
  wire                system_cores_1_logic_cpu_debugBus_ebreak;
  wire                system_cores_1_logic_cpu_debugBus_redo;
  wire                system_cores_1_logic_cpu_debugBus_regSuccess;
  wire                system_cores_1_logic_cpu_debugBus_resume_rsp_valid;
  wire                system_cores_1_logic_cpu_debugBus_hartToDm_valid;
  wire       [3:0]    system_cores_1_logic_cpu_debugBus_hartToDm_payload_address;
  wire       [31:0]   system_cores_1_logic_cpu_debugBus_hartToDm_payload_data;
  wire                system_cores_1_logic_cpu_FpuPlugin_port_cmd_valid;
  wire       [3:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_opcode;
  wire       [1:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_arg;
  wire       [4:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs1;
  wire       [4:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs2;
  wire       [4:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs3;
  wire       [4:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rd;
  wire       [0:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_format;
  wire       [2:0]    system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_roundMode;
  wire                system_cores_1_logic_cpu_FpuPlugin_port_commit_valid;
  wire       [3:0]    system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_opcode;
  wire       [4:0]    system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_rd;
  wire                system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_write;
  wire       [63:0]   system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_value;
  wire                system_cores_1_logic_cpu_FpuPlugin_port_rsp_ready;
  wire                system_cores_1_logic_cpu_CfuPlugin_bus_cmd_valid;
  wire       [9:0]    system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_function_id;
  wire       [31:0]   system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_0;
  wire       [31:0]   system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_1;
  wire                system_cores_1_logic_cpu_CfuPlugin_bus_rsp_ready;
  wire                system_cores_1_logic_cpu_iBus_cmd_valid;
  wire       [31:0]   system_cores_1_logic_cpu_iBus_cmd_payload_address;
  wire       [2:0]    system_cores_1_logic_cpu_iBus_cmd_payload_size;
  wire                system_cores_1_logic_cpu_stoptime;
  wire                system_fpu_logic_io_port_0_cmd_ready;
  wire                system_fpu_logic_io_port_0_commit_ready;
  wire                system_fpu_logic_io_port_0_rsp_valid;
  wire       [63:0]   system_fpu_logic_io_port_0_rsp_payload_value;
  wire                system_fpu_logic_io_port_0_rsp_payload_NV;
  wire                system_fpu_logic_io_port_0_rsp_payload_NX;
  wire                system_fpu_logic_io_port_0_completion_valid;
  wire                system_fpu_logic_io_port_0_completion_payload_flags_NX;
  wire                system_fpu_logic_io_port_0_completion_payload_flags_UF;
  wire                system_fpu_logic_io_port_0_completion_payload_flags_OF;
  wire                system_fpu_logic_io_port_0_completion_payload_flags_DZ;
  wire                system_fpu_logic_io_port_0_completion_payload_flags_NV;
  wire                system_fpu_logic_io_port_0_completion_payload_written;
  wire                system_fpu_logic_io_port_1_cmd_ready;
  wire                system_fpu_logic_io_port_1_commit_ready;
  wire                system_fpu_logic_io_port_1_rsp_valid;
  wire       [63:0]   system_fpu_logic_io_port_1_rsp_payload_value;
  wire                system_fpu_logic_io_port_1_rsp_payload_NV;
  wire                system_fpu_logic_io_port_1_rsp_payload_NX;
  wire                system_fpu_logic_io_port_1_completion_valid;
  wire                system_fpu_logic_io_port_1_completion_payload_flags_NX;
  wire                system_fpu_logic_io_port_1_completion_payload_flags_UF;
  wire                system_fpu_logic_io_port_1_completion_payload_flags_OF;
  wire                system_fpu_logic_io_port_1_completion_payload_flags_DZ;
  wire                system_fpu_logic_io_port_1_completion_payload_flags_NV;
  wire                system_fpu_logic_io_port_1_completion_payload_written;
  wire                system_riscvJtag_debug_logic_dm_io_ctrl_cmd_ready;
  wire                system_riscvJtag_debug_logic_dm_io_ctrl_rsp_valid;
  wire                system_riscvJtag_debug_logic_dm_io_ctrl_rsp_payload_error;
  wire       [31:0]   system_riscvJtag_debug_logic_dm_io_ctrl_rsp_payload_data;
  wire                system_riscvJtag_debug_logic_dm_io_ndmreset;
  wire                system_riscvJtag_debug_logic_dm_io_harts_0_resume_cmd_valid;
  wire                system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_valid;
  wire       [1:0]    system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_op;
  wire       [4:0]    system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_address;
  wire       [31:0]   system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_data;
  wire       [2:0]    system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_size;
  wire                system_riscvJtag_debug_logic_dm_io_harts_0_haltReq;
  wire                system_riscvJtag_debug_logic_dm_io_harts_0_ackReset;
  wire                system_riscvJtag_debug_logic_dm_io_harts_1_resume_cmd_valid;
  wire                system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_valid;
  wire       [1:0]    system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_op;
  wire       [4:0]    system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_address;
  wire       [31:0]   system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_data;
  wire       [2:0]    system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_size;
  wire                system_riscvJtag_debug_logic_dm_io_harts_1_haltReq;
  wire                system_riscvJtag_debug_logic_dm_io_harts_1_ackReset;
  wire                io_asyncReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire                debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire                peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire                ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire                userInterruptA_buffercc_io_dataOut;
  wire                userInterruptD_buffercc_io_dataOut;
  wire                userInterruptC_buffercc_io_dataOut;
  wire                userInterruptB_buffercc_io_dataOut;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_push_ready;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_valid;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_payload;
  wire       [5:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_occupancy;
  wire       [5:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_availability;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_push_ready;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_valid;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_payload;
  wire       [5:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_occupancy;
  wire       [5:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_availability;
  wire                system_coreStopTime_buffercc_io_dataOut;
  wire                system_riscvJtag_debug_systemReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire                system_riscvJtag_hard_noTap_tunnel_io_instruction_tdo;
  wire                system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_valid;
  wire                system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_write;
  wire       [31:0]   system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_data;
  wire       [6:0]    system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_address;
  wire                system_fabric_iBus_bmb_arbiter_io_inputs_0_cmd_ready;
  wire                system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_valid;
  wire                system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data;
  wire                system_fabric_iBus_bmb_arbiter_io_inputs_1_cmd_ready;
  wire                system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_valid;
  wire                system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data;
  wire                system_fabric_iBus_bmb_arbiter_io_output_cmd_valid;
  wire                system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_length;
  wire                system_fabric_iBus_bmb_arbiter_io_output_rsp_ready;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_input_cmd_ready;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_valid;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_data;
  wire       [4:0]    system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_context;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_input_inv_valid;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_all;
  wire       [31:0]   system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_address;
  wire       [5:0]    system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_length;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_source;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_input_ack_ready;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_input_sync_valid;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_monitor_io_input_sync_payload_source;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_valid;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_mask;
  wire       [43:0]   system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_context;
  wire                system_fabric_invalidationMonitor_logic_monitor_io_output_rsp_ready;
  wire                system_fabric_exclusiveMonitor_logic_io_input_cmd_ready;
  wire                system_fabric_exclusiveMonitor_logic_io_input_rsp_valid;
  wire                system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_opcode;
  wire                system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_context;
  wire                system_fabric_exclusiveMonitor_logic_io_input_inv_valid;
  wire                system_fabric_exclusiveMonitor_logic_io_input_inv_payload_all;
  wire       [31:0]   system_fabric_exclusiveMonitor_logic_io_input_inv_payload_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_logic_io_input_inv_payload_length;
  wire       [0:0]    system_fabric_exclusiveMonitor_logic_io_input_inv_payload_source;
  wire                system_fabric_exclusiveMonitor_logic_io_input_ack_ready;
  wire                system_fabric_exclusiveMonitor_logic_io_input_sync_valid;
  wire       [0:0]    system_fabric_exclusiveMonitor_logic_io_input_sync_payload_source;
  wire                system_fabric_exclusiveMonitor_logic_io_output_cmd_valid;
  wire                system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_mask;
  wire       [4:0]    system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_context;
  wire                system_fabric_exclusiveMonitor_logic_io_output_rsp_ready;
  wire                system_fabric_exclusiveMonitor_logic_io_output_inv_ready;
  wire                system_fabric_exclusiveMonitor_logic_io_output_ack_valid;
  wire                system_fabric_exclusiveMonitor_logic_io_output_sync_ready;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_cmd_ready;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_all;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_length;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_ack_ready;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_sync_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_cmd_ready;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_all;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_length;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_ack_ready;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_sync_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_mask;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_output_rsp_ready;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_output_inv_ready;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_output_ack_valid;
  wire                system_fabric_dBusCoherent_bmb_arbiter_io_output_sync_ready;
  wire                system_fabric_iBus_bmb_decoder_io_input_cmd_ready;
  wire                system_fabric_iBus_bmb_decoder_io_input_rsp_valid;
  wire                system_fabric_iBus_bmb_decoder_io_input_rsp_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_data;
  wire                system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_valid;
  wire                system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_length;
  wire                system_fabric_iBus_bmb_decoder_io_outputs_0_rsp_ready;
  wire                system_bridge_bmb_arbiter_io_inputs_0_cmd_ready;
  wire                system_bridge_bmb_arbiter_io_inputs_0_rsp_valid;
  wire                system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_last;
  wire       [0:0]    system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_context;
  wire                system_bridge_bmb_arbiter_io_inputs_1_cmd_ready;
  wire                system_bridge_bmb_arbiter_io_inputs_1_rsp_valid;
  wire                system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_last;
  wire       [0:0]    system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data;
  wire                system_bridge_bmb_arbiter_io_output_cmd_valid;
  wire                system_bridge_bmb_arbiter_io_output_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_arbiter_io_output_rsp_ready;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_input_cmd_ready;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_valid;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_last;
  wire       [1:0]    system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_opcode;
  wire       [127:0]  system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_data;
  wire       [45:0]   system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_context;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_valid;
  wire       [31:0]   system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_size;
  wire       [3:0]    system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_cache;
  wire       [2:0]    system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_prot;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_write;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_valid;
  wire       [127:0]  system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_strb;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_last;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_output_b_ready;
  wire                system_ddr_ddrLogic_bmbToAxiBridge_io_output_r_ready;
  wire                system_ddr_ddrLogic_cc_fifo_io_input_cmd_ready;
  wire                system_ddr_ddrLogic_cc_fifo_io_input_rsp_valid;
  wire                system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_last;
  wire       [1:0]    system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_opcode;
  wire       [127:0]  system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_data;
  wire       [45:0]   system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_context;
  wire                system_ddr_ddrLogic_cc_fifo_io_output_cmd_valid;
  wire                system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_last;
  wire       [1:0]    system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_length;
  wire       [127:0]  system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_data;
  wire       [15:0]   system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_mask;
  wire       [45:0]   system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_context;
  wire                system_ddr_ddrLogic_cc_fifo_io_output_rsp_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_ar_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_valid;
  wire       [127:0]  system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_data;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_resp;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_last;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_ar_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_valid;
  wire       [127:0]  system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_data;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_resp;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_last;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_ar_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_valid;
  wire       [127:0]  system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_data;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_resp;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_last;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_valid;
  wire       [31:0]   system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_prot;
  wire                system_ddr_ddrLogic_arbiterAxi4Read_io_output_r_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_aw_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_w_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_valid;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_payload_resp;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_aw_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_w_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_valid;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_payload_resp;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_aw_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_w_ready;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_valid;
  wire       [5:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_payload_resp;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_valid;
  wire       [31:0]   system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_prot;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_valid;
  wire       [127:0]  system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_strb;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_last;
  wire                system_ddr_ddrLogic_arbiterAxi4Write_io_output_b_ready;
  wire                ddrCd_logic_outputReset_buffercc_io_dataOut;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_input_ar_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_input_aw_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_input_w_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_valid;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_output_r_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_io_output_b_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_ar_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_aw_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_w_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_valid;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_valid;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_r_ready;
  wire                system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_b_ready;
  wire                ddrCd_logic_outputReset_buffercc_1_io_dataOut;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_input_ar_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_input_aw_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_input_w_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_valid;
  wire       [63:0]   system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_valid;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_valid;
  wire       [63:0]   system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_data;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_output_r_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_io_output_b_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_ar_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_aw_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_w_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_valid;
  wire       [63:0]   system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_valid;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_valid;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_valid;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_r_ready;
  wire                system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_b_ready;
  wire                system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_push_ready;
  wire                system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_valid;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_occupancy;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_availability;
  wire                system_axiA_logic_bmbToAxiBridge_io_input_cmd_ready;
  wire                system_axiA_logic_bmbToAxiBridge_io_input_rsp_valid;
  wire                system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_last;
  wire       [1:0]    system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_data;
  wire       [44:0]   system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_context;
  wire                system_axiA_logic_bmbToAxiBridge_io_output_arw_valid;
  wire       [31:0]   system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_addr;
  wire       [7:0]    system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_len;
  wire       [2:0]    system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_size;
  wire       [3:0]    system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_cache;
  wire       [2:0]    system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_prot;
  wire                system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_write;
  wire                system_axiA_logic_bmbToAxiBridge_io_output_w_valid;
  wire       [31:0]   system_axiA_logic_bmbToAxiBridge_io_output_w_payload_data;
  wire       [3:0]    system_axiA_logic_bmbToAxiBridge_io_output_w_payload_strb;
  wire                system_axiA_logic_bmbToAxiBridge_io_output_w_payload_last;
  wire                system_axiA_logic_bmbToAxiBridge_io_output_b_ready;
  wire                system_axiA_logic_bmbToAxiBridge_io_output_r_ready;
  wire                system_bridge_bmb_decoder_io_input_cmd_ready;
  wire                system_bridge_bmb_decoder_io_input_rsp_valid;
  wire                system_bridge_bmb_decoder_io_input_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_decoder_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_decoder_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_decoder_io_input_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_decoder_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_decoder_io_outputs_0_cmd_valid;
  wire                system_bridge_bmb_decoder_io_outputs_0_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_context;
  wire                system_bridge_bmb_decoder_io_outputs_0_rsp_ready;
  wire                system_bridge_bmb_decoder_io_outputs_1_cmd_valid;
  wire                system_bridge_bmb_decoder_io_outputs_1_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_context;
  wire                system_bridge_bmb_decoder_io_outputs_1_rsp_ready;
  wire                system_bridge_bmb_decoder_io_outputs_2_cmd_valid;
  wire                system_bridge_bmb_decoder_io_outputs_2_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_context;
  wire                system_bridge_bmb_decoder_io_outputs_2_rsp_ready;
  wire                system_bridge_bmb_decoder_io_outputs_3_cmd_valid;
  wire                system_bridge_bmb_decoder_io_outputs_3_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_context;
  wire                system_bridge_bmb_decoder_io_outputs_3_rsp_ready;
  wire                system_bridge_bmb_upSizer_io_input_cmd_ready;
  wire                system_bridge_bmb_upSizer_io_input_rsp_valid;
  wire                system_bridge_bmb_upSizer_io_input_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_upSizer_io_output_cmd_valid;
  wire                system_bridge_bmb_upSizer_io_output_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_length;
  wire       [127:0]  system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_data;
  wire       [15:0]   system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_mask;
  wire       [45:0]   system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_upSizer_io_output_rsp_ready;
  wire                system_bridge_bmb_downSizer_io_input_cmd_ready;
  wire                system_bridge_bmb_downSizer_io_input_rsp_valid;
  wire                system_bridge_bmb_downSizer_io_input_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_downSizer_io_output_cmd_valid;
  wire                system_bridge_bmb_downSizer_io_output_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_length;
  wire       [31:0]   system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_data;
  wire       [3:0]    system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_mask;
  wire       [44:0]   system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_downSizer_io_output_rsp_ready;
  wire                system_bridge_bmb_crossClock_io_input_cmd_ready;
  wire                system_bridge_bmb_crossClock_io_input_rsp_valid;
  wire                system_bridge_bmb_crossClock_io_input_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_data;
  wire       [44:0]   system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_crossClock_io_output_cmd_valid;
  wire                system_bridge_bmb_crossClock_io_output_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_length;
  wire       [31:0]   system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_data;
  wire       [3:0]    system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_mask;
  wire       [44:0]   system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_crossClock_io_output_rsp_ready;
  wire                system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1;
  wire                system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1;
  wire                system_ramA_logic_io_bus_cmd_ready;
  wire                system_ramA_logic_io_bus_rsp_valid;
  wire                system_ramA_logic_io_bus_rsp_payload_last;
  wire       [0:0]    system_ramA_logic_io_bus_rsp_payload_fragment_opcode;
  wire       [63:0]   system_ramA_logic_io_bus_rsp_payload_fragment_data;
  wire       [47:0]   system_ramA_logic_io_bus_rsp_payload_fragment_context;
  wire                system_bridge_bmb_downSizer_1_io_input_cmd_ready;
  wire                system_bridge_bmb_downSizer_1_io_input_rsp_valid;
  wire                system_bridge_bmb_downSizer_1_io_input_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_downSizer_1_io_output_cmd_valid;
  wire                system_bridge_bmb_downSizer_1_io_output_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_length;
  wire       [31:0]   system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_data;
  wire       [3:0]    system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_mask;
  wire       [44:0]   system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_downSizer_1_io_output_rsp_ready;
  wire                system_bridge_bmb_unburstify_io_input_cmd_ready;
  wire                system_bridge_bmb_unburstify_io_input_rsp_valid;
  wire                system_bridge_bmb_unburstify_io_input_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_data;
  wire       [44:0]   system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_unburstify_io_output_cmd_valid;
  wire                system_bridge_bmb_unburstify_io_output_cmd_payload_last;
  wire       [0:0]    system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_address;
  wire       [1:0]    system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_length;
  wire       [31:0]   system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_data;
  wire       [3:0]    system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_mask;
  wire       [48:0]   system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_unburstify_io_output_rsp_ready;
  wire                system_bridge_bmb_crossClock_1_io_input_cmd_ready;
  wire                system_bridge_bmb_crossClock_1_io_input_rsp_valid;
  wire                system_bridge_bmb_crossClock_1_io_input_rsp_payload_last;
  wire       [0:0]    system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_data;
  wire       [48:0]   system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_crossClock_1_io_output_cmd_valid;
  wire                system_bridge_bmb_crossClock_1_io_output_cmd_payload_last;
  wire       [0:0]    system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_address;
  wire       [1:0]    system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_length;
  wire       [31:0]   system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_data;
  wire       [3:0]    system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_mask;
  wire       [48:0]   system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_crossClock_1_io_output_rsp_ready;
  wire                system_bridge_bmb_unburstify_1_io_input_cmd_ready;
  wire                system_bridge_bmb_unburstify_1_io_input_rsp_valid;
  wire                system_bridge_bmb_unburstify_1_io_input_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_context;
  wire                system_bridge_bmb_unburstify_1_io_output_cmd_valid;
  wire                system_bridge_bmb_unburstify_1_io_output_cmd_payload_last;
  wire       [0:0]    system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_address;
  wire       [2:0]    system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_mask;
  wire       [47:0]   system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_context;
  wire                system_bridge_bmb_unburstify_1_io_output_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_input_cmd_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_input_rsp_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_data;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_0_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_1_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_2_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_3_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_4_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_5_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_6_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_7_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_8_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_9_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_10_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_11_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_12_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_13_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_14_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_15_rsp_ready;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_valid;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_decoder_io_outputs_16_rsp_ready;
  wire                system_clint_logic_io_bus_cmd_ready;
  wire                system_clint_logic_io_bus_rsp_valid;
  wire                system_clint_logic_io_bus_rsp_payload_last;
  wire       [0:0]    system_clint_logic_io_bus_rsp_payload_fragment_opcode;
  wire       [31:0]   system_clint_logic_io_bus_rsp_payload_fragment_data;
  wire       [48:0]   system_clint_logic_io_bus_rsp_payload_fragment_context;
  wire       [1:0]    system_clint_logic_io_timerInterrupt;
  wire       [1:0]    system_clint_logic_io_softwareInterrupt;
  wire       [63:0]   system_clint_logic_io_time;
  wire                system_uart_0_io_logic_io_bus_cmd_ready;
  wire                system_uart_0_io_logic_io_bus_rsp_valid;
  wire                system_uart_0_io_logic_io_bus_rsp_payload_last;
  wire       [0:0]    system_uart_0_io_logic_io_bus_rsp_payload_fragment_opcode;
  wire       [31:0]   system_uart_0_io_logic_io_bus_rsp_payload_fragment_data;
  wire       [48:0]   system_uart_0_io_logic_io_bus_rsp_payload_fragment_context;
  wire                system_uart_0_io_logic_io_uart_txd;
  wire                system_uart_0_io_logic_io_interrupt;
  wire                system_spi_0_io_logic_io_ctrl_cmd_ready;
  wire                system_spi_0_io_logic_io_ctrl_rsp_valid;
  wire                system_spi_0_io_logic_io_ctrl_rsp_payload_last;
  wire       [0:0]    system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_data;
  wire       [48:0]   system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_context;
  wire       [0:0]    system_spi_0_io_logic_io_spi_sclk_write;
  wire       [0:0]    system_spi_0_io_logic_io_spi_ss;
  wire       [0:0]    system_spi_0_io_logic_io_spi_data_0_write;
  wire                system_spi_0_io_logic_io_spi_data_0_writeEnable;
  wire       [0:0]    system_spi_0_io_logic_io_spi_data_1_write;
  wire                system_spi_0_io_logic_io_spi_data_1_writeEnable;
  wire       [0:0]    system_spi_0_io_logic_io_spi_data_2_write;
  wire                system_spi_0_io_logic_io_spi_data_2_writeEnable;
  wire       [0:0]    system_spi_0_io_logic_io_spi_data_3_write;
  wire                system_spi_0_io_logic_io_spi_data_3_writeEnable;
  wire                system_spi_0_io_logic_io_interrupt;
  wire                system_spi_1_io_logic_io_ctrl_cmd_ready;
  wire                system_spi_1_io_logic_io_ctrl_rsp_valid;
  wire                system_spi_1_io_logic_io_ctrl_rsp_payload_last;
  wire       [0:0]    system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_data;
  wire       [48:0]   system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_context;
  wire       [0:0]    system_spi_1_io_logic_io_spi_sclk_write;
  wire       [0:0]    system_spi_1_io_logic_io_spi_ss;
  wire       [0:0]    system_spi_1_io_logic_io_spi_data_0_write;
  wire                system_spi_1_io_logic_io_spi_data_0_writeEnable;
  wire       [0:0]    system_spi_1_io_logic_io_spi_data_1_write;
  wire                system_spi_1_io_logic_io_spi_data_1_writeEnable;
  wire       [0:0]    system_spi_1_io_logic_io_spi_data_2_write;
  wire                system_spi_1_io_logic_io_spi_data_2_writeEnable;
  wire       [0:0]    system_spi_1_io_logic_io_spi_data_3_write;
  wire                system_spi_1_io_logic_io_spi_data_3_writeEnable;
  wire                system_spi_1_io_logic_io_interrupt;
  wire                system_i2c_0_io_logic_io_ctrl_cmd_ready;
  wire                system_i2c_0_io_logic_io_ctrl_rsp_valid;
  wire                system_i2c_0_io_logic_io_ctrl_rsp_payload_last;
  wire       [0:0]    system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_data;
  wire       [48:0]   system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_context;
  wire                system_i2c_0_io_logic_io_i2c_scl_write;
  wire                system_i2c_0_io_logic_io_i2c_sda_write;
  wire                system_i2c_0_io_logic_io_interrupt;
  wire                system_i2c_2_io_logic_io_ctrl_cmd_ready;
  wire                system_i2c_2_io_logic_io_ctrl_rsp_valid;
  wire                system_i2c_2_io_logic_io_ctrl_rsp_payload_last;
  wire       [0:0]    system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_data;
  wire       [48:0]   system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_context;
  wire                system_i2c_2_io_logic_io_i2c_scl_write;
  wire                system_i2c_2_io_logic_io_i2c_sda_write;
  wire                system_i2c_2_io_logic_io_interrupt;
  wire                system_i2c_1_io_logic_io_ctrl_cmd_ready;
  wire                system_i2c_1_io_logic_io_ctrl_rsp_valid;
  wire                system_i2c_1_io_logic_io_ctrl_rsp_payload_last;
  wire       [0:0]    system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_data;
  wire       [48:0]   system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_context;
  wire                system_i2c_1_io_logic_io_i2c_scl_write;
  wire                system_i2c_1_io_logic_io_i2c_sda_write;
  wire                system_i2c_1_io_logic_io_interrupt;
  wire                system_userTimer_1_logic_io_ctrl_cmd_ready;
  wire                system_userTimer_1_logic_io_ctrl_rsp_valid;
  wire                system_userTimer_1_logic_io_ctrl_rsp_payload_last;
  wire       [0:0]    system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_data;
  wire       [48:0]   system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_context;
  wire       [0:0]    system_userTimer_1_logic_io_interrupts;
  wire                system_userTimer_0_logic_io_ctrl_cmd_ready;
  wire                system_userTimer_0_logic_io_ctrl_rsp_valid;
  wire                system_userTimer_0_logic_io_ctrl_rsp_payload_last;
  wire       [0:0]    system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_opcode;
  wire       [31:0]   system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_data;
  wire       [48:0]   system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_context;
  wire       [0:0]    system_userTimer_0_logic_io_interrupts;
  wire       [3:0]    system_gpio_0_io_logic_io_gpio_write;
  wire       [3:0]    system_gpio_0_io_logic_io_gpio_writeEnable;
  wire                system_gpio_0_io_logic_io_bus_cmd_ready;
  wire                system_gpio_0_io_logic_io_bus_rsp_valid;
  wire                system_gpio_0_io_logic_io_bus_rsp_payload_last;
  wire       [0:0]    system_gpio_0_io_logic_io_bus_rsp_payload_fragment_opcode;
  wire       [31:0]   system_gpio_0_io_logic_io_bus_rsp_payload_fragment_data;
  wire       [48:0]   system_gpio_0_io_logic_io_bus_rsp_payload_fragment_context;
  wire       [3:0]    system_gpio_0_io_logic_io_interrupt;
  wire                system_watchdog_logic_logic_io_bus_cmd_ready;
  wire                system_watchdog_logic_logic_io_bus_rsp_valid;
  wire                system_watchdog_logic_logic_io_bus_rsp_payload_last;
  wire       [0:0]    system_watchdog_logic_logic_io_bus_rsp_payload_fragment_opcode;
  wire       [31:0]   system_watchdog_logic_logic_io_bus_rsp_payload_fragment_data;
  wire       [48:0]   system_watchdog_logic_logic_io_bus_rsp_payload_fragment_context;
  wire       [1:0]    system_watchdog_logic_logic_io_panics;
  wire                io_apbSlave_2_logic_io_input_cmd_ready;
  wire                io_apbSlave_2_logic_io_input_rsp_valid;
  wire                io_apbSlave_2_logic_io_input_rsp_payload_last;
  wire       [0:0]    io_apbSlave_2_logic_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_2_logic_io_input_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_2_logic_io_input_rsp_payload_fragment_context;
  wire       [15:0]   io_apbSlave_2_logic_io_output_PADDR;
  wire       [0:0]    io_apbSlave_2_logic_io_output_PSEL;
  wire                io_apbSlave_2_logic_io_output_PENABLE;
  wire                io_apbSlave_2_logic_io_output_PWRITE;
  wire       [31:0]   io_apbSlave_2_logic_io_output_PWDATA;
  wire                io_apbSlave_1_logic_io_input_cmd_ready;
  wire                io_apbSlave_1_logic_io_input_rsp_valid;
  wire                io_apbSlave_1_logic_io_input_rsp_payload_last;
  wire       [0:0]    io_apbSlave_1_logic_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_1_logic_io_input_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_1_logic_io_input_rsp_payload_fragment_context;
  wire       [15:0]   io_apbSlave_1_logic_io_output_PADDR;
  wire       [0:0]    io_apbSlave_1_logic_io_output_PSEL;
  wire                io_apbSlave_1_logic_io_output_PENABLE;
  wire                io_apbSlave_1_logic_io_output_PWRITE;
  wire       [31:0]   io_apbSlave_1_logic_io_output_PWDATA;
  wire                io_apbSlave_4_logic_io_input_cmd_ready;
  wire                io_apbSlave_4_logic_io_input_rsp_valid;
  wire                io_apbSlave_4_logic_io_input_rsp_payload_last;
  wire       [0:0]    io_apbSlave_4_logic_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_4_logic_io_input_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_4_logic_io_input_rsp_payload_fragment_context;
  wire       [15:0]   io_apbSlave_4_logic_io_output_PADDR;
  wire       [0:0]    io_apbSlave_4_logic_io_output_PSEL;
  wire                io_apbSlave_4_logic_io_output_PENABLE;
  wire                io_apbSlave_4_logic_io_output_PWRITE;
  wire       [31:0]   io_apbSlave_4_logic_io_output_PWDATA;
  wire                io_apbSlave_0_logic_io_input_cmd_ready;
  wire                io_apbSlave_0_logic_io_input_rsp_valid;
  wire                io_apbSlave_0_logic_io_input_rsp_payload_last;
  wire       [0:0]    io_apbSlave_0_logic_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_0_logic_io_input_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_0_logic_io_input_rsp_payload_fragment_context;
  wire       [15:0]   io_apbSlave_0_logic_io_output_PADDR;
  wire       [0:0]    io_apbSlave_0_logic_io_output_PSEL;
  wire                io_apbSlave_0_logic_io_output_PENABLE;
  wire                io_apbSlave_0_logic_io_output_PWRITE;
  wire       [31:0]   io_apbSlave_0_logic_io_output_PWDATA;
  wire                io_apbSlave_3_logic_io_input_cmd_ready;
  wire                io_apbSlave_3_logic_io_input_rsp_valid;
  wire                io_apbSlave_3_logic_io_input_rsp_payload_last;
  wire       [0:0]    io_apbSlave_3_logic_io_input_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_3_logic_io_input_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_3_logic_io_input_rsp_payload_fragment_context;
  wire       [15:0]   io_apbSlave_3_logic_io_output_PADDR;
  wire       [0:0]    io_apbSlave_3_logic_io_output_PSEL;
  wire                io_apbSlave_3_logic_io_output_PENABLE;
  wire                io_apbSlave_3_logic_io_output_PWRITE;
  wire       [31:0]   io_apbSlave_3_logic_io_output_PWDATA;
  wire                io_time_sync_cc_io_input_ready;
  wire                io_time_sync_cc_io_output_valid;
  wire       [63:0]   io_time_sync_cc_io_output_payload;
  wire                io_time_sync_cc_1_io_input_ready;
  wire                io_time_sync_cc_1_io_output_valid;
  wire       [63:0]   io_time_sync_cc_1_io_output_payload;
  wire                bufferCC_74_io_dataOut;
  wire                bufferCC_75_io_dataOut;
  wire                bufferCC_76_io_dataOut;
  wire                bufferCC_77_io_dataOut;
  wire                system_cores_0_externalInterrupt_plic_target_iep_regNext_buffercc_io_dataOut;
  wire                system_cores_1_externalInterrupt_plic_target_iep_regNext_buffercc_io_dataOut;
  wire       [31:0]   _zz_dBus_inv_payload_fragment_address;
  wire       [5:0]    _zz_dBus_inv_payload_fragment_address_1;
  wire       [31:0]   _zz_dBus_inv_payload_fragment_address_2;
  wire       [5:0]    _zz_dBus_inv_payload_fragment_address_3;
  reg                 system_coreStopTime;
  wire                system_cores_0_debugRiscv_halted;
  wire                system_cores_1_debugRiscv_halted;
  wire                system_riscvJtag_debug_systemReset;
  reg                 debugCd_logic_inputResetTrigger;
  reg                 debugCd_logic_outputResetUnbuffered;
  reg        [11:0]   debugCd_logic_holdingLogic_resetCounter;
  wire                when_ClockDomainGenerator_l222;
  reg                 debugCd_logic_outputReset;
  reg                 ddrCd_logic_inputResetTrigger;
  reg                 ddrCd_logic_outputResetUnbuffered;
  reg        [5:0]    ddrCd_logic_holdingLogic_resetCounter;
  wire                when_ClockDomainGenerator_l222_1;
  reg                 ddrCd_logic_outputReset;
  reg                 peripheralCd_logic_inputResetTrigger;
  reg                 peripheralCd_logic_outputResetUnbuffered;
  reg        [5:0]    peripheralCd_logic_holdingLogic_resetCounter;
  wire                when_ClockDomainGenerator_l222_2;
  reg                 peripheralCd_logic_outputReset;
  wire                io_asyncReset_asyncAssertSyncDeassert;
  wire                debugCd_logic_inputResetAdapter_stuff_syncTrigger;
  wire                debugCd_logic_outputReset_asyncAssertSyncDeassert;
  reg                 systemCd_logic_inputResetTrigger;
  reg                 systemCd_logic_outputResetUnbuffered;
  reg        [5:0]    systemCd_logic_holdingLogic_resetCounter;
  wire                when_ClockDomainGenerator_l222_3;
  reg                 systemCd_logic_outputReset;
  wire                peripheralCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                ddrCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                userInterruptA_interrupt;
  wire                userInterruptD_interrupt;
  wire                userInterruptC_interrupt;
  wire                userInterruptB_interrupt;
  wire       [1:0]    userInterruptA_interrupt_plic_gateway_priority;
  reg                 userInterruptA_interrupt_plic_gateway_ip;
  reg                 userInterruptA_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21;
  wire       [1:0]    userInterruptD_interrupt_plic_gateway_priority;
  reg                 userInterruptD_interrupt_plic_gateway_ip;
  reg                 userInterruptD_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_1;
  wire       [1:0]    userInterruptC_interrupt_plic_gateway_priority;
  reg                 userInterruptC_interrupt_plic_gateway_ip;
  reg                 userInterruptC_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_2;
  wire       [1:0]    userInterruptB_interrupt_plic_gateway_priority;
  reg                 userInterruptB_interrupt_plic_gateway_ip;
  reg                 userInterruptB_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_3;
  wire                system_cores_0_debugRiscv_running;
  wire                system_cores_0_debugRiscv_unavailable;
  wire                system_cores_0_debugRiscv_exception;
  wire                system_cores_0_debugRiscv_commit;
  wire                system_cores_0_debugRiscv_ebreak;
  wire                system_cores_0_debugRiscv_redo;
  wire                system_cores_0_debugRiscv_regSuccess;
  wire                system_cores_0_debugRiscv_ackReset;
  wire                system_cores_0_debugRiscv_haveReset;
  wire                system_cores_0_debugRiscv_resume_cmd_valid;
  wire                system_cores_0_debugRiscv_resume_rsp_valid;
  wire                system_cores_0_debugRiscv_haltReq;
  wire                system_cores_0_debugRiscv_dmToHart_valid;
  wire       [1:0]    system_cores_0_debugRiscv_dmToHart_payload_op;
  wire       [4:0]    system_cores_0_debugRiscv_dmToHart_payload_address;
  wire       [31:0]   system_cores_0_debugRiscv_dmToHart_payload_data;
  wire       [2:0]    system_cores_0_debugRiscv_dmToHart_payload_size;
  wire                system_cores_0_debugRiscv_hartToDm_valid;
  wire       [3:0]    system_cores_0_debugRiscv_hartToDm_payload_address;
  wire       [31:0]   system_cores_0_debugRiscv_hartToDm_payload_data;
  wire                system_cores_0_iBus_cmd_valid;
  wire                system_cores_0_iBus_cmd_ready;
  wire                system_cores_0_iBus_cmd_payload_last;
  wire       [0:0]    system_cores_0_iBus_cmd_payload_fragment_opcode;
  wire       [31:0]   system_cores_0_iBus_cmd_payload_fragment_address;
  wire       [5:0]    system_cores_0_iBus_cmd_payload_fragment_length;
  wire                system_cores_0_iBus_rsp_valid;
  wire                system_cores_0_iBus_rsp_ready;
  wire                system_cores_0_iBus_rsp_payload_last;
  wire       [0:0]    system_cores_0_iBus_rsp_payload_fragment_opcode;
  wire       [63:0]   system_cores_0_iBus_rsp_payload_fragment_data;
  wire                dBus_Bridge_bus_cmd_valid;
  reg                 dBus_Bridge_bus_cmd_ready;
  wire                dBus_Bridge_bus_cmd_payload_last;
  wire       [0:0]    dBus_Bridge_bus_cmd_payload_fragment_opcode;
  wire                dBus_Bridge_bus_cmd_payload_fragment_exclusive;
  wire       [31:0]   dBus_Bridge_bus_cmd_payload_fragment_address;
  wire       [5:0]    dBus_Bridge_bus_cmd_payload_fragment_length;
  wire       [63:0]   dBus_Bridge_bus_cmd_payload_fragment_data;
  wire       [7:0]    dBus_Bridge_bus_cmd_payload_fragment_mask;
  wire       [3:0]    dBus_Bridge_bus_cmd_payload_fragment_context;
  wire                dBus_Bridge_bus_rsp_valid;
  wire                dBus_Bridge_bus_rsp_ready;
  wire                dBus_Bridge_bus_rsp_payload_last;
  wire       [0:0]    dBus_Bridge_bus_rsp_payload_fragment_opcode;
  wire                dBus_Bridge_bus_rsp_payload_fragment_exclusive;
  wire       [63:0]   dBus_Bridge_bus_rsp_payload_fragment_data;
  wire       [3:0]    dBus_Bridge_bus_rsp_payload_fragment_context;
  wire                dBus_Bridge_bus_inv_valid;
  wire                dBus_Bridge_bus_inv_ready;
  wire                dBus_Bridge_bus_inv_payload_all;
  wire       [31:0]   dBus_Bridge_bus_inv_payload_address;
  wire       [5:0]    dBus_Bridge_bus_inv_payload_length;
  wire                dBus_Bridge_bus_ack_valid;
  reg                 dBus_Bridge_bus_ack_ready;
  wire                dBus_Bridge_bus_sync_valid;
  wire                dBus_Bridge_bus_sync_ready;
  reg                 _zz_dBus_cmd_ready;
  wire                dBus_Bridge_withWriteBuffer_buffer_stream_valid;
  wire                dBus_Bridge_withWriteBuffer_buffer_stream_ready;
  reg                 _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid;
  wire                when_Stream_l375;
  reg        [31:0]   dBus_Bridge_withWriteBuffer_buffer_address;
  reg        [5:0]    dBus_Bridge_withWriteBuffer_buffer_length;
  reg                 dBus_Bridge_withWriteBuffer_buffer_write;
  reg                 dBus_Bridge_withWriteBuffer_buffer_exclusive;
  reg        [63:0]   dBus_Bridge_withWriteBuffer_buffer_data;
  reg        [7:0]    dBus_Bridge_withWriteBuffer_buffer_mask;
  reg                 dBus_Bridge_withWriteBuffer_aggregationEnabled;
  reg        [3:0]    dBus_Bridge_withWriteBuffer_aggregationCounter;
  wire                dBus_Bridge_withWriteBuffer_aggregationCounterFull;
  reg        [5:0]    dBus_Bridge_withWriteBuffer_timer;
  wire                dBus_Bridge_withWriteBuffer_timerFull;
  wire                dBus_Bridge_withWriteBuffer_hit;
  wire                dBus_Bridge_withWriteBuffer_canAggregate;
  wire                dBus_Bridge_withWriteBuffer_doFlush;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_busCmdContext_rspCount;
  reg                 dBus_Bridge_withWriteBuffer_halt;
  wire                dBus_cmd_fire;
  wire                when_DataCache_l465;
  wire                dBus_Bridge_bus_cmd_fire;
  wire                when_DataCache_l468;
  wire                when_DataCache_l493;
  wire                when_DataCache_l493_1;
  wire                when_DataCache_l493_2;
  wire                when_DataCache_l493_3;
  wire                when_DataCache_l493_4;
  wire                when_DataCache_l493_5;
  wire                when_DataCache_l493_6;
  wire                when_DataCache_l493_7;
  reg        [5:0]    _zz_dBus_Bridge_withWriteBuffer_buffer_length;
  wire                when_DataCache_l506;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_rspCtx_rspCount;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_valid;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_ready;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_payload;
  wire                when_DataCache_l523;
  wire                io_pop_s2mPipe_valid;
  reg                 io_pop_s2mPipe_ready;
  wire       [3:0]    io_pop_s2mPipe_payload;
  reg                 io_pop_rValidN;
  reg        [3:0]    io_pop_rData;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_valid;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_ready;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_payload;
  reg                 io_pop_s2mPipe_rValid;
  reg        [3:0]    io_pop_s2mPipe_rData;
  wire                when_Stream_l375_1;
  wire                dBus_Bridge_bus_sync_fire;
  wire                when_Stream_l445;
  reg                 dBus_ack_thrown_valid;
  wire                dBus_ack_thrown_ready;
  wire                dBus_ack_thrown_payload_last;
  wire                dBus_ack_thrown_payload_fragment_hit;
  wire                system_cores_1_debugRiscv_running;
  wire                system_cores_1_debugRiscv_unavailable;
  wire                system_cores_1_debugRiscv_exception;
  wire                system_cores_1_debugRiscv_commit;
  wire                system_cores_1_debugRiscv_ebreak;
  wire                system_cores_1_debugRiscv_redo;
  wire                system_cores_1_debugRiscv_regSuccess;
  wire                system_cores_1_debugRiscv_ackReset;
  wire                system_cores_1_debugRiscv_haveReset;
  wire                system_cores_1_debugRiscv_resume_cmd_valid;
  wire                system_cores_1_debugRiscv_resume_rsp_valid;
  wire                system_cores_1_debugRiscv_haltReq;
  wire                system_cores_1_debugRiscv_dmToHart_valid;
  wire       [1:0]    system_cores_1_debugRiscv_dmToHart_payload_op;
  wire       [4:0]    system_cores_1_debugRiscv_dmToHart_payload_address;
  wire       [31:0]   system_cores_1_debugRiscv_dmToHart_payload_data;
  wire       [2:0]    system_cores_1_debugRiscv_dmToHart_payload_size;
  wire                system_cores_1_debugRiscv_hartToDm_valid;
  wire       [3:0]    system_cores_1_debugRiscv_hartToDm_payload_address;
  wire       [31:0]   system_cores_1_debugRiscv_hartToDm_payload_data;
  wire                system_cores_1_iBus_cmd_valid;
  wire                system_cores_1_iBus_cmd_ready;
  wire                system_cores_1_iBus_cmd_payload_last;
  wire       [0:0]    system_cores_1_iBus_cmd_payload_fragment_opcode;
  wire       [31:0]   system_cores_1_iBus_cmd_payload_fragment_address;
  wire       [5:0]    system_cores_1_iBus_cmd_payload_fragment_length;
  wire                system_cores_1_iBus_rsp_valid;
  wire                system_cores_1_iBus_rsp_ready;
  wire                system_cores_1_iBus_rsp_payload_last;
  wire       [0:0]    system_cores_1_iBus_rsp_payload_fragment_opcode;
  wire       [63:0]   system_cores_1_iBus_rsp_payload_fragment_data;
  wire                dBus_Bridge_bus_cmd_valid_1;
  reg                 dBus_Bridge_bus_cmd_ready_1;
  wire                dBus_Bridge_bus_cmd_payload_last_1;
  wire       [0:0]    dBus_Bridge_bus_cmd_payload_fragment_opcode_1;
  wire                dBus_Bridge_bus_cmd_payload_fragment_exclusive_1;
  wire       [31:0]   dBus_Bridge_bus_cmd_payload_fragment_address_1;
  wire       [5:0]    dBus_Bridge_bus_cmd_payload_fragment_length_1;
  wire       [63:0]   dBus_Bridge_bus_cmd_payload_fragment_data_1;
  wire       [7:0]    dBus_Bridge_bus_cmd_payload_fragment_mask_1;
  wire       [3:0]    dBus_Bridge_bus_cmd_payload_fragment_context_1;
  wire                dBus_Bridge_bus_rsp_valid_1;
  wire                dBus_Bridge_bus_rsp_ready_1;
  wire                dBus_Bridge_bus_rsp_payload_last_1;
  wire       [0:0]    dBus_Bridge_bus_rsp_payload_fragment_opcode_1;
  wire                dBus_Bridge_bus_rsp_payload_fragment_exclusive_1;
  wire       [63:0]   dBus_Bridge_bus_rsp_payload_fragment_data_1;
  wire       [3:0]    dBus_Bridge_bus_rsp_payload_fragment_context_1;
  wire                dBus_Bridge_bus_inv_valid_1;
  wire                dBus_Bridge_bus_inv_ready_1;
  wire                dBus_Bridge_bus_inv_payload_all_1;
  wire       [31:0]   dBus_Bridge_bus_inv_payload_address_1;
  wire       [5:0]    dBus_Bridge_bus_inv_payload_length_1;
  wire                dBus_Bridge_bus_ack_valid_1;
  reg                 dBus_Bridge_bus_ack_ready_1;
  wire                dBus_Bridge_bus_sync_valid_1;
  wire                dBus_Bridge_bus_sync_ready_1;
  reg                 _zz_dBus_cmd_ready_1;
  wire                dBus_Bridge_withWriteBuffer_buffer_stream_valid_1;
  wire                dBus_Bridge_withWriteBuffer_buffer_stream_ready_1;
  reg                 _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid_1;
  wire                when_Stream_l375_2;
  reg        [31:0]   dBus_Bridge_withWriteBuffer_buffer_address_1;
  reg        [5:0]    dBus_Bridge_withWriteBuffer_buffer_length_1;
  reg                 dBus_Bridge_withWriteBuffer_buffer_write_1;
  reg                 dBus_Bridge_withWriteBuffer_buffer_exclusive_1;
  reg        [63:0]   dBus_Bridge_withWriteBuffer_buffer_data_1;
  reg        [7:0]    dBus_Bridge_withWriteBuffer_buffer_mask_1;
  reg                 dBus_Bridge_withWriteBuffer_aggregationEnabled_1;
  reg        [3:0]    dBus_Bridge_withWriteBuffer_aggregationCounter_1;
  wire                dBus_Bridge_withWriteBuffer_aggregationCounterFull_1;
  reg        [5:0]    dBus_Bridge_withWriteBuffer_timer_1;
  wire                dBus_Bridge_withWriteBuffer_timerFull_1;
  wire                dBus_Bridge_withWriteBuffer_hit_1;
  wire                dBus_Bridge_withWriteBuffer_canAggregate_1;
  wire                dBus_Bridge_withWriteBuffer_doFlush_1;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_busCmdContext_rspCount_1;
  reg                 dBus_Bridge_withWriteBuffer_halt_1;
  wire                dBus_cmd_fire_1;
  wire                when_DataCache_l465_1;
  wire                dBus_Bridge_bus_cmd_fire_1;
  wire                when_DataCache_l468_1;
  wire                when_DataCache_l493_8;
  wire                when_DataCache_l493_9;
  wire                when_DataCache_l493_10;
  wire                when_DataCache_l493_11;
  wire                when_DataCache_l493_12;
  wire                when_DataCache_l493_13;
  wire                when_DataCache_l493_14;
  wire                when_DataCache_l493_15;
  reg        [5:0]    _zz_dBus_Bridge_withWriteBuffer_buffer_length_1;
  wire                when_DataCache_l506_1;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_rspCtx_rspCount_1;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_valid_1;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_ready_1;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_payload_1;
  wire                when_DataCache_l523_1;
  wire                io_pop_s2mPipe_valid_1;
  reg                 io_pop_s2mPipe_ready_1;
  wire       [3:0]    io_pop_s2mPipe_payload_1;
  reg                 io_pop_rValidN_1;
  reg        [3:0]    io_pop_rData_1;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_valid_1;
  wire                dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_ready_1;
  wire       [3:0]    dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_payload_1;
  reg                 io_pop_s2mPipe_rValid_1;
  reg        [3:0]    io_pop_s2mPipe_rData_1;
  wire                when_Stream_l375_3;
  wire                dBus_Bridge_bus_sync_fire_1;
  wire                when_Stream_l445_1;
  reg                 dBus_ack_thrown_valid_1;
  wire                dBus_ack_thrown_ready_1;
  wire                dBus_ack_thrown_payload_last_1;
  wire                dBus_ack_thrown_payload_fragment_hit_1;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_valid;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_ready;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_length;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_valid;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_data;
  reg                 _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready;
  wire                system_cores_0_iBus_cmd_combStage_valid;
  wire                system_cores_0_iBus_cmd_combStage_ready;
  wire                system_cores_0_iBus_cmd_combStage_payload_last;
  wire       [0:0]    system_cores_0_iBus_cmd_combStage_payload_fragment_opcode;
  wire       [31:0]   system_cores_0_iBus_cmd_combStage_payload_fragment_address;
  wire       [5:0]    system_cores_0_iBus_cmd_combStage_payload_fragment_length;
  wire                _zz_system_cores_0_iBus_rsp_valid;
  reg                 _zz_system_cores_0_iBus_rsp_valid_1;
  reg                 _zz_system_cores_0_iBus_rsp_payload_last;
  reg        [0:0]    _zz_system_cores_0_iBus_rsp_payload_fragment_opcode;
  reg        [63:0]   _zz_system_cores_0_iBus_rsp_payload_fragment_data;
  wire                when_Stream_l375_4;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready;
  wire                system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data;
  reg                 _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready;
  wire                system_cores_1_iBus_cmd_combStage_valid;
  wire                system_cores_1_iBus_cmd_combStage_ready;
  wire                system_cores_1_iBus_cmd_combStage_payload_last;
  wire       [0:0]    system_cores_1_iBus_cmd_combStage_payload_fragment_opcode;
  wire       [31:0]   system_cores_1_iBus_cmd_combStage_payload_fragment_address;
  wire       [5:0]    system_cores_1_iBus_cmd_combStage_payload_fragment_length;
  wire                _zz_system_cores_1_iBus_rsp_valid;
  reg                 _zz_system_cores_1_iBus_rsp_valid_1;
  reg                 _zz_system_cores_1_iBus_rsp_payload_last;
  reg        [0:0]    _zz_system_cores_1_iBus_rsp_payload_fragment_opcode;
  reg        [63:0]   _zz_system_cores_1_iBus_rsp_payload_fragment_data;
  wire                when_Stream_l375_5;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_mask;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_all;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_length;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_ack_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_ack_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready;
  reg                 _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready;
  reg                 _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready;
  wire                dBus_Bridge_bus_cmd_m2sPipe_valid;
  wire                dBus_Bridge_bus_cmd_m2sPipe_ready;
  wire                dBus_Bridge_bus_cmd_m2sPipe_payload_last;
  wire       [0:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_opcode;
  wire                dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_exclusive;
  wire       [31:0]   dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_address;
  wire       [5:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_length;
  wire       [63:0]   dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_data;
  wire       [7:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_mask;
  wire       [3:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_context;
  reg                 dBus_Bridge_bus_cmd_rValid;
  reg                 dBus_Bridge_bus_cmd_rData_last;
  reg        [0:0]    dBus_Bridge_bus_cmd_rData_fragment_opcode;
  reg                 dBus_Bridge_bus_cmd_rData_fragment_exclusive;
  reg        [31:0]   dBus_Bridge_bus_cmd_rData_fragment_address;
  reg        [5:0]    dBus_Bridge_bus_cmd_rData_fragment_length;
  reg        [63:0]   dBus_Bridge_bus_cmd_rData_fragment_data;
  reg        [7:0]    dBus_Bridge_bus_cmd_rData_fragment_mask;
  reg        [3:0]    dBus_Bridge_bus_cmd_rData_fragment_context;
  wire                when_Stream_l375_6;
  wire                _zz_dBus_Bridge_bus_inv_valid;
  reg                 _zz_dBus_Bridge_bus_inv_valid_1;
  reg                 _zz_dBus_Bridge_bus_inv_payload_all;
  reg        [31:0]   _zz_dBus_Bridge_bus_inv_payload_address;
  reg        [5:0]    _zz_dBus_Bridge_bus_inv_payload_length;
  wire                when_Stream_l375_7;
  wire                dBus_Bridge_bus_ack_m2sPipe_valid;
  wire                dBus_Bridge_bus_ack_m2sPipe_ready;
  reg                 dBus_Bridge_bus_ack_rValid;
  wire                when_Stream_l375_8;
  wire                _zz_dBus_Bridge_bus_sync_valid;
  reg                 _zz_dBus_Bridge_bus_sync_valid_1;
  wire                when_Stream_l375_9;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_mask;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_all;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_length;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_ack_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_ack_ready;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_valid;
  wire                system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready;
  reg                 _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready;
  reg                 _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready;
  wire                dBus_Bridge_bus_cmd_m2sPipe_valid_1;
  wire                dBus_Bridge_bus_cmd_m2sPipe_ready_1;
  wire                dBus_Bridge_bus_cmd_m2sPipe_payload_last_1;
  wire       [0:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_opcode_1;
  wire                dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_exclusive_1;
  wire       [31:0]   dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_address_1;
  wire       [5:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_length_1;
  wire       [63:0]   dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_data_1;
  wire       [7:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_mask_1;
  wire       [3:0]    dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_context_1;
  reg                 dBus_Bridge_bus_cmd_rValid_1;
  reg                 dBus_Bridge_bus_cmd_rData_last_1;
  reg        [0:0]    dBus_Bridge_bus_cmd_rData_fragment_opcode_1;
  reg                 dBus_Bridge_bus_cmd_rData_fragment_exclusive_1;
  reg        [31:0]   dBus_Bridge_bus_cmd_rData_fragment_address_1;
  reg        [5:0]    dBus_Bridge_bus_cmd_rData_fragment_length_1;
  reg        [63:0]   dBus_Bridge_bus_cmd_rData_fragment_data_1;
  reg        [7:0]    dBus_Bridge_bus_cmd_rData_fragment_mask_1;
  reg        [3:0]    dBus_Bridge_bus_cmd_rData_fragment_context_1;
  wire                when_Stream_l375_10;
  wire                _zz_dBus_Bridge_bus_inv_valid_2;
  reg                 _zz_dBus_Bridge_bus_inv_valid_3;
  reg                 _zz_dBus_Bridge_bus_inv_payload_all_1;
  reg        [31:0]   _zz_dBus_Bridge_bus_inv_payload_address_1;
  reg        [5:0]    _zz_dBus_Bridge_bus_inv_payload_length_1;
  wire                when_Stream_l375_11;
  wire                dBus_Bridge_bus_ack_m2sPipe_valid_1;
  wire                dBus_Bridge_bus_ack_m2sPipe_ready_1;
  reg                 dBus_Bridge_bus_ack_rValid_1;
  wire                when_Stream_l375_12;
  wire                _zz_dBus_Bridge_bus_sync_valid_2;
  reg                 _zz_dBus_Bridge_bus_sync_valid_3;
  wire                when_Stream_l375_13;
  wire                system_peripheralStopTime;
  wire                FpuPlugin_port_commit_m2sPipe_valid;
  wire                FpuPlugin_port_commit_m2sPipe_ready;
  wire       [3:0]    FpuPlugin_port_commit_m2sPipe_payload_opcode;
  wire       [4:0]    FpuPlugin_port_commit_m2sPipe_payload_rd;
  wire                FpuPlugin_port_commit_m2sPipe_payload_write;
  wire       [63:0]   FpuPlugin_port_commit_m2sPipe_payload_value;
  reg                 FpuPlugin_port_commit_rValid;
  reg        [3:0]    FpuPlugin_port_commit_rData_opcode;
  reg        [4:0]    FpuPlugin_port_commit_rData_rd;
  reg                 FpuPlugin_port_commit_rData_write;
  reg        [63:0]   FpuPlugin_port_commit_rData_value;
  wire                when_Stream_l375_14;
  reg                 io_port_0_completion_regNext_valid;
  reg                 io_port_0_completion_regNext_payload_flags_NX;
  reg                 io_port_0_completion_regNext_payload_flags_UF;
  reg                 io_port_0_completion_regNext_payload_flags_OF;
  reg                 io_port_0_completion_regNext_payload_flags_DZ;
  reg                 io_port_0_completion_regNext_payload_flags_NV;
  reg                 io_port_0_completion_regNext_payload_written;
  wire                io_port_0_rsp_s2mPipe_valid;
  wire                io_port_0_rsp_s2mPipe_ready;
  wire       [63:0]   io_port_0_rsp_s2mPipe_payload_value;
  wire                io_port_0_rsp_s2mPipe_payload_NV;
  wire                io_port_0_rsp_s2mPipe_payload_NX;
  reg                 io_port_0_rsp_rValidN;
  reg        [63:0]   io_port_0_rsp_rData_value;
  reg                 io_port_0_rsp_rData_NV;
  reg                 io_port_0_rsp_rData_NX;
  wire                FpuPlugin_port_commit_m2sPipe_valid_1;
  wire                FpuPlugin_port_commit_m2sPipe_ready_1;
  wire       [3:0]    FpuPlugin_port_commit_m2sPipe_payload_opcode_1;
  wire       [4:0]    FpuPlugin_port_commit_m2sPipe_payload_rd_1;
  wire                FpuPlugin_port_commit_m2sPipe_payload_write_1;
  wire       [63:0]   FpuPlugin_port_commit_m2sPipe_payload_value_1;
  reg                 FpuPlugin_port_commit_rValid_1;
  reg        [3:0]    FpuPlugin_port_commit_rData_opcode_1;
  reg        [4:0]    FpuPlugin_port_commit_rData_rd_1;
  reg                 FpuPlugin_port_commit_rData_write_1;
  reg        [63:0]   FpuPlugin_port_commit_rData_value_1;
  wire                when_Stream_l375_15;
  reg                 io_port_1_completion_regNext_valid;
  reg                 io_port_1_completion_regNext_payload_flags_NX;
  reg                 io_port_1_completion_regNext_payload_flags_UF;
  reg                 io_port_1_completion_regNext_payload_flags_OF;
  reg                 io_port_1_completion_regNext_payload_flags_DZ;
  reg                 io_port_1_completion_regNext_payload_flags_NV;
  reg                 io_port_1_completion_regNext_payload_written;
  wire                io_port_1_rsp_s2mPipe_valid;
  wire                io_port_1_rsp_s2mPipe_ready;
  wire       [63:0]   io_port_1_rsp_s2mPipe_payload_value;
  wire                io_port_1_rsp_s2mPipe_payload_NV;
  wire                io_port_1_rsp_s2mPipe_payload_NX;
  reg                 io_port_1_rsp_rValidN;
  reg        [63:0]   io_port_1_rsp_rData_value;
  reg                 io_port_1_rsp_rData_NV;
  reg                 io_port_1_rsp_rData_NX;
  reg                 io_harts_0_dmToHart_regNext_valid;
  reg        [1:0]    io_harts_0_dmToHart_regNext_payload_op;
  reg        [4:0]    io_harts_0_dmToHart_regNext_payload_address;
  reg        [31:0]   io_harts_0_dmToHart_regNext_payload_data;
  reg        [2:0]    io_harts_0_dmToHart_regNext_payload_size;
  reg                 io_harts_1_dmToHart_regNext_valid;
  reg        [1:0]    io_harts_1_dmToHart_regNext_payload_op;
  reg        [4:0]    io_harts_1_dmToHart_regNext_payload_address;
  reg        [31:0]   io_harts_1_dmToHart_regNext_payload_data;
  reg        [2:0]    io_harts_1_dmToHart_regNext_payload_size;
  reg                 _zz_1;
  wire                system_riscvJtag_debug_systemReset_asyncAssertSyncDeassert;
  wire                system_fabric_iBus_bmb_cmd_valid;
  reg                 system_fabric_iBus_bmb_cmd_ready;
  wire                system_fabric_iBus_bmb_cmd_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_iBus_bmb_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_iBus_bmb_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_iBus_bmb_cmd_payload_fragment_length;
  wire                system_fabric_iBus_bmb_rsp_valid;
  wire                system_fabric_iBus_bmb_rsp_ready;
  wire                system_fabric_iBus_bmb_rsp_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_iBus_bmb_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_iBus_bmb_rsp_payload_fragment_data;
  wire                system_fabric_invalidationMonitor_logic_input_cmd_valid;
  wire                system_fabric_invalidationMonitor_logic_input_cmd_ready;
  wire                system_fabric_invalidationMonitor_logic_input_cmd_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_mask;
  wire       [4:0]    system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_context;
  wire                system_fabric_invalidationMonitor_logic_input_rsp_valid;
  wire                system_fabric_invalidationMonitor_logic_input_rsp_ready;
  wire                system_fabric_invalidationMonitor_logic_input_rsp_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_data;
  wire       [4:0]    system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_context;
  wire                system_fabric_invalidationMonitor_logic_input_inv_valid;
  wire                system_fabric_invalidationMonitor_logic_input_inv_ready;
  wire                system_fabric_invalidationMonitor_logic_input_inv_payload_all;
  wire       [31:0]   system_fabric_invalidationMonitor_logic_input_inv_payload_address;
  wire       [5:0]    system_fabric_invalidationMonitor_logic_input_inv_payload_length;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_input_inv_payload_source;
  wire                system_fabric_invalidationMonitor_logic_input_ack_valid;
  wire                system_fabric_invalidationMonitor_logic_input_ack_ready;
  wire                system_fabric_invalidationMonitor_logic_input_sync_valid;
  wire                system_fabric_invalidationMonitor_logic_input_sync_ready;
  wire       [0:0]    system_fabric_invalidationMonitor_logic_input_sync_payload_source;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [4:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [4:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_ready;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all;
  wire       [31:0]   system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address;
  wire       [5:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_valid;
  reg                 system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_valid;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_ready;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_payload_source;
  wire                _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid;
  wire                _zz_system_fabric_invalidationMonitor_logic_input_inv_ready;
  wire                _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all;
  wire       [31:0]   _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address;
  wire       [5:0]    _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length;
  wire       [0:0]    _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_valid;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_ready;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_opcode;
  wire       [31:0]   system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_address;
  wire       [5:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_length;
  wire       [63:0]   system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_data;
  wire       [7:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_mask;
  wire       [4:0]    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_context;
  reg                 _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1;
  reg                 _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all_1;
  reg        [31:0]   _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address_1;
  reg        [5:0]    _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length_1;
  reg        [0:0]    _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source_1;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_m2sPipe_valid;
  wire                system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_m2sPipe_ready;
  reg                 system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_rValid;
  wire                when_Stream_l375_16;
  wire                system_fabric_invalidationMonitor_output_connector_decoder_cmd_valid;
  wire                system_fabric_invalidationMonitor_output_connector_decoder_cmd_ready;
  wire                system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_mask;
  wire       [43:0]   system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_context;
  wire                system_fabric_invalidationMonitor_output_connector_decoder_rsp_valid;
  wire                system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready;
  wire                system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_last;
  wire       [0:0]    system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_data;
  wire       [43:0]   system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_context;
  reg                 _zz_system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready;
  wire                io_output_cmd_s2mPipe_valid;
  reg                 io_output_cmd_s2mPipe_ready;
  wire                io_output_cmd_s2mPipe_payload_last;
  wire       [0:0]    io_output_cmd_s2mPipe_payload_fragment_source;
  wire       [0:0]    io_output_cmd_s2mPipe_payload_fragment_opcode;
  wire       [31:0]   io_output_cmd_s2mPipe_payload_fragment_address;
  wire       [5:0]    io_output_cmd_s2mPipe_payload_fragment_length;
  wire       [63:0]   io_output_cmd_s2mPipe_payload_fragment_data;
  wire       [7:0]    io_output_cmd_s2mPipe_payload_fragment_mask;
  wire       [43:0]   io_output_cmd_s2mPipe_payload_fragment_context;
  reg                 io_output_cmd_rValidN;
  reg                 io_output_cmd_rData_last;
  reg        [0:0]    io_output_cmd_rData_fragment_source;
  reg        [0:0]    io_output_cmd_rData_fragment_opcode;
  reg        [31:0]   io_output_cmd_rData_fragment_address;
  reg        [5:0]    io_output_cmd_rData_fragment_length;
  reg        [63:0]   io_output_cmd_rData_fragment_data;
  reg        [7:0]    io_output_cmd_rData_fragment_mask;
  reg        [43:0]   io_output_cmd_rData_fragment_context;
  wire                io_output_cmd_s2mPipe_m2sPipe_valid;
  wire                io_output_cmd_s2mPipe_m2sPipe_ready;
  wire                io_output_cmd_s2mPipe_m2sPipe_payload_last;
  wire       [0:0]    io_output_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  wire       [0:0]    io_output_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   io_output_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  wire       [5:0]    io_output_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  wire       [63:0]   io_output_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  wire       [7:0]    io_output_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  wire       [43:0]   io_output_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  reg                 io_output_cmd_s2mPipe_rValid;
  reg                 io_output_cmd_s2mPipe_rData_last;
  reg        [0:0]    io_output_cmd_s2mPipe_rData_fragment_source;
  reg        [0:0]    io_output_cmd_s2mPipe_rData_fragment_opcode;
  reg        [31:0]   io_output_cmd_s2mPipe_rData_fragment_address;
  reg        [5:0]    io_output_cmd_s2mPipe_rData_fragment_length;
  reg        [63:0]   io_output_cmd_s2mPipe_rData_fragment_data;
  reg        [7:0]    io_output_cmd_s2mPipe_rData_fragment_mask;
  reg        [43:0]   io_output_cmd_s2mPipe_rData_fragment_context;
  wire                when_Stream_l375_17;
  wire                _zz_when_Stream_l375;
  reg                 _zz_when_Stream_l375_1;
  reg                 _zz_io_output_rsp_payload_last;
  reg        [0:0]    _zz_io_output_rsp_payload_fragment_source;
  reg        [0:0]    _zz_io_output_rsp_payload_fragment_opcode;
  reg        [63:0]   _zz_io_output_rsp_payload_fragment_data;
  reg        [43:0]   _zz_io_output_rsp_payload_fragment_context;
  wire                when_Stream_l375_18;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [3:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_ready;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all;
  wire       [31:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_valid;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_valid;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_ready;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_payload_source;
  reg                 _zz_io_input_rsp_ready;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid;
  reg                 system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length;
  wire       [63:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data;
  wire       [7:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask;
  wire       [3:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context;
  reg                 system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN;
  reg                 system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source;
  reg        [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg                 system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_exclusive;
  reg        [31:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [5:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [63:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [7:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask;
  reg        [3:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  wire       [63:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  wire       [7:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  wire       [3:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  reg                 system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid;
  reg                 system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last;
  reg        [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source;
  reg        [0:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode;
  reg                 system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_exclusive;
  reg        [31:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address;
  reg        [5:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length;
  reg        [63:0]   system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data;
  reg        [7:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask;
  reg        [3:0]    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context;
  wire                when_Stream_l375_19;
  wire                _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  reg                 _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  reg                 _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  reg        [0:0]    _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  reg        [0:0]    _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  reg                 _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_exclusive;
  reg        [63:0]   _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  reg        [3:0]    _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                when_Stream_l375_20;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_combStage_valid;
  wire                system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_combStage_ready;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_cmd_valid;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_cmd_ready;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_mask;
  wire       [4:0]    system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_context;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_rsp_valid;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_rsp_ready;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_last;
  wire       [0:0]    system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_data;
  wire       [4:0]    system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_context;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_inv_valid;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_inv_ready;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_all;
  wire       [31:0]   system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_address;
  wire       [5:0]    system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_length;
  wire       [0:0]    system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_source;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_ack_valid;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_ack_ready;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_sync_valid;
  wire                system_fabric_exclusiveMonitor_output_connector_decoder_sync_ready;
  wire       [0:0]    system_fabric_exclusiveMonitor_output_connector_decoder_sync_payload_source;
  wire                system_fabric_dBusCoherent_bmb_cmd_valid;
  wire                system_fabric_dBusCoherent_bmb_cmd_ready;
  wire                system_fabric_dBusCoherent_bmb_cmd_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_cmd_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_cmd_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_dBusCoherent_bmb_cmd_payload_fragment_mask;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_cmd_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_rsp_valid;
  wire                system_fabric_dBusCoherent_bmb_rsp_ready;
  wire                system_fabric_dBusCoherent_bmb_rsp_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_rsp_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_rsp_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_inv_valid;
  wire                system_fabric_dBusCoherent_bmb_inv_ready;
  wire                system_fabric_dBusCoherent_bmb_inv_payload_all;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_inv_payload_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_inv_payload_length;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_inv_payload_source;
  wire                system_fabric_dBusCoherent_bmb_ack_valid;
  wire                system_fabric_dBusCoherent_bmb_ack_ready;
  wire                system_fabric_dBusCoherent_bmb_sync_valid;
  wire                system_fabric_dBusCoherent_bmb_sync_ready;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_sync_payload_source;
  wire                system_fabric_dBus_bmb_cmd_valid;
  wire                system_fabric_dBus_bmb_cmd_ready;
  wire                system_fabric_dBus_bmb_cmd_payload_last;
  wire       [0:0]    system_fabric_dBus_bmb_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_dBus_bmb_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_dBus_bmb_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_dBus_bmb_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_dBus_bmb_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_dBus_bmb_cmd_payload_fragment_mask;
  wire       [43:0]   system_fabric_dBus_bmb_cmd_payload_fragment_context;
  wire                system_fabric_dBus_bmb_rsp_valid;
  wire                system_fabric_dBus_bmb_rsp_ready;
  wire                system_fabric_dBus_bmb_rsp_payload_last;
  wire       [0:0]    system_fabric_dBus_bmb_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_dBus_bmb_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_dBus_bmb_rsp_payload_fragment_data;
  wire       [43:0]   system_fabric_dBus_bmb_rsp_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_cmd_valid;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_cmd_ready;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_exclusive;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_mask;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_rsp_valid;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_rsp_ready;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_last;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_opcode;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_exclusive;
  wire       [63:0]   system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_data;
  wire       [3:0]    system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_context;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_inv_valid;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_inv_ready;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_all;
  wire       [31:0]   system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_address;
  wire       [5:0]    system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_length;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_source;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_ack_valid;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_ack_ready;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_sync_valid;
  wire                system_fabric_dBusCoherent_bmb_connector_decoder_sync_ready;
  wire       [0:0]    system_fabric_dBusCoherent_bmb_connector_decoder_sync_payload_source;
  wire                system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  wire       [0:0]    system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [31:0]   system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [5:0]    system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [63:0]   system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [7:0]    system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [43:0]   system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [63:0]   system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [43:0]   system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_fabric_iBus_bmb_cmd_m2sPipe_valid;
  wire                system_fabric_iBus_bmb_cmd_m2sPipe_ready;
  wire                system_fabric_iBus_bmb_cmd_m2sPipe_payload_last;
  wire       [0:0]    system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_source;
  wire       [0:0]    system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_address;
  wire       [5:0]    system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_length;
  reg                 system_fabric_iBus_bmb_cmd_rValid;
  reg                 system_fabric_iBus_bmb_cmd_rData_last;
  reg        [0:0]    system_fabric_iBus_bmb_cmd_rData_fragment_source;
  reg        [0:0]    system_fabric_iBus_bmb_cmd_rData_fragment_opcode;
  reg        [31:0]   system_fabric_iBus_bmb_cmd_rData_fragment_address;
  reg        [5:0]    system_fabric_iBus_bmb_cmd_rData_fragment_length;
  wire                when_Stream_l375_21;
  wire                system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid;
  wire                system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready;
  wire                system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last;
  wire       [0:0]    system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_context;
  wire                system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid;
  wire                system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready;
  wire                system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last;
  wire       [0:0]    system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_context;
  wire                system_bridge_bmb_cmd_valid;
  wire                system_bridge_bmb_cmd_ready;
  wire                system_bridge_bmb_cmd_payload_last;
  wire       [1:0]    system_bridge_bmb_cmd_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_cmd_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_cmd_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_cmd_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_cmd_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_cmd_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_cmd_payload_fragment_context;
  wire                system_bridge_bmb_rsp_valid;
  wire                system_bridge_bmb_rsp_ready;
  wire                system_bridge_bmb_rsp_payload_last;
  wire       [1:0]    system_bridge_bmb_rsp_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_rsp_payload_fragment_opcode;
  wire       [63:0]   system_bridge_bmb_rsp_payload_fragment_data;
  wire       [43:0]   system_bridge_bmb_rsp_payload_fragment_context;
  reg                 _zz_io_input_rsp_ready_1;
  wire                io_output_cmd_m2sPipe_valid;
  wire                io_output_cmd_m2sPipe_ready;
  wire                io_output_cmd_m2sPipe_payload_last;
  wire       [1:0]    io_output_cmd_m2sPipe_payload_fragment_source;
  wire       [0:0]    io_output_cmd_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   io_output_cmd_m2sPipe_payload_fragment_address;
  wire       [5:0]    io_output_cmd_m2sPipe_payload_fragment_length;
  wire       [127:0]  io_output_cmd_m2sPipe_payload_fragment_data;
  wire       [15:0]   io_output_cmd_m2sPipe_payload_fragment_mask;
  wire       [45:0]   io_output_cmd_m2sPipe_payload_fragment_context;
  reg                 io_output_cmd_rValid;
  reg                 io_output_cmd_rData_last_1;
  reg        [1:0]    io_output_cmd_rData_fragment_source_1;
  reg        [0:0]    io_output_cmd_rData_fragment_opcode_1;
  reg        [31:0]   io_output_cmd_rData_fragment_address_1;
  reg        [5:0]    io_output_cmd_rData_fragment_length_1;
  reg        [127:0]  io_output_cmd_rData_fragment_data_1;
  reg        [15:0]   io_output_cmd_rData_fragment_mask_1;
  reg        [45:0]   io_output_cmd_rData_fragment_context_1;
  wire                when_Stream_l375_22;
  wire                _zz_when_Stream_l375_2;
  reg                 _zz_when_Stream_l375_3;
  reg                 _zz_io_output_rsp_payload_last_1;
  reg        [1:0]    _zz_io_output_rsp_payload_fragment_source_1;
  reg        [0:0]    _zz_io_output_rsp_payload_fragment_opcode_1;
  reg        [127:0]  _zz_io_output_rsp_payload_fragment_data_1;
  reg        [45:0]   _zz_io_output_rsp_payload_fragment_context_1;
  wire                when_Stream_l375_23;
  wire                system_ddr_ddrLogic_cpuAccess_arw_valid;
  wire                system_ddr_ddrLogic_cpuAccess_arw_ready;
  wire       [31:0]   system_ddr_ddrLogic_cpuAccess_arw_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_cpuAccess_arw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_cpuAccess_arw_payload_size;
  wire       [3:0]    system_ddr_ddrLogic_cpuAccess_arw_payload_cache;
  wire       [2:0]    system_ddr_ddrLogic_cpuAccess_arw_payload_prot;
  wire                system_ddr_ddrLogic_cpuAccess_arw_payload_write;
  wire                system_ddr_ddrLogic_cpuAccess_w_valid;
  wire                system_ddr_ddrLogic_cpuAccess_w_ready;
  wire       [127:0]  system_ddr_ddrLogic_cpuAccess_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_cpuAccess_w_payload_strb;
  wire                system_ddr_ddrLogic_cpuAccess_w_payload_last;
  wire                system_ddr_ddrLogic_cpuAccess_b_valid;
  wire                system_ddr_ddrLogic_cpuAccess_b_ready;
  wire       [1:0]    system_ddr_ddrLogic_cpuAccess_b_payload_resp;
  wire                system_ddr_ddrLogic_cpuAccess_r_valid;
  wire                system_ddr_ddrLogic_cpuAccess_r_ready;
  wire       [127:0]  system_ddr_ddrLogic_cpuAccess_r_payload_data;
  wire       [1:0]    system_ddr_ddrLogic_cpuAccess_r_payload_resp;
  wire                system_ddr_ddrLogic_cpuAccess_r_payload_last;
  wire                io_output_arw_s2mPipe_valid;
  reg                 io_output_arw_s2mPipe_ready;
  wire       [31:0]   io_output_arw_s2mPipe_payload_addr;
  wire       [7:0]    io_output_arw_s2mPipe_payload_len;
  wire       [2:0]    io_output_arw_s2mPipe_payload_size;
  wire       [3:0]    io_output_arw_s2mPipe_payload_cache;
  wire       [2:0]    io_output_arw_s2mPipe_payload_prot;
  wire                io_output_arw_s2mPipe_payload_write;
  reg                 io_output_arw_rValidN;
  reg        [31:0]   io_output_arw_rData_addr;
  reg        [7:0]    io_output_arw_rData_len;
  reg        [2:0]    io_output_arw_rData_size;
  reg        [3:0]    io_output_arw_rData_cache;
  reg        [2:0]    io_output_arw_rData_prot;
  reg                 io_output_arw_rData_write;
  wire                io_output_arw_s2mPipe_m2sPipe_valid;
  reg                 io_output_arw_s2mPipe_m2sPipe_ready;
  wire       [31:0]   io_output_arw_s2mPipe_m2sPipe_payload_addr;
  wire       [7:0]    io_output_arw_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    io_output_arw_s2mPipe_m2sPipe_payload_size;
  wire       [3:0]    io_output_arw_s2mPipe_m2sPipe_payload_cache;
  wire       [2:0]    io_output_arw_s2mPipe_m2sPipe_payload_prot;
  wire                io_output_arw_s2mPipe_m2sPipe_payload_write;
  reg                 io_output_arw_s2mPipe_rValid;
  reg        [31:0]   io_output_arw_s2mPipe_rData_addr;
  reg        [7:0]    io_output_arw_s2mPipe_rData_len;
  reg        [2:0]    io_output_arw_s2mPipe_rData_size;
  reg        [3:0]    io_output_arw_s2mPipe_rData_cache;
  reg        [2:0]    io_output_arw_s2mPipe_rData_prot;
  reg                 io_output_arw_s2mPipe_rData_write;
  wire                when_Stream_l375_24;
  wire                io_output_arw_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                io_output_arw_s2mPipe_m2sPipe_m2sPipe_ready;
  wire       [31:0]   io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_addr;
  wire       [7:0]    io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_len;
  wire       [2:0]    io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_size;
  wire       [3:0]    io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_cache;
  wire       [2:0]    io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_prot;
  wire                io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_write;
  reg                 io_output_arw_s2mPipe_m2sPipe_rValid;
  reg        [31:0]   io_output_arw_s2mPipe_m2sPipe_rData_addr;
  reg        [7:0]    io_output_arw_s2mPipe_m2sPipe_rData_len;
  reg        [2:0]    io_output_arw_s2mPipe_m2sPipe_rData_size;
  reg        [3:0]    io_output_arw_s2mPipe_m2sPipe_rData_cache;
  reg        [2:0]    io_output_arw_s2mPipe_m2sPipe_rData_prot;
  reg                 io_output_arw_s2mPipe_m2sPipe_rData_write;
  wire                when_Stream_l375_25;
  wire                io_output_w_s2mPipe_valid;
  reg                 io_output_w_s2mPipe_ready;
  wire       [127:0]  io_output_w_s2mPipe_payload_data;
  wire       [15:0]   io_output_w_s2mPipe_payload_strb;
  wire                io_output_w_s2mPipe_payload_last;
  reg                 io_output_w_rValidN;
  reg        [127:0]  io_output_w_rData_data;
  reg        [15:0]   io_output_w_rData_strb;
  reg                 io_output_w_rData_last;
  wire                io_output_w_s2mPipe_m2sPipe_valid;
  reg                 io_output_w_s2mPipe_m2sPipe_ready;
  wire       [127:0]  io_output_w_s2mPipe_m2sPipe_payload_data;
  wire       [15:0]   io_output_w_s2mPipe_m2sPipe_payload_strb;
  wire                io_output_w_s2mPipe_m2sPipe_payload_last;
  reg                 io_output_w_s2mPipe_rValid;
  reg        [127:0]  io_output_w_s2mPipe_rData_data;
  reg        [15:0]   io_output_w_s2mPipe_rData_strb;
  reg                 io_output_w_s2mPipe_rData_last;
  wire                when_Stream_l375_26;
  wire                io_output_w_s2mPipe_m2sPipe_m2sPipe_valid;
  wire                io_output_w_s2mPipe_m2sPipe_m2sPipe_ready;
  wire       [127:0]  io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_data;
  wire       [15:0]   io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_strb;
  wire                io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_last;
  reg                 io_output_w_s2mPipe_m2sPipe_rValid;
  reg        [127:0]  io_output_w_s2mPipe_m2sPipe_rData_data;
  reg        [15:0]   io_output_w_s2mPipe_m2sPipe_rData_strb;
  reg                 io_output_w_s2mPipe_m2sPipe_rData_last;
  wire                when_Stream_l375_27;
  wire                system_ddr_ddrLogic_cpuAccess_b_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_cpuAccess_b_s2mPipe_ready;
  wire       [1:0]    system_ddr_ddrLogic_cpuAccess_b_s2mPipe_payload_resp;
  reg                 system_ddr_ddrLogic_cpuAccess_b_rValidN;
  reg        [1:0]    system_ddr_ddrLogic_cpuAccess_b_rData_resp;
  wire                system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_ready;
  wire       [1:0]    system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_payload_resp;
  reg                 system_ddr_ddrLogic_cpuAccess_b_s2mPipe_rValid;
  reg        [1:0]    system_ddr_ddrLogic_cpuAccess_b_s2mPipe_rData_resp;
  wire                when_Stream_l375_28;
  wire                system_ddr_ddrLogic_cpuAccess_r_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_cpuAccess_r_s2mPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_data;
  wire       [1:0]    system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_resp;
  wire                system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_last;
  reg                 system_ddr_ddrLogic_cpuAccess_r_rValidN;
  reg        [127:0]  system_ddr_ddrLogic_cpuAccess_r_rData_data;
  reg        [1:0]    system_ddr_ddrLogic_cpuAccess_r_rData_resp;
  reg                 system_ddr_ddrLogic_cpuAccess_r_rData_last;
  wire                system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_data;
  wire       [1:0]    system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_resp;
  wire                system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_last;
  reg                 system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rValid;
  reg        [127:0]  system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_data;
  reg        [1:0]    system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_resp;
  reg                 system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_last;
  wire                when_Stream_l375_29;
  wire       [3:0]    _zz_io_inputs_0_ar_payload_region;
  wire       [3:0]    _zz_io_inputs_0_aw_payload_region;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_b_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_b_ready;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_r_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_r_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_last;
  wire                io_ddrMasters_1_aw_s2mPipe_valid;
  reg                 io_ddrMasters_1_aw_s2mPipe_ready;
  wire       [31:0]   io_ddrMasters_1_aw_s2mPipe_payload_addr;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_payload_id;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_payload_region;
  wire       [7:0]    io_ddrMasters_1_aw_s2mPipe_payload_len;
  wire       [2:0]    io_ddrMasters_1_aw_s2mPipe_payload_size;
  wire       [1:0]    io_ddrMasters_1_aw_s2mPipe_payload_burst;
  wire       [0:0]    io_ddrMasters_1_aw_s2mPipe_payload_lock;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_payload_cache;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_payload_qos;
  wire       [2:0]    io_ddrMasters_1_aw_s2mPipe_payload_prot;
  reg                 io_ddrMasters_1_aw_rValidN;
  reg        [31:0]   io_ddrMasters_1_aw_rData_addr;
  reg        [3:0]    io_ddrMasters_1_aw_rData_id;
  reg        [3:0]    io_ddrMasters_1_aw_rData_region;
  reg        [7:0]    io_ddrMasters_1_aw_rData_len;
  reg        [2:0]    io_ddrMasters_1_aw_rData_size;
  reg        [1:0]    io_ddrMasters_1_aw_rData_burst;
  reg        [0:0]    io_ddrMasters_1_aw_rData_lock;
  reg        [3:0]    io_ddrMasters_1_aw_rData_cache;
  reg        [3:0]    io_ddrMasters_1_aw_rData_qos;
  reg        [2:0]    io_ddrMasters_1_aw_rData_prot;
  wire                io_ddrMasters_1_aw_s2mPipe_m2sPipe_valid;
  wire                io_ddrMasters_1_aw_s2mPipe_m2sPipe_ready;
  wire       [31:0]   io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_addr;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_id;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_region;
  wire       [7:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_burst;
  wire       [0:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_lock;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_cache;
  wire       [3:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_qos;
  wire       [2:0]    io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_prot;
  reg                 io_ddrMasters_1_aw_s2mPipe_rValid;
  reg        [31:0]   io_ddrMasters_1_aw_s2mPipe_rData_addr;
  reg        [3:0]    io_ddrMasters_1_aw_s2mPipe_rData_id;
  reg        [3:0]    io_ddrMasters_1_aw_s2mPipe_rData_region;
  reg        [7:0]    io_ddrMasters_1_aw_s2mPipe_rData_len;
  reg        [2:0]    io_ddrMasters_1_aw_s2mPipe_rData_size;
  reg        [1:0]    io_ddrMasters_1_aw_s2mPipe_rData_burst;
  reg        [0:0]    io_ddrMasters_1_aw_s2mPipe_rData_lock;
  reg        [3:0]    io_ddrMasters_1_aw_s2mPipe_rData_cache;
  reg        [3:0]    io_ddrMasters_1_aw_s2mPipe_rData_qos;
  reg        [2:0]    io_ddrMasters_1_aw_s2mPipe_rData_prot;
  wire                when_Stream_l375_30;
  wire                io_ddrMasters_1_ar_halfPipe_valid;
  wire                io_ddrMasters_1_ar_halfPipe_ready;
  wire       [31:0]   io_ddrMasters_1_ar_halfPipe_payload_addr;
  wire       [3:0]    io_ddrMasters_1_ar_halfPipe_payload_id;
  wire       [3:0]    io_ddrMasters_1_ar_halfPipe_payload_region;
  wire       [7:0]    io_ddrMasters_1_ar_halfPipe_payload_len;
  wire       [2:0]    io_ddrMasters_1_ar_halfPipe_payload_size;
  wire       [1:0]    io_ddrMasters_1_ar_halfPipe_payload_burst;
  wire       [0:0]    io_ddrMasters_1_ar_halfPipe_payload_lock;
  wire       [3:0]    io_ddrMasters_1_ar_halfPipe_payload_cache;
  wire       [3:0]    io_ddrMasters_1_ar_halfPipe_payload_qos;
  wire       [2:0]    io_ddrMasters_1_ar_halfPipe_payload_prot;
  reg                 io_ddrMasters_1_ar_rValid;
  wire                io_ddrMasters_1_ar_halfPipe_fire;
  reg        [31:0]   io_ddrMasters_1_ar_rData_addr;
  reg        [3:0]    io_ddrMasters_1_ar_rData_id;
  reg        [3:0]    io_ddrMasters_1_ar_rData_region;
  reg        [7:0]    io_ddrMasters_1_ar_rData_len;
  reg        [2:0]    io_ddrMasters_1_ar_rData_size;
  reg        [1:0]    io_ddrMasters_1_ar_rData_burst;
  reg        [0:0]    io_ddrMasters_1_ar_rData_lock;
  reg        [3:0]    io_ddrMasters_1_ar_rData_cache;
  reg        [3:0]    io_ddrMasters_1_ar_rData_qos;
  reg        [2:0]    io_ddrMasters_1_ar_rData_prot;
  wire                io_ddrMasters_1_w_s2mPipe_valid;
  reg                 io_ddrMasters_1_w_s2mPipe_ready;
  wire       [31:0]   io_ddrMasters_1_w_s2mPipe_payload_data;
  wire       [3:0]    io_ddrMasters_1_w_s2mPipe_payload_strb;
  wire                io_ddrMasters_1_w_s2mPipe_payload_last;
  reg                 io_ddrMasters_1_w_rValidN;
  reg        [31:0]   io_ddrMasters_1_w_rData_data;
  reg        [3:0]    io_ddrMasters_1_w_rData_strb;
  reg                 io_ddrMasters_1_w_rData_last;
  wire                io_ddrMasters_1_w_s2mPipe_m2sPipe_valid;
  wire                io_ddrMasters_1_w_s2mPipe_m2sPipe_ready;
  wire       [31:0]   io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_data;
  wire       [3:0]    io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_strb;
  wire                io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_last;
  reg                 io_ddrMasters_1_w_s2mPipe_rValid;
  reg        [31:0]   io_ddrMasters_1_w_s2mPipe_rData_data;
  reg        [3:0]    io_ddrMasters_1_w_s2mPipe_rData_strb;
  reg                 io_ddrMasters_1_w_s2mPipe_rData_last;
  wire                when_Stream_l375_31;
  wire                io_input_r_m2sPipe_valid;
  wire                io_input_r_m2sPipe_ready;
  wire       [31:0]   io_input_r_m2sPipe_payload_data;
  wire       [3:0]    io_input_r_m2sPipe_payload_id;
  wire       [1:0]    io_input_r_m2sPipe_payload_resp;
  wire                io_input_r_m2sPipe_payload_last;
  reg                 io_input_r_rValid;
  reg        [31:0]   io_input_r_rData_data;
  reg        [3:0]    io_input_r_rData_id;
  reg        [1:0]    io_input_r_rData_resp;
  reg                 io_input_r_rData_last;
  wire                when_Stream_l375_32;
  wire                io_input_b_s2mPipe_valid;
  reg                 io_input_b_s2mPipe_ready;
  wire       [3:0]    io_input_b_s2mPipe_payload_id;
  wire       [1:0]    io_input_b_s2mPipe_payload_resp;
  reg                 io_input_b_rValidN;
  reg        [3:0]    io_input_b_rData_id;
  reg        [1:0]    io_input_b_rData_resp;
  wire                io_input_b_s2mPipe_m2sPipe_valid;
  wire                io_input_b_s2mPipe_m2sPipe_ready;
  wire       [3:0]    io_input_b_s2mPipe_m2sPipe_payload_id;
  wire       [1:0]    io_input_b_s2mPipe_m2sPipe_payload_resp;
  reg                 io_input_b_s2mPipe_rValid;
  reg        [3:0]    io_input_b_s2mPipe_rData_id;
  reg        [1:0]    io_input_b_s2mPipe_rData_resp;
  wire                when_Stream_l375_33;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_ready;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_prot;
  reg                 system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rValid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_fire;
  reg        [31:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_addr;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_prot;
  reg                 system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rValid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_fire;
  reg        [31:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_addr;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_prot;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_data;
  reg        [15:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_strb;
  reg                 system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_last;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rValid;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_data;
  reg        [15:0]   system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_strb;
  reg                 system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_last;
  wire                when_Stream_l375_34;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_data;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_resp;
  reg                 system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_last;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rValid;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_data;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_resp;
  reg                 system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_last;
  wire                when_Stream_l375_35;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_ready;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_payload_resp;
  reg                 system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rValid;
  wire                system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_fire;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rData_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_b_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_b_ready;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_r_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_r_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_last;
  wire                io_ddrMasters_0_aw_s2mPipe_valid;
  reg                 io_ddrMasters_0_aw_s2mPipe_ready;
  wire       [31:0]   io_ddrMasters_0_aw_s2mPipe_payload_addr;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_payload_id;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_payload_region;
  wire       [7:0]    io_ddrMasters_0_aw_s2mPipe_payload_len;
  wire       [2:0]    io_ddrMasters_0_aw_s2mPipe_payload_size;
  wire       [1:0]    io_ddrMasters_0_aw_s2mPipe_payload_burst;
  wire       [0:0]    io_ddrMasters_0_aw_s2mPipe_payload_lock;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_payload_cache;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_payload_qos;
  wire       [2:0]    io_ddrMasters_0_aw_s2mPipe_payload_prot;
  reg                 io_ddrMasters_0_aw_rValidN;
  reg        [31:0]   io_ddrMasters_0_aw_rData_addr;
  reg        [3:0]    io_ddrMasters_0_aw_rData_id;
  reg        [3:0]    io_ddrMasters_0_aw_rData_region;
  reg        [7:0]    io_ddrMasters_0_aw_rData_len;
  reg        [2:0]    io_ddrMasters_0_aw_rData_size;
  reg        [1:0]    io_ddrMasters_0_aw_rData_burst;
  reg        [0:0]    io_ddrMasters_0_aw_rData_lock;
  reg        [3:0]    io_ddrMasters_0_aw_rData_cache;
  reg        [3:0]    io_ddrMasters_0_aw_rData_qos;
  reg        [2:0]    io_ddrMasters_0_aw_rData_prot;
  wire                io_ddrMasters_0_aw_s2mPipe_m2sPipe_valid;
  wire                io_ddrMasters_0_aw_s2mPipe_m2sPipe_ready;
  wire       [31:0]   io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_addr;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_id;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_region;
  wire       [7:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_burst;
  wire       [0:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_lock;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_cache;
  wire       [3:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_qos;
  wire       [2:0]    io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_prot;
  reg                 io_ddrMasters_0_aw_s2mPipe_rValid;
  reg        [31:0]   io_ddrMasters_0_aw_s2mPipe_rData_addr;
  reg        [3:0]    io_ddrMasters_0_aw_s2mPipe_rData_id;
  reg        [3:0]    io_ddrMasters_0_aw_s2mPipe_rData_region;
  reg        [7:0]    io_ddrMasters_0_aw_s2mPipe_rData_len;
  reg        [2:0]    io_ddrMasters_0_aw_s2mPipe_rData_size;
  reg        [1:0]    io_ddrMasters_0_aw_s2mPipe_rData_burst;
  reg        [0:0]    io_ddrMasters_0_aw_s2mPipe_rData_lock;
  reg        [3:0]    io_ddrMasters_0_aw_s2mPipe_rData_cache;
  reg        [3:0]    io_ddrMasters_0_aw_s2mPipe_rData_qos;
  reg        [2:0]    io_ddrMasters_0_aw_s2mPipe_rData_prot;
  wire                when_Stream_l375_36;
  wire                io_ddrMasters_0_ar_halfPipe_valid;
  wire                io_ddrMasters_0_ar_halfPipe_ready;
  wire       [31:0]   io_ddrMasters_0_ar_halfPipe_payload_addr;
  wire       [3:0]    io_ddrMasters_0_ar_halfPipe_payload_id;
  wire       [3:0]    io_ddrMasters_0_ar_halfPipe_payload_region;
  wire       [7:0]    io_ddrMasters_0_ar_halfPipe_payload_len;
  wire       [2:0]    io_ddrMasters_0_ar_halfPipe_payload_size;
  wire       [1:0]    io_ddrMasters_0_ar_halfPipe_payload_burst;
  wire       [0:0]    io_ddrMasters_0_ar_halfPipe_payload_lock;
  wire       [3:0]    io_ddrMasters_0_ar_halfPipe_payload_cache;
  wire       [3:0]    io_ddrMasters_0_ar_halfPipe_payload_qos;
  wire       [2:0]    io_ddrMasters_0_ar_halfPipe_payload_prot;
  reg                 io_ddrMasters_0_ar_rValid;
  wire                io_ddrMasters_0_ar_halfPipe_fire;
  reg        [31:0]   io_ddrMasters_0_ar_rData_addr;
  reg        [3:0]    io_ddrMasters_0_ar_rData_id;
  reg        [3:0]    io_ddrMasters_0_ar_rData_region;
  reg        [7:0]    io_ddrMasters_0_ar_rData_len;
  reg        [2:0]    io_ddrMasters_0_ar_rData_size;
  reg        [1:0]    io_ddrMasters_0_ar_rData_burst;
  reg        [0:0]    io_ddrMasters_0_ar_rData_lock;
  reg        [3:0]    io_ddrMasters_0_ar_rData_cache;
  reg        [3:0]    io_ddrMasters_0_ar_rData_qos;
  reg        [2:0]    io_ddrMasters_0_ar_rData_prot;
  wire                io_ddrMasters_0_w_s2mPipe_valid;
  reg                 io_ddrMasters_0_w_s2mPipe_ready;
  wire       [63:0]   io_ddrMasters_0_w_s2mPipe_payload_data;
  wire       [7:0]    io_ddrMasters_0_w_s2mPipe_payload_strb;
  wire                io_ddrMasters_0_w_s2mPipe_payload_last;
  reg                 io_ddrMasters_0_w_rValidN;
  reg        [63:0]   io_ddrMasters_0_w_rData_data;
  reg        [7:0]    io_ddrMasters_0_w_rData_strb;
  reg                 io_ddrMasters_0_w_rData_last;
  wire                io_ddrMasters_0_w_s2mPipe_m2sPipe_valid;
  wire                io_ddrMasters_0_w_s2mPipe_m2sPipe_ready;
  wire       [63:0]   io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_data;
  wire       [7:0]    io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_strb;
  wire                io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_last;
  reg                 io_ddrMasters_0_w_s2mPipe_rValid;
  reg        [63:0]   io_ddrMasters_0_w_s2mPipe_rData_data;
  reg        [7:0]    io_ddrMasters_0_w_s2mPipe_rData_strb;
  reg                 io_ddrMasters_0_w_s2mPipe_rData_last;
  wire                when_Stream_l375_37;
  wire                io_input_r_m2sPipe_valid_1;
  wire                io_input_r_m2sPipe_ready_1;
  wire       [63:0]   io_input_r_m2sPipe_payload_data_1;
  wire       [3:0]    io_input_r_m2sPipe_payload_id_1;
  wire       [1:0]    io_input_r_m2sPipe_payload_resp_1;
  wire                io_input_r_m2sPipe_payload_last_1;
  reg                 io_input_r_rValid_1;
  reg        [63:0]   io_input_r_rData_data_1;
  reg        [3:0]    io_input_r_rData_id_1;
  reg        [1:0]    io_input_r_rData_resp_1;
  reg                 io_input_r_rData_last_1;
  wire                when_Stream_l375_38;
  wire                io_input_b_s2mPipe_valid_1;
  reg                 io_input_b_s2mPipe_ready_1;
  wire       [3:0]    io_input_b_s2mPipe_payload_id_1;
  wire       [1:0]    io_input_b_s2mPipe_payload_resp_1;
  reg                 io_input_b_rValidN_1;
  reg        [3:0]    io_input_b_rData_id_1;
  reg        [1:0]    io_input_b_rData_resp_1;
  wire                io_input_b_s2mPipe_m2sPipe_valid_1;
  wire                io_input_b_s2mPipe_m2sPipe_ready_1;
  wire       [3:0]    io_input_b_s2mPipe_m2sPipe_payload_id_1;
  wire       [1:0]    io_input_b_s2mPipe_m2sPipe_payload_resp_1;
  reg                 io_input_b_s2mPipe_rValid_1;
  reg        [3:0]    io_input_b_s2mPipe_rData_id_1;
  reg        [1:0]    io_input_b_s2mPipe_rData_resp_1;
  wire                when_Stream_l375_39;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_ready;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_last;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_prot;
  reg                 system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rValid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_fire;
  reg        [31:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_addr;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_addr;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_prot;
  reg                 system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rValid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_fire;
  reg        [31:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_addr;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_prot;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_data;
  reg        [15:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_strb;
  reg                 system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_last;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_strb;
  wire                system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rValid;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_data;
  reg        [15:0]   system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_strb;
  reg                 system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_last;
  wire                when_Stream_l375_40;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_data;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_resp;
  reg                 system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_last;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_ready;
  wire       [127:0]  system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_data;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_resp;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_last;
  reg                 system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rValid;
  reg        [127:0]  system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_data;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_resp;
  reg                 system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_last;
  wire                when_Stream_l375_41;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_valid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_ready;
  wire       [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_payload_resp;
  reg                 system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rValid;
  wire                system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_fire;
  reg        [3:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rData_resp;
  wire                system_ddr_ddrLogic_ddrAAxi4_aw_valid;
  wire                system_ddr_ddrLogic_ddrAAxi4_aw_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAAxi4_aw_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_aw_payload_prot;
  reg                 system_ddr_ddrLogic_ddrAAxi4_w_valid;
  wire                system_ddr_ddrLogic_ddrAAxi4_w_ready;
  wire       [127:0]  system_ddr_ddrLogic_ddrAAxi4_w_payload_data;
  wire       [15:0]   system_ddr_ddrLogic_ddrAAxi4_w_payload_strb;
  reg                 system_ddr_ddrLogic_ddrAAxi4_w_payload_last;
  wire                system_ddr_ddrLogic_ddrAAxi4_b_valid;
  wire                system_ddr_ddrLogic_ddrAAxi4_b_ready;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_b_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_b_payload_resp;
  wire                system_ddr_ddrLogic_ddrAAxi4_ar_valid;
  wire                system_ddr_ddrLogic_ddrAAxi4_ar_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAAxi4_ar_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_payload_prot;
  wire                system_ddr_ddrLogic_ddrAAxi4_r_valid;
  wire                system_ddr_ddrLogic_ddrAAxi4_r_ready;
  wire       [127:0]  system_ddr_ddrLogic_ddrAAxi4_r_payload_data;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_r_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_r_payload_resp;
  wire                system_ddr_ddrLogic_ddrAAxi4_r_payload_last;
  wire                io_output_aw_s2mPipe_valid;
  reg                 io_output_aw_s2mPipe_ready;
  wire       [31:0]   io_output_aw_s2mPipe_payload_addr;
  wire       [7:0]    io_output_aw_s2mPipe_payload_id;
  wire       [3:0]    io_output_aw_s2mPipe_payload_region;
  wire       [7:0]    io_output_aw_s2mPipe_payload_len;
  wire       [2:0]    io_output_aw_s2mPipe_payload_size;
  wire       [1:0]    io_output_aw_s2mPipe_payload_burst;
  wire       [0:0]    io_output_aw_s2mPipe_payload_lock;
  wire       [3:0]    io_output_aw_s2mPipe_payload_cache;
  wire       [3:0]    io_output_aw_s2mPipe_payload_qos;
  wire       [2:0]    io_output_aw_s2mPipe_payload_prot;
  reg                 io_output_aw_rValidN;
  reg        [31:0]   io_output_aw_rData_addr;
  reg        [7:0]    io_output_aw_rData_id;
  reg        [3:0]    io_output_aw_rData_region;
  reg        [7:0]    io_output_aw_rData_len;
  reg        [2:0]    io_output_aw_rData_size;
  reg        [1:0]    io_output_aw_rData_burst;
  reg        [0:0]    io_output_aw_rData_lock;
  reg        [3:0]    io_output_aw_rData_cache;
  reg        [3:0]    io_output_aw_rData_qos;
  reg        [2:0]    io_output_aw_rData_prot;
  wire                io_output_aw_s2mPipe_m2sPipe_valid;
  wire                io_output_aw_s2mPipe_m2sPipe_ready;
  wire       [31:0]   io_output_aw_s2mPipe_m2sPipe_payload_addr;
  wire       [7:0]    io_output_aw_s2mPipe_m2sPipe_payload_id;
  wire       [3:0]    io_output_aw_s2mPipe_m2sPipe_payload_region;
  wire       [7:0]    io_output_aw_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    io_output_aw_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    io_output_aw_s2mPipe_m2sPipe_payload_burst;
  wire       [0:0]    io_output_aw_s2mPipe_m2sPipe_payload_lock;
  wire       [3:0]    io_output_aw_s2mPipe_m2sPipe_payload_cache;
  wire       [3:0]    io_output_aw_s2mPipe_m2sPipe_payload_qos;
  wire       [2:0]    io_output_aw_s2mPipe_m2sPipe_payload_prot;
  reg                 io_output_aw_s2mPipe_rValid;
  reg        [31:0]   io_output_aw_s2mPipe_rData_addr;
  reg        [7:0]    io_output_aw_s2mPipe_rData_id;
  reg        [3:0]    io_output_aw_s2mPipe_rData_region;
  reg        [7:0]    io_output_aw_s2mPipe_rData_len;
  reg        [2:0]    io_output_aw_s2mPipe_rData_size;
  reg        [1:0]    io_output_aw_s2mPipe_rData_burst;
  reg        [0:0]    io_output_aw_s2mPipe_rData_lock;
  reg        [3:0]    io_output_aw_s2mPipe_rData_cache;
  reg        [3:0]    io_output_aw_s2mPipe_rData_qos;
  reg        [2:0]    io_output_aw_s2mPipe_rData_prot;
  wire                when_Stream_l375_42;
  wire                io_output_ar_s2mPipe_valid;
  reg                 io_output_ar_s2mPipe_ready;
  wire       [31:0]   io_output_ar_s2mPipe_payload_addr;
  wire       [7:0]    io_output_ar_s2mPipe_payload_id;
  wire       [3:0]    io_output_ar_s2mPipe_payload_region;
  wire       [7:0]    io_output_ar_s2mPipe_payload_len;
  wire       [2:0]    io_output_ar_s2mPipe_payload_size;
  wire       [1:0]    io_output_ar_s2mPipe_payload_burst;
  wire       [0:0]    io_output_ar_s2mPipe_payload_lock;
  wire       [3:0]    io_output_ar_s2mPipe_payload_cache;
  wire       [3:0]    io_output_ar_s2mPipe_payload_qos;
  wire       [2:0]    io_output_ar_s2mPipe_payload_prot;
  reg                 io_output_ar_rValidN;
  reg        [31:0]   io_output_ar_rData_addr;
  reg        [7:0]    io_output_ar_rData_id;
  reg        [3:0]    io_output_ar_rData_region;
  reg        [7:0]    io_output_ar_rData_len;
  reg        [2:0]    io_output_ar_rData_size;
  reg        [1:0]    io_output_ar_rData_burst;
  reg        [0:0]    io_output_ar_rData_lock;
  reg        [3:0]    io_output_ar_rData_cache;
  reg        [3:0]    io_output_ar_rData_qos;
  reg        [2:0]    io_output_ar_rData_prot;
  wire                io_output_ar_s2mPipe_m2sPipe_valid;
  wire                io_output_ar_s2mPipe_m2sPipe_ready;
  wire       [31:0]   io_output_ar_s2mPipe_m2sPipe_payload_addr;
  wire       [7:0]    io_output_ar_s2mPipe_m2sPipe_payload_id;
  wire       [3:0]    io_output_ar_s2mPipe_m2sPipe_payload_region;
  wire       [7:0]    io_output_ar_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    io_output_ar_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    io_output_ar_s2mPipe_m2sPipe_payload_burst;
  wire       [0:0]    io_output_ar_s2mPipe_m2sPipe_payload_lock;
  wire       [3:0]    io_output_ar_s2mPipe_m2sPipe_payload_cache;
  wire       [3:0]    io_output_ar_s2mPipe_m2sPipe_payload_qos;
  wire       [2:0]    io_output_ar_s2mPipe_m2sPipe_payload_prot;
  reg                 io_output_ar_s2mPipe_rValid;
  reg        [31:0]   io_output_ar_s2mPipe_rData_addr;
  reg        [7:0]    io_output_ar_s2mPipe_rData_id;
  reg        [3:0]    io_output_ar_s2mPipe_rData_region;
  reg        [7:0]    io_output_ar_s2mPipe_rData_len;
  reg        [2:0]    io_output_ar_s2mPipe_rData_size;
  reg        [1:0]    io_output_ar_s2mPipe_rData_burst;
  reg        [0:0]    io_output_ar_s2mPipe_rData_lock;
  reg        [3:0]    io_output_ar_s2mPipe_rData_cache;
  reg        [3:0]    io_output_ar_s2mPipe_rData_qos;
  reg        [2:0]    io_output_ar_s2mPipe_rData_prot;
  wire                when_Stream_l375_43;
  wire                io_output_w_m2sPipe_valid;
  wire                io_output_w_m2sPipe_ready;
  wire       [127:0]  io_output_w_m2sPipe_payload_data;
  wire       [15:0]   io_output_w_m2sPipe_payload_strb;
  wire                io_output_w_m2sPipe_payload_last;
  reg                 io_output_w_rValid;
  reg        [127:0]  io_output_w_rData_data_1;
  reg        [15:0]   io_output_w_rData_strb_1;
  reg                 io_output_w_rData_last_1;
  wire                when_Stream_l375_44;
  wire                system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_ready;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_payload_resp;
  reg                 system_ddr_ddrLogic_ddrAAxi4_b_rValidN;
  reg        [7:0]    system_ddr_ddrLogic_ddrAAxi4_b_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_ddrAAxi4_b_rData_resp;
  wire                system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_ready;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_payload_id;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_payload_resp;
  reg                 system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rValid;
  reg        [7:0]    system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rData_id;
  reg        [1:0]    system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rData_resp;
  wire                when_Stream_l375_45;
  reg        [4:0]    system_ddr_ddrLogic_ddrAReset_counter;
  reg                 system_ddr_ddrLogic_ddrAReset_resetUnbuffered;
  wire       [4:0]    _zz_when_TrionDdrGenerator_l257;
  wire                when_TrionDdrGenerator_l257;
  reg                 system_ddr_ddrLogic_ddrAReset_reset;
  wire                system_ddr_ddrLogic_ddrAToAxi4_ioAw_valid;
  wire                system_ddr_ddrLogic_ddrAToAxi4_ioAw_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_prot;
  wire                system_ddr_ddrLogic_ddrAToAxi4_patchAw_valid;
  wire                system_ddr_ddrLogic_ddrAToAxi4_patchAw_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_prot;
  wire                system_ddr_ddrLogic_ddrAAxi4_aw_fire;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_a2wPayload_len;
  wire                system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_valid;
  wire                system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_ready;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_payload_len;
  wire                io_pop_s2mPipe_valid_2;
  reg                 io_pop_s2mPipe_ready_2;
  wire       [7:0]    io_pop_s2mPipe_payload_len;
  reg                 io_pop_rValidN_2;
  reg        [7:0]    io_pop_rData_len;
  wire                system_ddr_ddrLogic_ddrAToAxi4_widStream_valid;
  wire                system_ddr_ddrLogic_ddrAToAxi4_widStream_ready;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_widStream_payload_len;
  reg                 io_pop_s2mPipe_rValid_2;
  reg        [7:0]    io_pop_s2mPipe_rData_len;
  wire                when_Stream_l375_46;
  wire                system_ddr_ddrLogic_ddrAAxi4_w_fire;
  reg        [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ddrA_wCounter;
  reg                 ddrCd_logic_outputReset_regNext;
  wire                when_TrionDdrGenerator_l363;
  wire                system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_prot;
  reg                 system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN;
  reg        [31:0]   system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_addr;
  reg        [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_prot;
  wire                system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_prot;
  reg                 system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rValid;
  reg        [31:0]   system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_addr;
  reg        [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_prot;
  wire                when_Stream_l375_47;
  wire                system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_valid;
  reg                 system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_prot;
  reg                 system_ddr_ddrLogic_ddrAAxi4_ar_rValidN;
  reg        [31:0]   system_ddr_ddrLogic_ddrAAxi4_ar_rData_addr;
  reg        [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_rData_prot;
  wire                system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_valid;
  wire                system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_ready;
  wire       [31:0]   system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_addr;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_id;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_region;
  wire       [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_len;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_size;
  wire       [1:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_burst;
  wire       [0:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_lock;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_cache;
  wire       [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_qos;
  wire       [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_prot;
  reg                 system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rValid;
  reg        [31:0]   system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_addr;
  reg        [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_id;
  reg        [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_region;
  reg        [7:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_len;
  reg        [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_size;
  reg        [1:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_burst;
  reg        [0:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_lock;
  reg        [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_cache;
  reg        [3:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_qos;
  reg        [2:0]    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_prot;
  wire                when_Stream_l375_48;
  wire                _zz_io_ddrA_w_valid;
  wire                io_ddrA_r_m2sPipe_valid;
  wire                io_ddrA_r_m2sPipe_ready;
  wire       [127:0]  io_ddrA_r_m2sPipe_payload_data;
  wire       [7:0]    io_ddrA_r_m2sPipe_payload_id;
  wire       [1:0]    io_ddrA_r_m2sPipe_payload_resp;
  wire                io_ddrA_r_m2sPipe_payload_last;
  reg                 io_ddrA_r_rValid;
  reg        [127:0]  io_ddrA_r_rData_data;
  reg        [7:0]    io_ddrA_r_rData_id;
  reg        [1:0]    io_ddrA_r_rData_resp;
  reg                 io_ddrA_r_rData_last;
  wire                when_Stream_l375_49;
  wire                io_ddrA_b_s2mPipe_valid;
  reg                 io_ddrA_b_s2mPipe_ready;
  wire       [7:0]    io_ddrA_b_s2mPipe_payload_id;
  wire       [1:0]    io_ddrA_b_s2mPipe_payload_resp;
  reg                 io_ddrA_b_rValidN;
  reg        [7:0]    io_ddrA_b_rData_id;
  reg        [1:0]    io_ddrA_b_rData_resp;
  wire                io_ddrA_b_s2mPipe_m2sPipe_valid;
  wire                io_ddrA_b_s2mPipe_m2sPipe_ready;
  wire       [7:0]    io_ddrA_b_s2mPipe_m2sPipe_payload_id;
  wire       [1:0]    io_ddrA_b_s2mPipe_m2sPipe_payload_resp;
  reg                 io_ddrA_b_s2mPipe_rValid;
  reg        [7:0]    io_ddrA_b_s2mPipe_rData_id;
  reg        [1:0]    io_ddrA_b_s2mPipe_rData_resp;
  wire                when_Stream_l375_50;
  reg                 ddrCd_logic_outputReset_regNext_1;
  wire                system_axiA_logic_axiAAdapted_aw_valid;
  wire                system_axiA_logic_axiAAdapted_aw_ready;
  wire       [31:0]   system_axiA_logic_axiAAdapted_aw_payload_addr;
  wire       [7:0]    system_axiA_logic_axiAAdapted_aw_payload_id;
  wire       [3:0]    system_axiA_logic_axiAAdapted_aw_payload_region;
  wire       [7:0]    system_axiA_logic_axiAAdapted_aw_payload_len;
  wire       [2:0]    system_axiA_logic_axiAAdapted_aw_payload_size;
  wire       [1:0]    system_axiA_logic_axiAAdapted_aw_payload_burst;
  wire       [0:0]    system_axiA_logic_axiAAdapted_aw_payload_lock;
  wire       [3:0]    system_axiA_logic_axiAAdapted_aw_payload_cache;
  wire       [3:0]    system_axiA_logic_axiAAdapted_aw_payload_qos;
  wire       [2:0]    system_axiA_logic_axiAAdapted_aw_payload_prot;
  wire                system_axiA_logic_axiAAdapted_w_valid;
  wire                system_axiA_logic_axiAAdapted_w_ready;
  wire       [31:0]   system_axiA_logic_axiAAdapted_w_payload_data;
  wire       [3:0]    system_axiA_logic_axiAAdapted_w_payload_strb;
  wire                system_axiA_logic_axiAAdapted_w_payload_last;
  wire                system_axiA_logic_axiAAdapted_b_valid;
  wire                system_axiA_logic_axiAAdapted_b_ready;
  wire       [7:0]    system_axiA_logic_axiAAdapted_b_payload_id;
  wire       [1:0]    system_axiA_logic_axiAAdapted_b_payload_resp;
  wire                system_axiA_logic_axiAAdapted_ar_valid;
  wire                system_axiA_logic_axiAAdapted_ar_ready;
  wire       [31:0]   system_axiA_logic_axiAAdapted_ar_payload_addr;
  wire       [7:0]    system_axiA_logic_axiAAdapted_ar_payload_id;
  wire       [3:0]    system_axiA_logic_axiAAdapted_ar_payload_region;
  wire       [7:0]    system_axiA_logic_axiAAdapted_ar_payload_len;
  wire       [2:0]    system_axiA_logic_axiAAdapted_ar_payload_size;
  wire       [1:0]    system_axiA_logic_axiAAdapted_ar_payload_burst;
  wire       [0:0]    system_axiA_logic_axiAAdapted_ar_payload_lock;
  wire       [3:0]    system_axiA_logic_axiAAdapted_ar_payload_cache;
  wire       [3:0]    system_axiA_logic_axiAAdapted_ar_payload_qos;
  wire       [2:0]    system_axiA_logic_axiAAdapted_ar_payload_prot;
  wire                system_axiA_logic_axiAAdapted_r_valid;
  wire                system_axiA_logic_axiAAdapted_r_ready;
  wire       [31:0]   system_axiA_logic_axiAAdapted_r_payload_data;
  wire       [7:0]    system_axiA_logic_axiAAdapted_r_payload_id;
  wire       [1:0]    system_axiA_logic_axiAAdapted_r_payload_resp;
  wire                system_axiA_logic_axiAAdapted_r_payload_last;
  wire       [3:0]    _zz_system_axiA_logic_axiAAdapted_ar_payload_region;
  wire       [3:0]    _zz_system_axiA_logic_axiAAdapted_aw_payload_region;
  wire                axiA_r_m2sPipe_valid;
  wire                axiA_r_m2sPipe_ready;
  wire       [31:0]   axiA_r_m2sPipe_payload_data;
  wire       [7:0]    axiA_r_m2sPipe_payload_id;
  wire       [1:0]    axiA_r_m2sPipe_payload_resp;
  wire                axiA_r_m2sPipe_payload_last;
  reg                 axiA_r_rValid;
  reg        [31:0]   axiA_r_rData_data;
  reg        [7:0]    axiA_r_rData_id;
  reg        [1:0]    axiA_r_rData_resp;
  reg                 axiA_r_rData_last;
  wire                when_Stream_l375_51;
  wire                system_bridge_bmb_cmd_s2mPipe_valid;
  reg                 system_bridge_bmb_cmd_s2mPipe_ready;
  wire                system_bridge_bmb_cmd_s2mPipe_payload_last;
  wire       [1:0]    system_bridge_bmb_cmd_s2mPipe_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_cmd_s2mPipe_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_cmd_s2mPipe_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_cmd_s2mPipe_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_cmd_s2mPipe_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_cmd_s2mPipe_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_cmd_s2mPipe_payload_fragment_context;
  reg                 system_bridge_bmb_cmd_rValidN;
  reg                 system_bridge_bmb_cmd_rData_last;
  reg        [1:0]    system_bridge_bmb_cmd_rData_fragment_source;
  reg        [0:0]    system_bridge_bmb_cmd_rData_fragment_opcode;
  reg        [31:0]   system_bridge_bmb_cmd_rData_fragment_address;
  reg        [5:0]    system_bridge_bmb_cmd_rData_fragment_length;
  reg        [63:0]   system_bridge_bmb_cmd_rData_fragment_data;
  reg        [7:0]    system_bridge_bmb_cmd_rData_fragment_mask;
  reg        [43:0]   system_bridge_bmb_cmd_rData_fragment_context;
  wire                system_bridge_bmb_cmd_s2mPipe_m2sPipe_valid;
  wire                system_bridge_bmb_cmd_s2mPipe_m2sPipe_ready;
  wire                system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_last;
  wire       [1:0]    system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  wire       [0:0]    system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  wire       [5:0]    system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  wire       [63:0]   system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  wire       [7:0]    system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  wire       [43:0]   system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  reg                 system_bridge_bmb_cmd_s2mPipe_rValid;
  reg                 system_bridge_bmb_cmd_s2mPipe_rData_last;
  reg        [1:0]    system_bridge_bmb_cmd_s2mPipe_rData_fragment_source;
  reg        [0:0]    system_bridge_bmb_cmd_s2mPipe_rData_fragment_opcode;
  reg        [31:0]   system_bridge_bmb_cmd_s2mPipe_rData_fragment_address;
  reg        [5:0]    system_bridge_bmb_cmd_s2mPipe_rData_fragment_length;
  reg        [63:0]   system_bridge_bmb_cmd_s2mPipe_rData_fragment_data;
  reg        [7:0]    system_bridge_bmb_cmd_s2mPipe_rData_fragment_mask;
  reg        [43:0]   system_bridge_bmb_cmd_s2mPipe_rData_fragment_context;
  wire                when_Stream_l375_52;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [1:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  wire       [0:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [31:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [5:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [127:0]  system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [15:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [45:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [1:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [127:0]  system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [45:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  reg                 _zz_io_input_rsp_ready_2;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid;
  reg                 system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last;
  wire       [1:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source;
  wire       [0:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode;
  wire       [31:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address;
  wire       [5:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length;
  wire       [127:0]  system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data;
  wire       [15:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask;
  wire       [45:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context;
  reg                 system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN;
  reg                 system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [1:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source;
  reg        [0:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [31:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [5:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [127:0]  system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [15:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask;
  reg        [45:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready;
  wire                system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last;
  wire       [1:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  wire       [0:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  wire       [5:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  wire       [127:0]  system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  wire       [15:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  wire       [45:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  reg                 system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid;
  reg                 system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last;
  reg        [1:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source;
  reg        [0:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode;
  reg        [31:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address;
  reg        [5:0]    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length;
  reg        [127:0]  system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data;
  reg        [15:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask;
  reg        [45:0]   system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context;
  wire                when_Stream_l375_53;
  wire                _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  reg                 _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  reg                 _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  reg        [1:0]    _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  reg        [0:0]    _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  reg        [127:0]  _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  reg        [45:0]   _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                when_Stream_l375_54;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [1:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  wire       [0:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [5:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [3:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [44:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [1:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [44:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                _zz_io_input_rsp_ready_3;
  wire                _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [1:0]    _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  wire       [0:0]    _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [44:0]   _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid;
  reg                 system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last;
  wire       [1:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source;
  wire       [0:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode;
  wire       [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address;
  wire       [5:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length;
  wire       [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data;
  wire       [3:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask;
  wire       [44:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context;
  reg                 system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN;
  reg                 system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [1:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source;
  reg        [0:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [5:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [3:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask;
  reg        [44:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready;
  wire                system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last;
  wire       [1:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  wire       [0:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  wire       [5:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  wire       [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  wire       [3:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  wire       [44:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  reg                 system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid;
  reg                 system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last;
  reg        [1:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source;
  reg        [0:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode;
  reg        [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address;
  reg        [5:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length;
  reg        [31:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data;
  reg        [3:0]    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask;
  reg        [44:0]   system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context;
  wire                when_Stream_l375_55;
  reg                 _zz_2;
  reg                 _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1;
  reg                 _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_2;
  reg        [1:0]    _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source_1;
  reg        [0:0]    _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode_1;
  reg        [31:0]   _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data_1;
  reg        [44:0]   _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context_1;
  wire                _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  reg                 _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_2;
  reg                 _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_3;
  reg        [1:0]    _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source_2;
  reg        [0:0]    _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode_2;
  reg        [31:0]   _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data_2;
  reg        [44:0]   _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context_2;
  wire                when_Stream_l375_56;
  wire       [1:0]    system_axiA_interrupt_plic_gateway_priority;
  reg                 system_axiA_interrupt_plic_gateway_ip;
  reg                 system_axiA_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_4;
  wire                system_bmbPeripheral_bmb_cmd_valid;
  wire                system_bmbPeripheral_bmb_cmd_ready;
  wire                system_bmbPeripheral_bmb_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_rsp_valid;
  wire                system_bmbPeripheral_bmb_rsp_ready;
  wire                system_bmbPeripheral_bmb_rsp_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_rsp_payload_fragment_opcode;
  wire       [31:0]   system_bmbPeripheral_bmb_rsp_payload_fragment_data;
  wire       [48:0]   system_bmbPeripheral_bmb_rsp_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [10:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [2:0]    system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [63:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [7:0]    system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  wire       [47:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [63:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [47:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  reg                 _zz_io_bus_rsp_ready;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_valid;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_ready;
  wire                system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_last;
  wire       [0:0]    system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_opcode;
  wire       [10:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_address;
  wire       [2:0]    system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_length;
  wire       [63:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_data;
  wire       [7:0]    system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_mask;
  wire       [47:0]   system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_context;
  wire                _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  reg                 _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  reg                 _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  reg        [0:0]    _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  reg        [63:0]   _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  reg        [47:0]   _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                when_Stream_l375_57;
  wire                _zz_io_input_rsp_ready_4;
  wire                system_bmbPeripheral_bmb_cmd_combStage_valid;
  wire                system_bmbPeripheral_bmb_cmd_combStage_ready;
  wire                system_bmbPeripheral_bmb_cmd_combStage_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_data;
  wire       [3:0]    system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_mask;
  wire       [48:0]   system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_context;
  wire                _zz_system_bmbPeripheral_bmb_rsp_valid;
  reg                 _zz_system_bmbPeripheral_bmb_rsp_valid_1;
  reg                 _zz_system_bmbPeripheral_bmb_rsp_payload_last;
  reg        [0:0]    _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_data;
  reg        [48:0]   _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_context;
  wire                system_userTimer_1_interrupts_0;
  wire                system_userTimer_0_interrupts_0;
  wire                system_gpio_0_io_interrupts_0;
  wire                system_gpio_0_io_interrupts_1;
  wire                system_gpio_0_io_interrupts_2;
  wire                system_gpio_0_io_interrupts_3;
  wire                _zz_system_watchdog_logic_panics_0_plic_gateway_ip;
  wire                system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [15:0]   system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [5:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                _zz_io_bus_rsp_ready_1;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [5:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [5:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire                _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  reg                 _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  reg                 _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  reg        [0:0]    _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  reg        [48:0]   _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire       [1:0]    system_uart_0_io_interrupt_plic_gateway_priority;
  reg                 system_uart_0_io_interrupt_plic_gateway_ip;
  reg                 system_uart_0_io_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_5;
  wire       [1:0]    system_spi_0_io_interrupt_plic_gateway_priority;
  reg                 system_spi_0_io_interrupt_plic_gateway_ip;
  reg                 system_spi_0_io_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_6;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [11:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [11:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [11:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire       [1:0]    system_spi_1_io_interrupt_plic_gateway_priority;
  reg                 system_spi_1_io_interrupt_plic_gateway_ip;
  reg                 system_spi_1_io_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_7;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [11:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [11:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [11:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [7:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [7:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [7:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire       [1:0]    system_i2c_0_io_interrupt_plic_gateway_priority;
  reg                 system_i2c_0_io_interrupt_plic_gateway_ip;
  reg                 system_i2c_0_io_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_8;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [7:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [7:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [7:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire       [1:0]    system_i2c_2_io_interrupt_plic_gateway_priority;
  reg                 system_i2c_2_io_interrupt_plic_gateway_ip;
  reg                 system_i2c_2_io_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_9;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [7:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [7:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [7:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire       [1:0]    system_i2c_1_io_interrupt_plic_gateway_priority;
  reg                 system_i2c_1_io_interrupt_plic_gateway_ip;
  reg                 system_i2c_1_io_interrupt_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_10;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [7:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [7:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [7:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire       [1:0]    system_userTimer_1_interrupts_0_plic_gateway_priority;
  reg                 system_userTimer_1_interrupts_0_plic_gateway_ip;
  reg                 system_userTimer_1_interrupts_0_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_11;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [7:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last;
  wire       [0:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode;
  wire       [7:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address;
  wire       [1:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length;
  wire       [31:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data;
  wire       [48:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context;
  reg                 system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  wire                system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire;
  reg                 system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  reg        [0:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  reg        [7:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  reg        [1:0]    system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  reg        [31:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  reg        [48:0]   system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  wire       [1:0]    system_userTimer_0_interrupts_0_plic_gateway_priority;
  reg                 system_userTimer_0_interrupts_0_plic_gateway_ip;
  reg                 system_userTimer_0_interrupts_0_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_12;
  wire                system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [7:0]    system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire       [1:0]    system_gpio_0_io_interrupts_0_plic_gateway_priority;
  reg                 system_gpio_0_io_interrupts_0_plic_gateway_ip;
  reg                 system_gpio_0_io_interrupts_0_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_13;
  wire       [1:0]    system_gpio_0_io_interrupts_1_plic_gateway_priority;
  reg                 system_gpio_0_io_interrupts_1_plic_gateway_ip;
  reg                 system_gpio_0_io_interrupts_1_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_14;
  wire                system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [7:0]    system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire       [1:0]    system_watchdog_logic_panics_0_plic_gateway_priority;
  reg                 system_watchdog_logic_panics_0_plic_gateway_ip;
  reg                 system_watchdog_logic_panics_0_plic_gateway_waitCompletion;
  wire                when_PlicGateway_l21_15;
  wire                io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [15:0]   io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [15:0]   io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [15:0]   io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [15:0]   io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [15:0]   io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_1;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_1;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_1;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_1;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_1;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_1;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_1;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_1;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_1;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_1;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_1;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_1;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_1;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_1;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_2;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_2;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_2;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_2;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_2;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_2;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_2;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_2;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_2;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_2;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_2;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_2;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_2;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_2;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_3;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_3;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_3;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_3;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_3;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_3;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_3;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_3;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_3;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_3;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_3;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_3;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_3;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_3;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_4;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_4;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_4;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_4;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_4;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_4;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_4;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_4;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_4;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_4;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_4;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_4;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_4;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_4;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_5;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_5;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_5;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_5;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_5;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_5;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_5;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_5;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_5;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_5;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_5;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_5;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_5;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_5;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_6;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_6;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_6;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_6;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_6;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_6;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_6;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_6;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_6;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_6;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_6;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_6;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_6;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_6;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_7;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_7;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_7;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_7;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_7;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_7;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_7;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_7;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_7;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_7;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_7;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_7;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_7;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_7;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_8;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_8;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_8;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_8;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_8;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_8;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_8;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_8;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_8;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_8;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_8;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_8;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_8;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_8;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_9;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_9;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_9;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_9;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_9;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_9;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_9;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_9;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_9;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_9;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_9;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_9;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_9;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_9;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_10;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_10;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_10;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_10;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_10;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_10;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_10;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_10;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_10;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_10;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_10;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_10;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_10;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_10;
  wire                system_plic_logic_bmb_cmd_valid;
  wire                system_plic_logic_bmb_cmd_ready;
  wire                system_plic_logic_bmb_cmd_payload_last;
  wire       [0:0]    system_plic_logic_bmb_cmd_payload_fragment_opcode;
  wire       [21:0]   system_plic_logic_bmb_cmd_payload_fragment_address;
  wire       [1:0]    system_plic_logic_bmb_cmd_payload_fragment_length;
  wire       [31:0]   system_plic_logic_bmb_cmd_payload_fragment_data;
  wire       [48:0]   system_plic_logic_bmb_cmd_payload_fragment_context;
  wire                system_plic_logic_bmb_rsp_valid;
  wire                system_plic_logic_bmb_rsp_ready;
  wire                system_plic_logic_bmb_rsp_payload_last;
  wire       [0:0]    system_plic_logic_bmb_rsp_payload_fragment_opcode;
  wire       [31:0]   system_plic_logic_bmb_rsp_payload_fragment_data;
  wire       [48:0]   system_plic_logic_bmb_rsp_payload_fragment_context;
  wire                system_plic_logic_bus_readErrorFlag;
  wire                system_plic_logic_bus_writeErrorFlag;
  reg                 system_plic_logic_bus_readHaltTrigger;
  wire                system_plic_logic_bus_writeHaltTrigger;
  wire                system_plic_logic_bus_rsp_valid;
  wire                system_plic_logic_bus_rsp_ready;
  wire                system_plic_logic_bus_rsp_payload_last;
  reg        [0:0]    system_plic_logic_bus_rsp_payload_fragment_opcode;
  reg        [31:0]   system_plic_logic_bus_rsp_payload_fragment_data;
  wire       [48:0]   system_plic_logic_bus_rsp_payload_fragment_context;
  wire                _zz_system_plic_logic_bus_rsp_ready;
  reg                 _zz_system_plic_logic_bus_rsp_ready_1;
  wire                _zz_system_plic_logic_bmb_rsp_valid;
  reg                 _zz_system_plic_logic_bmb_rsp_valid_1;
  reg                 _zz_system_plic_logic_bmb_rsp_payload_last;
  reg        [0:0]    _zz_system_plic_logic_bmb_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_system_plic_logic_bmb_rsp_payload_fragment_data;
  reg        [48:0]   _zz_system_plic_logic_bmb_rsp_payload_fragment_context;
  wire                when_Stream_l375_58;
  wire                system_plic_logic_bus_askWrite;
  wire                system_plic_logic_bus_askRead;
  wire                system_plic_logic_bmb_cmd_fire;
  wire                system_plic_logic_bus_doWrite;
  wire                system_plic_logic_bus_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  wire                system_cores_0_externalInterrupt_plic_target_ie_0;
  wire                system_cores_0_externalInterrupt_plic_target_ie_1;
  wire                system_cores_0_externalInterrupt_plic_target_ie_2;
  wire                system_cores_0_externalInterrupt_plic_target_ie_3;
  wire                system_cores_0_externalInterrupt_plic_target_ie_4;
  wire                system_cores_0_externalInterrupt_plic_target_ie_5;
  wire                system_cores_0_externalInterrupt_plic_target_ie_6;
  wire                system_cores_0_externalInterrupt_plic_target_ie_7;
  wire                system_cores_0_externalInterrupt_plic_target_ie_8;
  wire                system_cores_0_externalInterrupt_plic_target_ie_9;
  wire                system_cores_0_externalInterrupt_plic_target_ie_10;
  wire                system_cores_0_externalInterrupt_plic_target_ie_11;
  wire                system_cores_0_externalInterrupt_plic_target_ie_12;
  wire                system_cores_0_externalInterrupt_plic_target_ie_13;
  wire                system_cores_0_externalInterrupt_plic_target_ie_14;
  wire                system_cores_0_externalInterrupt_plic_target_ie_15;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_threshold;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_0_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_0_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_0_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_1_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_1_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_1_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_2_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_2_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_2_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_3_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_3_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_3_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_4_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_4_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_4_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_5_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_5_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_5_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_6_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_6_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_6_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_7_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_7_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_7_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_8_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_8_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_8_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_9_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_9_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_9_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_10_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_10_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_10_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_11_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_11_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_11_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_12_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_12_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_12_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_13_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_13_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_13_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_14_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_14_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_14_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_15_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_15_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_15_valid;
  wire       [1:0]    system_cores_0_externalInterrupt_plic_target_requests_16_priority;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_requests_16_id;
  wire                system_cores_0_externalInterrupt_plic_target_requests_16_valid;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_1;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_2;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_3;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_4;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_5;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_6;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_7;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_8;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_9;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_10;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_11;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_12;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_13;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_14;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_15;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_16;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_17;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_18;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_19;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_20;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_21;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_22;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_23;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_24;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_25;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_26;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_27;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_28;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_29;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_30;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_31;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_32;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_33;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_34;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_35;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_36;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_37;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_38;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_1;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_39;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_40;
  wire       [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_2;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_valid;
  wire                _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_3;
  reg        [1:0]    system_cores_0_externalInterrupt_plic_target_bestRequest_priority;
  reg        [5:0]    system_cores_0_externalInterrupt_plic_target_bestRequest_id;
  reg                 system_cores_0_externalInterrupt_plic_target_bestRequest_valid;
  wire                system_cores_0_externalInterrupt_plic_target_iep;
  wire       [5:0]    system_cores_0_externalInterrupt_plic_target_claim;
  wire                system_cores_1_externalInterrupt_plic_target_ie_0;
  wire                system_cores_1_externalInterrupt_plic_target_ie_1;
  wire                system_cores_1_externalInterrupt_plic_target_ie_2;
  wire                system_cores_1_externalInterrupt_plic_target_ie_3;
  wire                system_cores_1_externalInterrupt_plic_target_ie_4;
  wire                system_cores_1_externalInterrupt_plic_target_ie_5;
  wire                system_cores_1_externalInterrupt_plic_target_ie_6;
  wire                system_cores_1_externalInterrupt_plic_target_ie_7;
  wire                system_cores_1_externalInterrupt_plic_target_ie_8;
  wire                system_cores_1_externalInterrupt_plic_target_ie_9;
  wire                system_cores_1_externalInterrupt_plic_target_ie_10;
  wire                system_cores_1_externalInterrupt_plic_target_ie_11;
  wire                system_cores_1_externalInterrupt_plic_target_ie_12;
  wire                system_cores_1_externalInterrupt_plic_target_ie_13;
  wire                system_cores_1_externalInterrupt_plic_target_ie_14;
  wire                system_cores_1_externalInterrupt_plic_target_ie_15;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_threshold;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_0_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_0_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_0_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_1_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_1_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_1_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_2_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_2_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_2_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_3_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_3_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_3_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_4_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_4_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_4_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_5_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_5_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_5_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_6_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_6_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_6_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_7_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_7_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_7_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_8_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_8_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_8_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_9_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_9_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_9_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_10_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_10_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_10_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_11_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_11_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_11_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_12_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_12_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_12_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_13_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_13_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_13_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_14_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_14_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_14_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_15_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_15_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_15_valid;
  wire       [1:0]    system_cores_1_externalInterrupt_plic_target_requests_16_priority;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_requests_16_id;
  wire                system_cores_1_externalInterrupt_plic_target_requests_16_valid;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_1;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_2;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_3;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_4;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_5;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_6;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_7;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_8;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_9;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_10;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_11;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_12;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_13;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_14;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_15;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_16;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_17;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_18;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_19;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_20;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_21;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_22;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_23;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_24;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_25;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_26;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_27;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_28;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_29;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_30;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_31;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_32;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_33;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_34;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_35;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_36;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_37;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_38;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_1;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_39;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_40;
  wire       [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_2;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_valid;
  wire                _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_3;
  reg        [1:0]    system_cores_1_externalInterrupt_plic_target_bestRequest_priority;
  reg        [5:0]    system_cores_1_externalInterrupt_plic_target_bestRequest_id;
  reg                 system_cores_1_externalInterrupt_plic_target_bestRequest_valid;
  wire                system_cores_1_externalInterrupt_plic_target_iep;
  wire       [5:0]    system_cores_1_externalInterrupt_plic_target_claim;
  reg        [1:0]    _zz_userInterruptA_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_userInterruptD_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_userInterruptC_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_userInterruptB_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_axiA_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_uart_0_io_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_spi_0_io_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_spi_1_io_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_i2c_0_io_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_i2c_2_io_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_i2c_1_io_interrupt_plic_gateway_priority;
  reg        [1:0]    _zz_system_userTimer_1_interrupts_0_plic_gateway_priority;
  reg        [1:0]    _zz_system_userTimer_0_interrupts_0_plic_gateway_priority;
  reg        [1:0]    _zz_system_gpio_0_io_interrupts_0_plic_gateway_priority;
  reg        [1:0]    _zz_system_gpio_0_io_interrupts_1_plic_gateway_priority;
  reg        [1:0]    _zz_system_watchdog_logic_panics_0_plic_gateway_priority;
  reg                 system_plic_logic_bridge_claim_valid;
  reg        [5:0]    system_plic_logic_bridge_claim_payload;
  reg                 system_plic_logic_bridge_completion_valid;
  reg        [5:0]    system_plic_logic_bridge_completion_payload;
  reg                 system_plic_logic_bridge_coherencyStall_willIncrement;
  wire                system_plic_logic_bridge_coherencyStall_willClear;
  reg        [0:0]    system_plic_logic_bridge_coherencyStall_valueNext;
  reg        [0:0]    system_plic_logic_bridge_coherencyStall_value;
  wire                system_plic_logic_bridge_coherencyStall_willOverflowIfInc;
  wire                system_plic_logic_bridge_coherencyStall_willOverflow;
  wire                when_PlicMapper_l122;
  reg        [1:0]    _zz_system_cores_0_externalInterrupt_plic_target_threshold;
  reg                 system_plic_logic_bridge_targetMapping_0_targetCompletion_valid;
  wire       [5:0]    system_plic_logic_bridge_targetMapping_0_targetCompletion_payload;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_0;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_1;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_2;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_3;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_4;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_5;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_6;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_7;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_8;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_9;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_10;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_11;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_12;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_13;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_14;
  reg                 _zz_system_cores_0_externalInterrupt_plic_target_ie_15;
  reg        [1:0]    _zz_system_cores_1_externalInterrupt_plic_target_threshold;
  reg                 system_plic_logic_bridge_targetMapping_1_targetCompletion_valid;
  wire       [5:0]    system_plic_logic_bridge_targetMapping_1_targetCompletion_payload;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_0;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_1;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_2;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_3;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_4;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_5;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_6;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_7;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_8;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_9;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_10;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_11;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_12;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_13;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_14;
  reg                 _zz_system_cores_1_externalInterrupt_plic_target_ie_15;
  reg                 system_cores_0_externalInterrupt_plic_target_iep_regNext;
  reg                 system_cores_1_externalInterrupt_plic_target_iep_regNext;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_11;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_11;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_11;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_11;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_11;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_11;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_11;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_11;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_11;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_11;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_11;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_11;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_11;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_11;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_12;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_12;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_12;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_12;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_12;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_12;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_12;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_12;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_12;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_12;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_12;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_12;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_12;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_12;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_13;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_13;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_13;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_13;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_13;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_13;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_13;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_13;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_13;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_13;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_13;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_13;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_13;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_13;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_14;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_14;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_14;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_14;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_14;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_14;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_14;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_14;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_14;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_14;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_14;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_14;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_14;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_14;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_15;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_15;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_15;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_15;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_15;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_15;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_15;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_15;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_15;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_15;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_15;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_15;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_15;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_15;
  wire                system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  wire                system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  wire                system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  wire       [0:0]    system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  wire       [21:0]   system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  wire       [1:0]    system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  wire       [31:0]   system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  wire       [48:0]   system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  wire                system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  wire                system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  wire                system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  wire       [0:0]    system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  wire       [31:0]   system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  wire       [48:0]   system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_valid_16;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_ready_16;
  wire                system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_16;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_16;
  wire       [23:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_16;
  wire       [1:0]    system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_16;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_16;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_16;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_valid_16;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_ready_16;
  wire                system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_16;
  wire       [0:0]    system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_16;
  wire       [31:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_16;
  wire       [48:0]   system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_16;
  wire                when_BmbSlaveFactory_l77;
  `ifndef SYNTHESIS
  reg [71:0] system_cores_0_debugRiscv_dmToHart_payload_op_string;
  reg [71:0] system_cores_1_debugRiscv_dmToHart_payload_op_string;
  reg [63:0] FpuPlugin_port_commit_m2sPipe_payload_opcode_string;
  reg [63:0] FpuPlugin_port_commit_rData_opcode_string;
  reg [63:0] FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string;
  reg [63:0] FpuPlugin_port_commit_rData_opcode_1_string;
  reg [71:0] io_harts_0_dmToHart_regNext_payload_op_string;
  reg [71:0] io_harts_1_dmToHart_regNext_payload_op_string;
  `endif


  assign io_ddrMasters_1_reset = io_ddrMasters_1_reset_read_buffer;
  assign io_ddrMasters_0_reset = io_ddrMasters_0_reset_read_buffer;
  assign _zz_dBus_inv_payload_fragment_address_1 = 6'h0;
  assign _zz_dBus_inv_payload_fragment_address = {26'd0, _zz_dBus_inv_payload_fragment_address_1};
  assign _zz_dBus_inv_payload_fragment_address_3 = 6'h0;
  assign _zz_dBus_inv_payload_fragment_address_2 = {26'd0, _zz_dBus_inv_payload_fragment_address_3};
  VexRiscv system_cores_0_logic_cpu (
    .dBus_cmd_valid                             (system_cores_0_logic_cpu_dBus_cmd_valid                                     ), //o
    .dBus_cmd_ready                             (_zz_dBus_cmd_ready                                                          ), //i
    .dBus_cmd_payload_wr                        (system_cores_0_logic_cpu_dBus_cmd_payload_wr                                ), //o
    .dBus_cmd_payload_uncached                  (system_cores_0_logic_cpu_dBus_cmd_payload_uncached                          ), //o
    .dBus_cmd_payload_address                   (system_cores_0_logic_cpu_dBus_cmd_payload_address[31:0]                     ), //o
    .dBus_cmd_payload_data                      (system_cores_0_logic_cpu_dBus_cmd_payload_data[63:0]                        ), //o
    .dBus_cmd_payload_mask                      (system_cores_0_logic_cpu_dBus_cmd_payload_mask[7:0]                         ), //o
    .dBus_cmd_payload_size                      (system_cores_0_logic_cpu_dBus_cmd_payload_size[2:0]                         ), //o
    .dBus_cmd_payload_exclusive                 (system_cores_0_logic_cpu_dBus_cmd_payload_exclusive                         ), //o
    .dBus_cmd_payload_last                      (system_cores_0_logic_cpu_dBus_cmd_payload_last                              ), //o
    .dBus_rsp_valid                             (dBus_Bridge_bus_rsp_valid                                                   ), //i
    .dBus_rsp_payload_aggregated                (dBus_Bridge_withWriteBuffer_rspCtx_rspCount[3:0]                            ), //i
    .dBus_rsp_payload_last                      (dBus_Bridge_bus_rsp_payload_last                                            ), //i
    .dBus_rsp_payload_data                      (dBus_Bridge_bus_rsp_payload_fragment_data[63:0]                             ), //i
    .dBus_rsp_payload_error                     (system_cores_0_logic_cpu_dBus_rsp_payload_error                             ), //i
    .dBus_rsp_payload_exclusive                 (dBus_Bridge_bus_rsp_payload_fragment_exclusive                              ), //i
    .dBus_inv_valid                             (dBus_Bridge_bus_inv_valid                                                   ), //i
    .dBus_inv_ready                             (system_cores_0_logic_cpu_dBus_inv_ready                                     ), //o
    .dBus_inv_payload_last                      (system_cores_0_logic_cpu_dBus_inv_payload_last                              ), //i
    .dBus_inv_payload_fragment_enable           (dBus_Bridge_bus_inv_payload_all                                             ), //i
    .dBus_inv_payload_fragment_address          (system_cores_0_logic_cpu_dBus_inv_payload_fragment_address[31:0]            ), //i
    .dBus_ack_valid                             (system_cores_0_logic_cpu_dBus_ack_valid                                     ), //o
    .dBus_ack_ready                             (system_cores_0_logic_cpu_dBus_ack_ready                                     ), //i
    .dBus_ack_payload_last                      (system_cores_0_logic_cpu_dBus_ack_payload_last                              ), //o
    .dBus_ack_payload_fragment_hit              (system_cores_0_logic_cpu_dBus_ack_payload_fragment_hit                      ), //o
    .dBus_sync_valid                            (dBus_Bridge_bus_sync_valid                                                  ), //i
    .dBus_sync_ready                            (system_cores_0_logic_cpu_dBus_sync_ready                                    ), //o
    .dBus_sync_payload_aggregated               (dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_payload[3:0]                  ), //i
    .timerInterrupt                             (bufferCC_74_io_dataOut                                                      ), //i
    .externalInterrupt                          (system_cores_0_externalInterrupt_plic_target_iep_regNext_buffercc_io_dataOut), //i
    .softwareInterrupt                          (bufferCC_75_io_dataOut                                                      ), //i
    .debugBus_halted                            (system_cores_0_logic_cpu_debugBus_halted                                    ), //o
    .debugBus_running                           (system_cores_0_logic_cpu_debugBus_running                                   ), //o
    .debugBus_unavailable                       (system_cores_0_logic_cpu_debugBus_unavailable                               ), //o
    .debugBus_exception                         (system_cores_0_logic_cpu_debugBus_exception                                 ), //o
    .debugBus_commit                            (system_cores_0_logic_cpu_debugBus_commit                                    ), //o
    .debugBus_ebreak                            (system_cores_0_logic_cpu_debugBus_ebreak                                    ), //o
    .debugBus_redo                              (system_cores_0_logic_cpu_debugBus_redo                                      ), //o
    .debugBus_regSuccess                        (system_cores_0_logic_cpu_debugBus_regSuccess                                ), //o
    .debugBus_ackReset                          (system_cores_0_debugRiscv_ackReset                                          ), //i
    .debugBus_haveReset                         (system_cores_0_logic_cpu_debugBus_haveReset                                 ), //o
    .debugBus_resume_cmd_valid                  (system_cores_0_debugRiscv_resume_cmd_valid                                  ), //i
    .debugBus_resume_rsp_valid                  (system_cores_0_logic_cpu_debugBus_resume_rsp_valid                          ), //o
    .debugBus_haltReq                           (system_cores_0_debugRiscv_haltReq                                           ), //i
    .debugBus_dmToHart_valid                    (system_cores_0_debugRiscv_dmToHart_valid                                    ), //i
    .debugBus_dmToHart_payload_op               (system_cores_0_debugRiscv_dmToHart_payload_op[1:0]                          ), //i
    .debugBus_dmToHart_payload_address          (system_cores_0_debugRiscv_dmToHart_payload_address[4:0]                     ), //i
    .debugBus_dmToHart_payload_data             (system_cores_0_debugRiscv_dmToHart_payload_data[31:0]                       ), //i
    .debugBus_dmToHart_payload_size             (system_cores_0_debugRiscv_dmToHart_payload_size[2:0]                        ), //i
    .debugBus_hartToDm_valid                    (system_cores_0_logic_cpu_debugBus_hartToDm_valid                            ), //o
    .debugBus_hartToDm_payload_address          (system_cores_0_logic_cpu_debugBus_hartToDm_payload_address[3:0]             ), //o
    .debugBus_hartToDm_payload_data             (system_cores_0_logic_cpu_debugBus_hartToDm_payload_data[31:0]               ), //o
    .FpuPlugin_port_cmd_valid                   (system_cores_0_logic_cpu_FpuPlugin_port_cmd_valid                           ), //o
    .FpuPlugin_port_cmd_ready                   (system_fpu_logic_io_port_0_cmd_ready                                        ), //i
    .FpuPlugin_port_cmd_payload_opcode          (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_opcode[3:0]             ), //o
    .FpuPlugin_port_cmd_payload_arg             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_arg[1:0]                ), //o
    .FpuPlugin_port_cmd_payload_rs1             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs1[4:0]                ), //o
    .FpuPlugin_port_cmd_payload_rs2             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs2[4:0]                ), //o
    .FpuPlugin_port_cmd_payload_rs3             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs3[4:0]                ), //o
    .FpuPlugin_port_cmd_payload_rd              (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rd[4:0]                 ), //o
    .FpuPlugin_port_cmd_payload_format          (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_format                  ), //o
    .FpuPlugin_port_cmd_payload_roundMode       (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_roundMode[2:0]          ), //o
    .FpuPlugin_port_commit_valid                (system_cores_0_logic_cpu_FpuPlugin_port_commit_valid                        ), //o
    .FpuPlugin_port_commit_ready                (system_cores_0_logic_cpu_FpuPlugin_port_commit_ready                        ), //i
    .FpuPlugin_port_commit_payload_opcode       (system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_opcode[3:0]          ), //o
    .FpuPlugin_port_commit_payload_rd           (system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_rd[4:0]              ), //o
    .FpuPlugin_port_commit_payload_write        (system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_write                ), //o
    .FpuPlugin_port_commit_payload_value        (system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_value[63:0]          ), //o
    .FpuPlugin_port_rsp_valid                   (io_port_0_rsp_s2mPipe_valid                                                 ), //i
    .FpuPlugin_port_rsp_ready                   (system_cores_0_logic_cpu_FpuPlugin_port_rsp_ready                           ), //o
    .FpuPlugin_port_rsp_payload_value           (io_port_0_rsp_s2mPipe_payload_value[63:0]                                   ), //i
    .FpuPlugin_port_rsp_payload_NV              (io_port_0_rsp_s2mPipe_payload_NV                                            ), //i
    .FpuPlugin_port_rsp_payload_NX              (io_port_0_rsp_s2mPipe_payload_NX                                            ), //i
    .FpuPlugin_port_completion_valid            (io_port_0_completion_regNext_valid                                          ), //i
    .FpuPlugin_port_completion_payload_flags_NX (io_port_0_completion_regNext_payload_flags_NX                               ), //i
    .FpuPlugin_port_completion_payload_flags_UF (io_port_0_completion_regNext_payload_flags_UF                               ), //i
    .FpuPlugin_port_completion_payload_flags_OF (io_port_0_completion_regNext_payload_flags_OF                               ), //i
    .FpuPlugin_port_completion_payload_flags_DZ (io_port_0_completion_regNext_payload_flags_DZ                               ), //i
    .FpuPlugin_port_completion_payload_flags_NV (io_port_0_completion_regNext_payload_flags_NV                               ), //i
    .FpuPlugin_port_completion_payload_written  (io_port_0_completion_regNext_payload_written                                ), //i
    .CfuPlugin_bus_cmd_valid                    (system_cores_0_logic_cpu_CfuPlugin_bus_cmd_valid                            ), //o
    .CfuPlugin_bus_cmd_ready                    (cpu0_customInstruction_cmd_ready                                            ), //i
    .CfuPlugin_bus_cmd_payload_function_id      (system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_function_id[9:0]         ), //o
    .CfuPlugin_bus_cmd_payload_inputs_0         (system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_0[31:0]           ), //o
    .CfuPlugin_bus_cmd_payload_inputs_1         (system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_1[31:0]           ), //o
    .CfuPlugin_bus_rsp_valid                    (cpu0_customInstruction_rsp_valid                                            ), //i
    .CfuPlugin_bus_rsp_ready                    (system_cores_0_logic_cpu_CfuPlugin_bus_rsp_ready                            ), //o
    .CfuPlugin_bus_rsp_payload_outputs_0        (cpu0_customInstruction_outputs_0[31:0]                                      ), //i
    .iBus_cmd_valid                             (system_cores_0_logic_cpu_iBus_cmd_valid                                     ), //o
    .iBus_cmd_ready                             (system_cores_0_iBus_cmd_ready                                               ), //i
    .iBus_cmd_payload_address                   (system_cores_0_logic_cpu_iBus_cmd_payload_address[31:0]                     ), //o
    .iBus_cmd_payload_size                      (system_cores_0_logic_cpu_iBus_cmd_payload_size[2:0]                         ), //o
    .iBus_rsp_valid                             (system_cores_0_iBus_rsp_valid                                               ), //i
    .iBus_rsp_payload_data                      (system_cores_0_iBus_rsp_payload_fragment_data[63:0]                         ), //i
    .iBus_rsp_payload_error                     (system_cores_0_logic_cpu_iBus_rsp_payload_error                             ), //i
    .systemCd_logic_outputReset                 (systemCd_logic_outputReset                                                  ), //i
    .stoptime                                   (system_cores_0_logic_cpu_stoptime                                           ), //o
    .io_systemClk                               (io_systemClk                                                                )  //i
  );
  VexRiscv_1 system_cores_1_logic_cpu (
    .dBus_cmd_valid                             (system_cores_1_logic_cpu_dBus_cmd_valid                                     ), //o
    .dBus_cmd_ready                             (_zz_dBus_cmd_ready_1                                                        ), //i
    .dBus_cmd_payload_wr                        (system_cores_1_logic_cpu_dBus_cmd_payload_wr                                ), //o
    .dBus_cmd_payload_uncached                  (system_cores_1_logic_cpu_dBus_cmd_payload_uncached                          ), //o
    .dBus_cmd_payload_address                   (system_cores_1_logic_cpu_dBus_cmd_payload_address[31:0]                     ), //o
    .dBus_cmd_payload_data                      (system_cores_1_logic_cpu_dBus_cmd_payload_data[63:0]                        ), //o
    .dBus_cmd_payload_mask                      (system_cores_1_logic_cpu_dBus_cmd_payload_mask[7:0]                         ), //o
    .dBus_cmd_payload_size                      (system_cores_1_logic_cpu_dBus_cmd_payload_size[2:0]                         ), //o
    .dBus_cmd_payload_exclusive                 (system_cores_1_logic_cpu_dBus_cmd_payload_exclusive                         ), //o
    .dBus_cmd_payload_last                      (system_cores_1_logic_cpu_dBus_cmd_payload_last                              ), //o
    .dBus_rsp_valid                             (dBus_Bridge_bus_rsp_valid_1                                                 ), //i
    .dBus_rsp_payload_aggregated                (dBus_Bridge_withWriteBuffer_rspCtx_rspCount_1[3:0]                          ), //i
    .dBus_rsp_payload_last                      (dBus_Bridge_bus_rsp_payload_last_1                                          ), //i
    .dBus_rsp_payload_data                      (dBus_Bridge_bus_rsp_payload_fragment_data_1[63:0]                           ), //i
    .dBus_rsp_payload_error                     (system_cores_1_logic_cpu_dBus_rsp_payload_error                             ), //i
    .dBus_rsp_payload_exclusive                 (dBus_Bridge_bus_rsp_payload_fragment_exclusive_1                            ), //i
    .dBus_inv_valid                             (dBus_Bridge_bus_inv_valid_1                                                 ), //i
    .dBus_inv_ready                             (system_cores_1_logic_cpu_dBus_inv_ready                                     ), //o
    .dBus_inv_payload_last                      (system_cores_1_logic_cpu_dBus_inv_payload_last                              ), //i
    .dBus_inv_payload_fragment_enable           (dBus_Bridge_bus_inv_payload_all_1                                           ), //i
    .dBus_inv_payload_fragment_address          (system_cores_1_logic_cpu_dBus_inv_payload_fragment_address[31:0]            ), //i
    .dBus_ack_valid                             (system_cores_1_logic_cpu_dBus_ack_valid                                     ), //o
    .dBus_ack_ready                             (system_cores_1_logic_cpu_dBus_ack_ready                                     ), //i
    .dBus_ack_payload_last                      (system_cores_1_logic_cpu_dBus_ack_payload_last                              ), //o
    .dBus_ack_payload_fragment_hit              (system_cores_1_logic_cpu_dBus_ack_payload_fragment_hit                      ), //o
    .dBus_sync_valid                            (dBus_Bridge_bus_sync_valid_1                                                ), //i
    .dBus_sync_ready                            (system_cores_1_logic_cpu_dBus_sync_ready                                    ), //o
    .dBus_sync_payload_aggregated               (dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_payload_1[3:0]                ), //i
    .timerInterrupt                             (bufferCC_76_io_dataOut                                                      ), //i
    .externalInterrupt                          (system_cores_1_externalInterrupt_plic_target_iep_regNext_buffercc_io_dataOut), //i
    .softwareInterrupt                          (bufferCC_77_io_dataOut                                                      ), //i
    .debugBus_halted                            (system_cores_1_logic_cpu_debugBus_halted                                    ), //o
    .debugBus_running                           (system_cores_1_logic_cpu_debugBus_running                                   ), //o
    .debugBus_unavailable                       (system_cores_1_logic_cpu_debugBus_unavailable                               ), //o
    .debugBus_exception                         (system_cores_1_logic_cpu_debugBus_exception                                 ), //o
    .debugBus_commit                            (system_cores_1_logic_cpu_debugBus_commit                                    ), //o
    .debugBus_ebreak                            (system_cores_1_logic_cpu_debugBus_ebreak                                    ), //o
    .debugBus_redo                              (system_cores_1_logic_cpu_debugBus_redo                                      ), //o
    .debugBus_regSuccess                        (system_cores_1_logic_cpu_debugBus_regSuccess                                ), //o
    .debugBus_ackReset                          (system_cores_1_debugRiscv_ackReset                                          ), //i
    .debugBus_haveReset                         (system_cores_1_logic_cpu_debugBus_haveReset                                 ), //o
    .debugBus_resume_cmd_valid                  (system_cores_1_debugRiscv_resume_cmd_valid                                  ), //i
    .debugBus_resume_rsp_valid                  (system_cores_1_logic_cpu_debugBus_resume_rsp_valid                          ), //o
    .debugBus_haltReq                           (system_cores_1_debugRiscv_haltReq                                           ), //i
    .debugBus_dmToHart_valid                    (system_cores_1_debugRiscv_dmToHart_valid                                    ), //i
    .debugBus_dmToHart_payload_op               (system_cores_1_debugRiscv_dmToHart_payload_op[1:0]                          ), //i
    .debugBus_dmToHart_payload_address          (system_cores_1_debugRiscv_dmToHart_payload_address[4:0]                     ), //i
    .debugBus_dmToHart_payload_data             (system_cores_1_debugRiscv_dmToHart_payload_data[31:0]                       ), //i
    .debugBus_dmToHart_payload_size             (system_cores_1_debugRiscv_dmToHart_payload_size[2:0]                        ), //i
    .debugBus_hartToDm_valid                    (system_cores_1_logic_cpu_debugBus_hartToDm_valid                            ), //o
    .debugBus_hartToDm_payload_address          (system_cores_1_logic_cpu_debugBus_hartToDm_payload_address[3:0]             ), //o
    .debugBus_hartToDm_payload_data             (system_cores_1_logic_cpu_debugBus_hartToDm_payload_data[31:0]               ), //o
    .FpuPlugin_port_cmd_valid                   (system_cores_1_logic_cpu_FpuPlugin_port_cmd_valid                           ), //o
    .FpuPlugin_port_cmd_ready                   (system_fpu_logic_io_port_1_cmd_ready                                        ), //i
    .FpuPlugin_port_cmd_payload_opcode          (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_opcode[3:0]             ), //o
    .FpuPlugin_port_cmd_payload_arg             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_arg[1:0]                ), //o
    .FpuPlugin_port_cmd_payload_rs1             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs1[4:0]                ), //o
    .FpuPlugin_port_cmd_payload_rs2             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs2[4:0]                ), //o
    .FpuPlugin_port_cmd_payload_rs3             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs3[4:0]                ), //o
    .FpuPlugin_port_cmd_payload_rd              (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rd[4:0]                 ), //o
    .FpuPlugin_port_cmd_payload_format          (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_format                  ), //o
    .FpuPlugin_port_cmd_payload_roundMode       (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_roundMode[2:0]          ), //o
    .FpuPlugin_port_commit_valid                (system_cores_1_logic_cpu_FpuPlugin_port_commit_valid                        ), //o
    .FpuPlugin_port_commit_ready                (system_cores_1_logic_cpu_FpuPlugin_port_commit_ready                        ), //i
    .FpuPlugin_port_commit_payload_opcode       (system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_opcode[3:0]          ), //o
    .FpuPlugin_port_commit_payload_rd           (system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_rd[4:0]              ), //o
    .FpuPlugin_port_commit_payload_write        (system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_write                ), //o
    .FpuPlugin_port_commit_payload_value        (system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_value[63:0]          ), //o
    .FpuPlugin_port_rsp_valid                   (io_port_1_rsp_s2mPipe_valid                                                 ), //i
    .FpuPlugin_port_rsp_ready                   (system_cores_1_logic_cpu_FpuPlugin_port_rsp_ready                           ), //o
    .FpuPlugin_port_rsp_payload_value           (io_port_1_rsp_s2mPipe_payload_value[63:0]                                   ), //i
    .FpuPlugin_port_rsp_payload_NV              (io_port_1_rsp_s2mPipe_payload_NV                                            ), //i
    .FpuPlugin_port_rsp_payload_NX              (io_port_1_rsp_s2mPipe_payload_NX                                            ), //i
    .FpuPlugin_port_completion_valid            (io_port_1_completion_regNext_valid                                          ), //i
    .FpuPlugin_port_completion_payload_flags_NX (io_port_1_completion_regNext_payload_flags_NX                               ), //i
    .FpuPlugin_port_completion_payload_flags_UF (io_port_1_completion_regNext_payload_flags_UF                               ), //i
    .FpuPlugin_port_completion_payload_flags_OF (io_port_1_completion_regNext_payload_flags_OF                               ), //i
    .FpuPlugin_port_completion_payload_flags_DZ (io_port_1_completion_regNext_payload_flags_DZ                               ), //i
    .FpuPlugin_port_completion_payload_flags_NV (io_port_1_completion_regNext_payload_flags_NV                               ), //i
    .FpuPlugin_port_completion_payload_written  (io_port_1_completion_regNext_payload_written                                ), //i
    .CfuPlugin_bus_cmd_valid                    (system_cores_1_logic_cpu_CfuPlugin_bus_cmd_valid                            ), //o
    .CfuPlugin_bus_cmd_ready                    (cpu1_customInstruction_cmd_ready                                            ), //i
    .CfuPlugin_bus_cmd_payload_function_id      (system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_function_id[9:0]         ), //o
    .CfuPlugin_bus_cmd_payload_inputs_0         (system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_0[31:0]           ), //o
    .CfuPlugin_bus_cmd_payload_inputs_1         (system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_1[31:0]           ), //o
    .CfuPlugin_bus_rsp_valid                    (cpu1_customInstruction_rsp_valid                                            ), //i
    .CfuPlugin_bus_rsp_ready                    (system_cores_1_logic_cpu_CfuPlugin_bus_rsp_ready                            ), //o
    .CfuPlugin_bus_rsp_payload_outputs_0        (cpu1_customInstruction_outputs_0[31:0]                                      ), //i
    .iBus_cmd_valid                             (system_cores_1_logic_cpu_iBus_cmd_valid                                     ), //o
    .iBus_cmd_ready                             (system_cores_1_iBus_cmd_ready                                               ), //i
    .iBus_cmd_payload_address                   (system_cores_1_logic_cpu_iBus_cmd_payload_address[31:0]                     ), //o
    .iBus_cmd_payload_size                      (system_cores_1_logic_cpu_iBus_cmd_payload_size[2:0]                         ), //o
    .iBus_rsp_valid                             (system_cores_1_iBus_rsp_valid                                               ), //i
    .iBus_rsp_payload_data                      (system_cores_1_iBus_rsp_payload_fragment_data[63:0]                         ), //i
    .iBus_rsp_payload_error                     (system_cores_1_logic_cpu_iBus_rsp_payload_error                             ), //i
    .systemCd_logic_outputReset                 (systemCd_logic_outputReset                                                  ), //i
    .stoptime                                   (system_cores_1_logic_cpu_stoptime                                           ), //o
    .io_systemClk                               (io_systemClk                                                                )  //i
  );
  FpuCore system_fpu_logic (
    .io_port_0_cmd_valid                   (system_cores_0_logic_cpu_FpuPlugin_port_cmd_valid                 ), //i
    .io_port_0_cmd_ready                   (system_fpu_logic_io_port_0_cmd_ready                              ), //o
    .io_port_0_cmd_payload_opcode          (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_opcode[3:0]   ), //i
    .io_port_0_cmd_payload_arg             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_arg[1:0]      ), //i
    .io_port_0_cmd_payload_rs1             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs1[4:0]      ), //i
    .io_port_0_cmd_payload_rs2             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs2[4:0]      ), //i
    .io_port_0_cmd_payload_rs3             (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rs3[4:0]      ), //i
    .io_port_0_cmd_payload_rd              (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_rd[4:0]       ), //i
    .io_port_0_cmd_payload_format          (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_format        ), //i
    .io_port_0_cmd_payload_roundMode       (system_cores_0_logic_cpu_FpuPlugin_port_cmd_payload_roundMode[2:0]), //i
    .io_port_0_commit_valid                (FpuPlugin_port_commit_m2sPipe_valid                               ), //i
    .io_port_0_commit_ready                (system_fpu_logic_io_port_0_commit_ready                           ), //o
    .io_port_0_commit_payload_opcode       (FpuPlugin_port_commit_m2sPipe_payload_opcode[3:0]                 ), //i
    .io_port_0_commit_payload_rd           (FpuPlugin_port_commit_m2sPipe_payload_rd[4:0]                     ), //i
    .io_port_0_commit_payload_write        (FpuPlugin_port_commit_m2sPipe_payload_write                       ), //i
    .io_port_0_commit_payload_value        (FpuPlugin_port_commit_m2sPipe_payload_value[63:0]                 ), //i
    .io_port_0_rsp_valid                   (system_fpu_logic_io_port_0_rsp_valid                              ), //o
    .io_port_0_rsp_ready                   (io_port_0_rsp_rValidN                                             ), //i
    .io_port_0_rsp_payload_value           (system_fpu_logic_io_port_0_rsp_payload_value[63:0]                ), //o
    .io_port_0_rsp_payload_NV              (system_fpu_logic_io_port_0_rsp_payload_NV                         ), //o
    .io_port_0_rsp_payload_NX              (system_fpu_logic_io_port_0_rsp_payload_NX                         ), //o
    .io_port_0_completion_valid            (system_fpu_logic_io_port_0_completion_valid                       ), //o
    .io_port_0_completion_payload_flags_NX (system_fpu_logic_io_port_0_completion_payload_flags_NX            ), //o
    .io_port_0_completion_payload_flags_UF (system_fpu_logic_io_port_0_completion_payload_flags_UF            ), //o
    .io_port_0_completion_payload_flags_OF (system_fpu_logic_io_port_0_completion_payload_flags_OF            ), //o
    .io_port_0_completion_payload_flags_DZ (system_fpu_logic_io_port_0_completion_payload_flags_DZ            ), //o
    .io_port_0_completion_payload_flags_NV (system_fpu_logic_io_port_0_completion_payload_flags_NV            ), //o
    .io_port_0_completion_payload_written  (system_fpu_logic_io_port_0_completion_payload_written             ), //o
    .io_port_1_cmd_valid                   (system_cores_1_logic_cpu_FpuPlugin_port_cmd_valid                 ), //i
    .io_port_1_cmd_ready                   (system_fpu_logic_io_port_1_cmd_ready                              ), //o
    .io_port_1_cmd_payload_opcode          (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_opcode[3:0]   ), //i
    .io_port_1_cmd_payload_arg             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_arg[1:0]      ), //i
    .io_port_1_cmd_payload_rs1             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs1[4:0]      ), //i
    .io_port_1_cmd_payload_rs2             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs2[4:0]      ), //i
    .io_port_1_cmd_payload_rs3             (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rs3[4:0]      ), //i
    .io_port_1_cmd_payload_rd              (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_rd[4:0]       ), //i
    .io_port_1_cmd_payload_format          (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_format        ), //i
    .io_port_1_cmd_payload_roundMode       (system_cores_1_logic_cpu_FpuPlugin_port_cmd_payload_roundMode[2:0]), //i
    .io_port_1_commit_valid                (FpuPlugin_port_commit_m2sPipe_valid_1                             ), //i
    .io_port_1_commit_ready                (system_fpu_logic_io_port_1_commit_ready                           ), //o
    .io_port_1_commit_payload_opcode       (FpuPlugin_port_commit_m2sPipe_payload_opcode_1[3:0]               ), //i
    .io_port_1_commit_payload_rd           (FpuPlugin_port_commit_m2sPipe_payload_rd_1[4:0]                   ), //i
    .io_port_1_commit_payload_write        (FpuPlugin_port_commit_m2sPipe_payload_write_1                     ), //i
    .io_port_1_commit_payload_value        (FpuPlugin_port_commit_m2sPipe_payload_value_1[63:0]               ), //i
    .io_port_1_rsp_valid                   (system_fpu_logic_io_port_1_rsp_valid                              ), //o
    .io_port_1_rsp_ready                   (io_port_1_rsp_rValidN                                             ), //i
    .io_port_1_rsp_payload_value           (system_fpu_logic_io_port_1_rsp_payload_value[63:0]                ), //o
    .io_port_1_rsp_payload_NV              (system_fpu_logic_io_port_1_rsp_payload_NV                         ), //o
    .io_port_1_rsp_payload_NX              (system_fpu_logic_io_port_1_rsp_payload_NX                         ), //o
    .io_port_1_completion_valid            (system_fpu_logic_io_port_1_completion_valid                       ), //o
    .io_port_1_completion_payload_flags_NX (system_fpu_logic_io_port_1_completion_payload_flags_NX            ), //o
    .io_port_1_completion_payload_flags_UF (system_fpu_logic_io_port_1_completion_payload_flags_UF            ), //o
    .io_port_1_completion_payload_flags_OF (system_fpu_logic_io_port_1_completion_payload_flags_OF            ), //o
    .io_port_1_completion_payload_flags_DZ (system_fpu_logic_io_port_1_completion_payload_flags_DZ            ), //o
    .io_port_1_completion_payload_flags_NV (system_fpu_logic_io_port_1_completion_payload_flags_NV            ), //o
    .io_port_1_completion_payload_written  (system_fpu_logic_io_port_1_completion_payload_written             ), //o
    .io_systemClk                          (io_systemClk                                                      ), //i
    .systemCd_logic_outputReset            (systemCd_logic_outputReset                                        )  //i
  );
  DebugModule system_riscvJtag_debug_logic_dm (
    .io_ctrl_cmd_valid                   (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_valid                     ), //i
    .io_ctrl_cmd_ready                   (system_riscvJtag_debug_logic_dm_io_ctrl_cmd_ready                       ), //o
    .io_ctrl_cmd_payload_write           (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_write             ), //i
    .io_ctrl_cmd_payload_data            (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_data[31:0]        ), //i
    .io_ctrl_cmd_payload_address         (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_address[6:0]      ), //i
    .io_ctrl_rsp_valid                   (system_riscvJtag_debug_logic_dm_io_ctrl_rsp_valid                       ), //o
    .io_ctrl_rsp_payload_error           (system_riscvJtag_debug_logic_dm_io_ctrl_rsp_payload_error               ), //o
    .io_ctrl_rsp_payload_data            (system_riscvJtag_debug_logic_dm_io_ctrl_rsp_payload_data[31:0]          ), //o
    .io_ndmreset                         (system_riscvJtag_debug_logic_dm_io_ndmreset                             ), //o
    .io_harts_0_halted                   (system_cores_0_debugRiscv_halted                                        ), //i
    .io_harts_0_running                  (system_cores_0_debugRiscv_running                                       ), //i
    .io_harts_0_unavailable              (system_cores_0_debugRiscv_unavailable                                   ), //i
    .io_harts_0_exception                (system_cores_0_debugRiscv_exception                                     ), //i
    .io_harts_0_commit                   (system_cores_0_debugRiscv_commit                                        ), //i
    .io_harts_0_ebreak                   (system_cores_0_debugRiscv_ebreak                                        ), //i
    .io_harts_0_redo                     (system_cores_0_debugRiscv_redo                                          ), //i
    .io_harts_0_regSuccess               (system_cores_0_debugRiscv_regSuccess                                    ), //i
    .io_harts_0_ackReset                 (system_riscvJtag_debug_logic_dm_io_harts_0_ackReset                     ), //o
    .io_harts_0_haveReset                (system_cores_0_debugRiscv_haveReset                                     ), //i
    .io_harts_0_resume_cmd_valid         (system_riscvJtag_debug_logic_dm_io_harts_0_resume_cmd_valid             ), //o
    .io_harts_0_resume_rsp_valid         (system_cores_0_debugRiscv_resume_rsp_valid                              ), //i
    .io_harts_0_haltReq                  (system_riscvJtag_debug_logic_dm_io_harts_0_haltReq                      ), //o
    .io_harts_0_dmToHart_valid           (system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_valid               ), //o
    .io_harts_0_dmToHart_payload_op      (system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_op[1:0]     ), //o
    .io_harts_0_dmToHart_payload_address (system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_address[4:0]), //o
    .io_harts_0_dmToHart_payload_data    (system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_data[31:0]  ), //o
    .io_harts_0_dmToHart_payload_size    (system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_size[2:0]   ), //o
    .io_harts_0_hartToDm_valid           (system_cores_0_debugRiscv_hartToDm_valid                                ), //i
    .io_harts_0_hartToDm_payload_address (system_cores_0_debugRiscv_hartToDm_payload_address[3:0]                 ), //i
    .io_harts_0_hartToDm_payload_data    (system_cores_0_debugRiscv_hartToDm_payload_data[31:0]                   ), //i
    .io_harts_1_halted                   (system_cores_1_debugRiscv_halted                                        ), //i
    .io_harts_1_running                  (system_cores_1_debugRiscv_running                                       ), //i
    .io_harts_1_unavailable              (system_cores_1_debugRiscv_unavailable                                   ), //i
    .io_harts_1_exception                (system_cores_1_debugRiscv_exception                                     ), //i
    .io_harts_1_commit                   (system_cores_1_debugRiscv_commit                                        ), //i
    .io_harts_1_ebreak                   (system_cores_1_debugRiscv_ebreak                                        ), //i
    .io_harts_1_redo                     (system_cores_1_debugRiscv_redo                                          ), //i
    .io_harts_1_regSuccess               (system_cores_1_debugRiscv_regSuccess                                    ), //i
    .io_harts_1_ackReset                 (system_riscvJtag_debug_logic_dm_io_harts_1_ackReset                     ), //o
    .io_harts_1_haveReset                (system_cores_1_debugRiscv_haveReset                                     ), //i
    .io_harts_1_resume_cmd_valid         (system_riscvJtag_debug_logic_dm_io_harts_1_resume_cmd_valid             ), //o
    .io_harts_1_resume_rsp_valid         (system_cores_1_debugRiscv_resume_rsp_valid                              ), //i
    .io_harts_1_haltReq                  (system_riscvJtag_debug_logic_dm_io_harts_1_haltReq                      ), //o
    .io_harts_1_dmToHart_valid           (system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_valid               ), //o
    .io_harts_1_dmToHart_payload_op      (system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_op[1:0]     ), //o
    .io_harts_1_dmToHart_payload_address (system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_address[4:0]), //o
    .io_harts_1_dmToHart_payload_data    (system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_data[31:0]  ), //o
    .io_harts_1_dmToHart_payload_size    (system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_size[2:0]   ), //o
    .io_harts_1_hartToDm_valid           (system_cores_1_debugRiscv_hartToDm_valid                                ), //i
    .io_harts_1_hartToDm_payload_address (system_cores_1_debugRiscv_hartToDm_payload_address[3:0]                 ), //i
    .io_harts_1_hartToDm_payload_data    (system_cores_1_debugRiscv_hartToDm_payload_data[31:0]                   ), //i
    .io_systemClk                        (io_systemClk                                                            ), //i
    .debugCd_logic_outputReset           (debugCd_logic_outputReset                                               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_56 io_asyncReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn     (io_asyncReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut    (io_asyncReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_systemClk  (io_systemClk                                             ), //i
    .io_asyncReset (io_asyncReset                                            )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_57 debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn                 (debugCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut                (debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_memoryClk              (io_memoryClk                                                         ), //i
    .debugCd_logic_outputReset (debugCd_logic_outputReset                                            )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_39 peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn                      (peripheralCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut                     (peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_systemClk                   (io_systemClk                                                              ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                                            )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_59 ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn               (ddrCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut              (ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_peripheralClk        (io_peripheralClk                                                   ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                                            )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_60 userInterruptA_buffercc (
    .io_dataIn                      (userInterruptA                    ), //i
    .io_dataOut                     (userInterruptA_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                  ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset    )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_60 userInterruptD_buffercc (
    .io_dataIn                      (userInterruptD                    ), //i
    .io_dataOut                     (userInterruptD_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                  ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset    )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_60 userInterruptC_buffercc (
    .io_dataIn                      (userInterruptC                    ), //i
    .io_dataOut                     (userInterruptC_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                  ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset    )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_60 userInterruptB_buffercc (
    .io_dataIn                      (userInterruptB                    ), //i
    .io_dataOut                     (userInterruptB_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                  ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset    )  //i
  );
  StreamFifo_15 dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo (
    .io_push_valid              (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_valid                    ), //i
    .io_push_ready              (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_push_ready       ), //o
    .io_push_payload            (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_payload[3:0]             ), //i
    .io_pop_valid               (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_valid        ), //o
    .io_pop_ready               (io_pop_rValidN                                                        ), //i
    .io_pop_payload             (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_payload[3:0] ), //o
    .io_flush                   (1'b0                                                                  ), //i
    .io_occupancy               (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_occupancy[5:0]   ), //o
    .io_availability            (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_availability[5:0]), //o
    .io_systemClk               (io_systemClk                                                          ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                                            )  //i
  );
  StreamFifo_15 dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1 (
    .io_push_valid              (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_valid_1                    ), //i
    .io_push_ready              (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_push_ready       ), //o
    .io_push_payload            (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_payload_1[3:0]             ), //i
    .io_pop_valid               (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_valid        ), //o
    .io_pop_ready               (io_pop_rValidN_1                                                        ), //i
    .io_pop_payload             (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_payload[3:0] ), //o
    .io_flush                   (1'b0                                                                    ), //i
    .io_occupancy               (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_occupancy[5:0]   ), //o
    .io_availability            (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_availability[5:0]), //o
    .io_systemClk               (io_systemClk                                                            ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                                              )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_60 system_coreStopTime_buffercc (
    .io_dataIn                      (system_coreStopTime                    ), //i
    .io_dataOut                     (system_coreStopTime_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                       ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset         )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_65 system_riscvJtag_debug_systemReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn                          (system_riscvJtag_debug_systemReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut                         (system_riscvJtag_debug_systemReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_memoryClk                       (io_memoryClk                                                                  ), //i
    .system_riscvJtag_debug_systemReset (system_riscvJtag_debug_systemReset                                            )  //i
  );
  DebugTransportModuleTunneled system_riscvJtag_hard_noTap_tunnel (
    .io_instruction_tdi         (jtagCtrl_tdi                                                      ), //i
    .io_instruction_enable      (jtagCtrl_enable                                                   ), //i
    .io_instruction_capture     (jtagCtrl_capture                                                  ), //i
    .io_instruction_shift       (jtagCtrl_shift                                                    ), //i
    .io_instruction_update      (jtagCtrl_update                                                   ), //i
    .io_instruction_reset       (jtagCtrl_reset                                                    ), //i
    .io_instruction_tdo         (system_riscvJtag_hard_noTap_tunnel_io_instruction_tdo             ), //o
    .io_bus_cmd_valid           (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_valid               ), //o
    .io_bus_cmd_ready           (system_riscvJtag_debug_logic_dm_io_ctrl_cmd_ready                 ), //i
    .io_bus_cmd_payload_write   (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_write       ), //o
    .io_bus_cmd_payload_data    (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_data[31:0]  ), //o
    .io_bus_cmd_payload_address (system_riscvJtag_hard_noTap_tunnel_io_bus_cmd_payload_address[6:0]), //o
    .io_bus_rsp_valid           (system_riscvJtag_debug_logic_dm_io_ctrl_rsp_valid                 ), //i
    .io_bus_rsp_payload_error   (system_riscvJtag_debug_logic_dm_io_ctrl_rsp_payload_error         ), //i
    .io_bus_rsp_payload_data    (system_riscvJtag_debug_logic_dm_io_ctrl_rsp_payload_data[31:0]    ), //i
    .jtagCtrl_tck               (jtagCtrl_tck                                                      ), //i
    .io_systemClk               (io_systemClk                                                      ), //i
    .debugCd_logic_outputReset  (debugCd_logic_outputReset                                         )  //i
  );
  BmbArbiter system_fabric_iBus_bmb_arbiter (
    .io_inputs_0_cmd_valid                    (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid                         ), //i
    .io_inputs_0_cmd_ready                    (system_fabric_iBus_bmb_arbiter_io_inputs_0_cmd_ready                                                  ), //o
    .io_inputs_0_cmd_payload_last             (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last                  ), //i
    .io_inputs_0_cmd_payload_fragment_opcode  (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode       ), //i
    .io_inputs_0_cmd_payload_fragment_address (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address[31:0]), //i
    .io_inputs_0_cmd_payload_fragment_length  (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length[5:0]  ), //i
    .io_inputs_0_rsp_valid                    (system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_valid                                                  ), //o
    .io_inputs_0_rsp_ready                    (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready                         ), //i
    .io_inputs_0_rsp_payload_last             (system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_last                                           ), //o
    .io_inputs_0_rsp_payload_fragment_opcode  (system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode                                ), //o
    .io_inputs_0_rsp_payload_fragment_data    (system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data[63:0]                            ), //o
    .io_inputs_1_cmd_valid                    (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_valid                         ), //i
    .io_inputs_1_cmd_ready                    (system_fabric_iBus_bmb_arbiter_io_inputs_1_cmd_ready                                                  ), //o
    .io_inputs_1_cmd_payload_last             (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_last                  ), //i
    .io_inputs_1_cmd_payload_fragment_opcode  (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_opcode       ), //i
    .io_inputs_1_cmd_payload_fragment_address (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_address[31:0]), //i
    .io_inputs_1_cmd_payload_fragment_length  (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_length[5:0]  ), //i
    .io_inputs_1_rsp_valid                    (system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_valid                                                  ), //o
    .io_inputs_1_rsp_ready                    (system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready                         ), //i
    .io_inputs_1_rsp_payload_last             (system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_last                                           ), //o
    .io_inputs_1_rsp_payload_fragment_opcode  (system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode                                ), //o
    .io_inputs_1_rsp_payload_fragment_data    (system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data[63:0]                            ), //o
    .io_output_cmd_valid                      (system_fabric_iBus_bmb_arbiter_io_output_cmd_valid                                                    ), //o
    .io_output_cmd_ready                      (system_fabric_iBus_bmb_cmd_ready                                                                      ), //i
    .io_output_cmd_payload_last               (system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_last                                             ), //o
    .io_output_cmd_payload_fragment_source    (system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_source                                  ), //o
    .io_output_cmd_payload_fragment_opcode    (system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_opcode                                  ), //o
    .io_output_cmd_payload_fragment_address   (system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_address[31:0]                           ), //o
    .io_output_cmd_payload_fragment_length    (system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_length[5:0]                             ), //o
    .io_output_rsp_valid                      (system_fabric_iBus_bmb_rsp_valid                                                                      ), //i
    .io_output_rsp_ready                      (system_fabric_iBus_bmb_arbiter_io_output_rsp_ready                                                    ), //o
    .io_output_rsp_payload_last               (system_fabric_iBus_bmb_rsp_payload_last                                                               ), //i
    .io_output_rsp_payload_fragment_source    (system_fabric_iBus_bmb_rsp_payload_fragment_source                                                    ), //i
    .io_output_rsp_payload_fragment_opcode    (system_fabric_iBus_bmb_rsp_payload_fragment_opcode                                                    ), //i
    .io_output_rsp_payload_fragment_data      (system_fabric_iBus_bmb_rsp_payload_fragment_data[63:0]                                                ), //i
    .io_systemClk                             (io_systemClk                                                                                          ), //i
    .systemCd_logic_outputReset               (systemCd_logic_outputReset                                                                            )  //i
  );
  BmbInvalidateMonitor system_fabric_invalidationMonitor_logic_monitor (
    .io_input_cmd_valid                     (system_fabric_invalidationMonitor_logic_input_cmd_valid                                     ), //i
    .io_input_cmd_ready                     (system_fabric_invalidationMonitor_logic_monitor_io_input_cmd_ready                          ), //o
    .io_input_cmd_payload_last              (system_fabric_invalidationMonitor_logic_input_cmd_payload_last                              ), //i
    .io_input_cmd_payload_fragment_source   (system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_source                   ), //i
    .io_input_cmd_payload_fragment_opcode   (system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_opcode                   ), //i
    .io_input_cmd_payload_fragment_address  (system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_address[31:0]            ), //i
    .io_input_cmd_payload_fragment_length   (system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_length[5:0]              ), //i
    .io_input_cmd_payload_fragment_data     (system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_data[63:0]               ), //i
    .io_input_cmd_payload_fragment_mask     (system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_mask[7:0]                ), //i
    .io_input_cmd_payload_fragment_context  (system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_context[4:0]             ), //i
    .io_input_rsp_valid                     (system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_valid                          ), //o
    .io_input_rsp_ready                     (system_fabric_invalidationMonitor_logic_input_rsp_ready                                     ), //i
    .io_input_rsp_payload_last              (system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_last                   ), //o
    .io_input_rsp_payload_fragment_source   (system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_source        ), //o
    .io_input_rsp_payload_fragment_opcode   (system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_opcode        ), //o
    .io_input_rsp_payload_fragment_data     (system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_data[63:0]    ), //o
    .io_input_rsp_payload_fragment_context  (system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_context[4:0]  ), //o
    .io_input_inv_valid                     (system_fabric_invalidationMonitor_logic_monitor_io_input_inv_valid                          ), //o
    .io_input_inv_ready                     (system_fabric_invalidationMonitor_logic_input_inv_ready                                     ), //i
    .io_input_inv_payload_all               (system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_all                    ), //o
    .io_input_inv_payload_address           (system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_address[31:0]          ), //o
    .io_input_inv_payload_length            (system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_length[5:0]            ), //o
    .io_input_inv_payload_source            (system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_source                 ), //o
    .io_input_ack_valid                     (system_fabric_invalidationMonitor_logic_input_ack_valid                                     ), //i
    .io_input_ack_ready                     (system_fabric_invalidationMonitor_logic_monitor_io_input_ack_ready                          ), //o
    .io_input_sync_valid                    (system_fabric_invalidationMonitor_logic_monitor_io_input_sync_valid                         ), //o
    .io_input_sync_ready                    (system_fabric_invalidationMonitor_logic_input_sync_ready                                    ), //i
    .io_input_sync_payload_source           (system_fabric_invalidationMonitor_logic_monitor_io_input_sync_payload_source                ), //o
    .io_output_cmd_valid                    (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_valid                         ), //o
    .io_output_cmd_ready                    (io_output_cmd_rValidN                                                                       ), //i
    .io_output_cmd_payload_last             (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_last                  ), //o
    .io_output_cmd_payload_fragment_source  (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_source       ), //o
    .io_output_cmd_payload_fragment_opcode  (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_opcode       ), //o
    .io_output_cmd_payload_fragment_address (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_address[31:0]), //o
    .io_output_cmd_payload_fragment_length  (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_length[5:0]  ), //o
    .io_output_cmd_payload_fragment_data    (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_data[63:0]   ), //o
    .io_output_cmd_payload_fragment_mask    (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_mask[7:0]    ), //o
    .io_output_cmd_payload_fragment_context (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_context[43:0]), //o
    .io_output_rsp_valid                    (_zz_when_Stream_l375                                                                        ), //i
    .io_output_rsp_ready                    (system_fabric_invalidationMonitor_logic_monitor_io_output_rsp_ready                         ), //o
    .io_output_rsp_payload_last             (_zz_io_output_rsp_payload_last                                                              ), //i
    .io_output_rsp_payload_fragment_source  (_zz_io_output_rsp_payload_fragment_source                                                   ), //i
    .io_output_rsp_payload_fragment_opcode  (_zz_io_output_rsp_payload_fragment_opcode                                                   ), //i
    .io_output_rsp_payload_fragment_data    (_zz_io_output_rsp_payload_fragment_data[63:0]                                               ), //i
    .io_output_rsp_payload_fragment_context (_zz_io_output_rsp_payload_fragment_context[43:0]                                            ), //i
    .io_systemClk                           (io_systemClk                                                                                ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                                                  )  //i
  );
  BmbExclusiveMonitor system_fabric_exclusiveMonitor_logic (
    .io_input_cmd_valid                      (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid                         ), //i
    .io_input_cmd_ready                      (system_fabric_exclusiveMonitor_logic_io_input_cmd_ready                                                                       ), //o
    .io_input_cmd_payload_last               (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last                  ), //i
    .io_input_cmd_payload_fragment_source    (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source       ), //i
    .io_input_cmd_payload_fragment_opcode    (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_exclusive (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_exclusive    ), //i
    .io_input_cmd_payload_fragment_address   (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address[31:0]), //i
    .io_input_cmd_payload_fragment_length    (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length[5:0]  ), //i
    .io_input_cmd_payload_fragment_data      (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data[63:0]   ), //i
    .io_input_cmd_payload_fragment_mask      (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask[7:0]    ), //i
    .io_input_cmd_payload_fragment_context   (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context[3:0] ), //i
    .io_input_rsp_valid                      (system_fabric_exclusiveMonitor_logic_io_input_rsp_valid                                                                       ), //o
    .io_input_rsp_ready                      (_zz_io_input_rsp_ready                                                                                                        ), //i
    .io_input_rsp_payload_last               (system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_last                                                                ), //o
    .io_input_rsp_payload_fragment_source    (system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_source                                                     ), //o
    .io_input_rsp_payload_fragment_opcode    (system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_opcode                                                     ), //o
    .io_input_rsp_payload_fragment_exclusive (system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_exclusive                                                  ), //o
    .io_input_rsp_payload_fragment_data      (system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_data[63:0]                                                 ), //o
    .io_input_rsp_payload_fragment_context   (system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_context[3:0]                                               ), //o
    .io_input_inv_valid                      (system_fabric_exclusiveMonitor_logic_io_input_inv_valid                                                                       ), //o
    .io_input_inv_ready                      (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_ready                                         ), //i
    .io_input_inv_payload_all                (system_fabric_exclusiveMonitor_logic_io_input_inv_payload_all                                                                 ), //o
    .io_input_inv_payload_address            (system_fabric_exclusiveMonitor_logic_io_input_inv_payload_address[31:0]                                                       ), //o
    .io_input_inv_payload_length             (system_fabric_exclusiveMonitor_logic_io_input_inv_payload_length[5:0]                                                         ), //o
    .io_input_inv_payload_source             (system_fabric_exclusiveMonitor_logic_io_input_inv_payload_source                                                              ), //o
    .io_input_ack_valid                      (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_combStage_valid                               ), //i
    .io_input_ack_ready                      (system_fabric_exclusiveMonitor_logic_io_input_ack_ready                                                                       ), //o
    .io_input_sync_valid                     (system_fabric_exclusiveMonitor_logic_io_input_sync_valid                                                                      ), //o
    .io_input_sync_ready                     (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_ready                                        ), //i
    .io_input_sync_payload_source            (system_fabric_exclusiveMonitor_logic_io_input_sync_payload_source                                                             ), //o
    .io_output_cmd_valid                     (system_fabric_exclusiveMonitor_logic_io_output_cmd_valid                                                                      ), //o
    .io_output_cmd_ready                     (system_fabric_exclusiveMonitor_output_connector_decoder_cmd_ready                                                             ), //i
    .io_output_cmd_payload_last              (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_last                                                               ), //o
    .io_output_cmd_payload_fragment_source   (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_source                                                    ), //o
    .io_output_cmd_payload_fragment_opcode   (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_opcode                                                    ), //o
    .io_output_cmd_payload_fragment_address  (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_address[31:0]                                             ), //o
    .io_output_cmd_payload_fragment_length   (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_length[5:0]                                               ), //o
    .io_output_cmd_payload_fragment_data     (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_data[63:0]                                                ), //o
    .io_output_cmd_payload_fragment_mask     (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_mask[7:0]                                                 ), //o
    .io_output_cmd_payload_fragment_context  (system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_context[4:0]                                              ), //o
    .io_output_rsp_valid                     (system_fabric_exclusiveMonitor_output_connector_decoder_rsp_valid                                                             ), //i
    .io_output_rsp_ready                     (system_fabric_exclusiveMonitor_logic_io_output_rsp_ready                                                                      ), //o
    .io_output_rsp_payload_last              (system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_last                                                      ), //i
    .io_output_rsp_payload_fragment_source   (system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_source                                           ), //i
    .io_output_rsp_payload_fragment_opcode   (system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_opcode                                           ), //i
    .io_output_rsp_payload_fragment_data     (system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_data[63:0]                                       ), //i
    .io_output_rsp_payload_fragment_context  (system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_context[4:0]                                     ), //i
    .io_output_inv_valid                     (system_fabric_exclusiveMonitor_output_connector_decoder_inv_valid                                                             ), //i
    .io_output_inv_ready                     (system_fabric_exclusiveMonitor_logic_io_output_inv_ready                                                                      ), //o
    .io_output_inv_payload_all               (system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_all                                                       ), //i
    .io_output_inv_payload_address           (system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_address[31:0]                                             ), //i
    .io_output_inv_payload_length            (system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_length[5:0]                                               ), //i
    .io_output_inv_payload_source            (system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_source                                                    ), //i
    .io_output_ack_valid                     (system_fabric_exclusiveMonitor_logic_io_output_ack_valid                                                                      ), //o
    .io_output_ack_ready                     (system_fabric_exclusiveMonitor_output_connector_decoder_ack_ready                                                             ), //i
    .io_output_sync_valid                    (system_fabric_exclusiveMonitor_output_connector_decoder_sync_valid                                                            ), //i
    .io_output_sync_ready                    (system_fabric_exclusiveMonitor_logic_io_output_sync_ready                                                                     ), //o
    .io_output_sync_payload_source           (system_fabric_exclusiveMonitor_output_connector_decoder_sync_payload_source                                                   ), //i
    .io_systemClk                            (io_systemClk                                                                                                                  ), //i
    .systemCd_logic_outputReset              (systemCd_logic_outputReset                                                                                                    )  //i
  );
  BmbArbiter_1 system_fabric_dBusCoherent_bmb_arbiter (
    .io_inputs_0_cmd_valid                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid                         ), //i
    .io_inputs_0_cmd_ready                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_cmd_ready                                                  ), //o
    .io_inputs_0_cmd_payload_last               (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last                  ), //i
    .io_inputs_0_cmd_payload_fragment_opcode    (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode       ), //i
    .io_inputs_0_cmd_payload_fragment_exclusive (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_exclusive    ), //i
    .io_inputs_0_cmd_payload_fragment_address   (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address[31:0]), //i
    .io_inputs_0_cmd_payload_fragment_length    (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length[5:0]  ), //i
    .io_inputs_0_cmd_payload_fragment_data      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_data[63:0]   ), //i
    .io_inputs_0_cmd_payload_fragment_mask      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_mask[7:0]    ), //i
    .io_inputs_0_cmd_payload_fragment_context   (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_context[3:0] ), //i
    .io_inputs_0_rsp_valid                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_valid                                                  ), //o
    .io_inputs_0_rsp_ready                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready                         ), //i
    .io_inputs_0_rsp_payload_last               (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_last                                           ), //o
    .io_inputs_0_rsp_payload_fragment_opcode    (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode                                ), //o
    .io_inputs_0_rsp_payload_fragment_exclusive (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_exclusive                             ), //o
    .io_inputs_0_rsp_payload_fragment_data      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data[63:0]                            ), //o
    .io_inputs_0_rsp_payload_fragment_context   (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_context[3:0]                          ), //o
    .io_inputs_0_inv_valid                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_valid                                                  ), //o
    .io_inputs_0_inv_ready                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready                         ), //i
    .io_inputs_0_inv_payload_all                (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_all                                            ), //o
    .io_inputs_0_inv_payload_address            (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_address[31:0]                                  ), //o
    .io_inputs_0_inv_payload_length             (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_length[5:0]                                    ), //o
    .io_inputs_0_ack_valid                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_ack_valid                         ), //i
    .io_inputs_0_ack_ready                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_ack_ready                                                  ), //o
    .io_inputs_0_sync_valid                     (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_sync_valid                                                 ), //o
    .io_inputs_0_sync_ready                     (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready                        ), //i
    .io_inputs_1_cmd_valid                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_valid                         ), //i
    .io_inputs_1_cmd_ready                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_cmd_ready                                                  ), //o
    .io_inputs_1_cmd_payload_last               (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_last                  ), //i
    .io_inputs_1_cmd_payload_fragment_opcode    (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_opcode       ), //i
    .io_inputs_1_cmd_payload_fragment_exclusive (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_exclusive    ), //i
    .io_inputs_1_cmd_payload_fragment_address   (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_address[31:0]), //i
    .io_inputs_1_cmd_payload_fragment_length    (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_length[5:0]  ), //i
    .io_inputs_1_cmd_payload_fragment_data      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_data[63:0]   ), //i
    .io_inputs_1_cmd_payload_fragment_mask      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_mask[7:0]    ), //i
    .io_inputs_1_cmd_payload_fragment_context   (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_context[3:0] ), //i
    .io_inputs_1_rsp_valid                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_valid                                                  ), //o
    .io_inputs_1_rsp_ready                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready                         ), //i
    .io_inputs_1_rsp_payload_last               (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_last                                           ), //o
    .io_inputs_1_rsp_payload_fragment_opcode    (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode                                ), //o
    .io_inputs_1_rsp_payload_fragment_exclusive (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_exclusive                             ), //o
    .io_inputs_1_rsp_payload_fragment_data      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data[63:0]                            ), //o
    .io_inputs_1_rsp_payload_fragment_context   (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_context[3:0]                          ), //o
    .io_inputs_1_inv_valid                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_valid                                                  ), //o
    .io_inputs_1_inv_ready                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready                         ), //i
    .io_inputs_1_inv_payload_all                (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_all                                            ), //o
    .io_inputs_1_inv_payload_address            (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_address[31:0]                                  ), //o
    .io_inputs_1_inv_payload_length             (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_length[5:0]                                    ), //o
    .io_inputs_1_ack_valid                      (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_ack_valid                         ), //i
    .io_inputs_1_ack_ready                      (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_ack_ready                                                  ), //o
    .io_inputs_1_sync_valid                     (system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_sync_valid                                                 ), //o
    .io_inputs_1_sync_ready                     (system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready                        ), //i
    .io_output_cmd_valid                        (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_valid                                                    ), //o
    .io_output_cmd_ready                        (system_fabric_dBusCoherent_bmb_cmd_ready                                                                      ), //i
    .io_output_cmd_payload_last                 (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_last                                             ), //o
    .io_output_cmd_payload_fragment_source      (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_source                                  ), //o
    .io_output_cmd_payload_fragment_opcode      (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_opcode                                  ), //o
    .io_output_cmd_payload_fragment_exclusive   (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_exclusive                               ), //o
    .io_output_cmd_payload_fragment_address     (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_address[31:0]                           ), //o
    .io_output_cmd_payload_fragment_length      (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_length[5:0]                             ), //o
    .io_output_cmd_payload_fragment_data        (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_data[63:0]                              ), //o
    .io_output_cmd_payload_fragment_mask        (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_mask[7:0]                               ), //o
    .io_output_cmd_payload_fragment_context     (system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_context[3:0]                            ), //o
    .io_output_rsp_valid                        (system_fabric_dBusCoherent_bmb_rsp_valid                                                                      ), //i
    .io_output_rsp_ready                        (system_fabric_dBusCoherent_bmb_arbiter_io_output_rsp_ready                                                    ), //o
    .io_output_rsp_payload_last                 (system_fabric_dBusCoherent_bmb_rsp_payload_last                                                               ), //i
    .io_output_rsp_payload_fragment_source      (system_fabric_dBusCoherent_bmb_rsp_payload_fragment_source                                                    ), //i
    .io_output_rsp_payload_fragment_opcode      (system_fabric_dBusCoherent_bmb_rsp_payload_fragment_opcode                                                    ), //i
    .io_output_rsp_payload_fragment_exclusive   (system_fabric_dBusCoherent_bmb_rsp_payload_fragment_exclusive                                                 ), //i
    .io_output_rsp_payload_fragment_data        (system_fabric_dBusCoherent_bmb_rsp_payload_fragment_data[63:0]                                                ), //i
    .io_output_rsp_payload_fragment_context     (system_fabric_dBusCoherent_bmb_rsp_payload_fragment_context[3:0]                                              ), //i
    .io_output_inv_valid                        (system_fabric_dBusCoherent_bmb_inv_valid                                                                      ), //i
    .io_output_inv_ready                        (system_fabric_dBusCoherent_bmb_arbiter_io_output_inv_ready                                                    ), //o
    .io_output_inv_payload_all                  (system_fabric_dBusCoherent_bmb_inv_payload_all                                                                ), //i
    .io_output_inv_payload_address              (system_fabric_dBusCoherent_bmb_inv_payload_address[31:0]                                                      ), //i
    .io_output_inv_payload_length               (system_fabric_dBusCoherent_bmb_inv_payload_length[5:0]                                                        ), //i
    .io_output_inv_payload_source               (system_fabric_dBusCoherent_bmb_inv_payload_source                                                             ), //i
    .io_output_ack_valid                        (system_fabric_dBusCoherent_bmb_arbiter_io_output_ack_valid                                                    ), //o
    .io_output_ack_ready                        (system_fabric_dBusCoherent_bmb_ack_ready                                                                      ), //i
    .io_output_sync_valid                       (system_fabric_dBusCoherent_bmb_sync_valid                                                                     ), //i
    .io_output_sync_ready                       (system_fabric_dBusCoherent_bmb_arbiter_io_output_sync_ready                                                   ), //o
    .io_output_sync_payload_source              (system_fabric_dBusCoherent_bmb_sync_payload_source                                                            ), //i
    .io_systemClk                               (io_systemClk                                                                                                  ), //i
    .systemCd_logic_outputReset                 (systemCd_logic_outputReset                                                                                    )  //i
  );
  BmbDecoder system_fabric_iBus_bmb_decoder (
    .io_input_cmd_valid                        (system_fabric_iBus_bmb_cmd_m2sPipe_valid                                      ), //i
    .io_input_cmd_ready                        (system_fabric_iBus_bmb_decoder_io_input_cmd_ready                             ), //o
    .io_input_cmd_payload_last                 (system_fabric_iBus_bmb_cmd_m2sPipe_payload_last                               ), //i
    .io_input_cmd_payload_fragment_source      (system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_source                    ), //i
    .io_input_cmd_payload_fragment_opcode      (system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_opcode                    ), //i
    .io_input_cmd_payload_fragment_address     (system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_address[31:0]             ), //i
    .io_input_cmd_payload_fragment_length      (system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_length[5:0]               ), //i
    .io_input_rsp_valid                        (system_fabric_iBus_bmb_decoder_io_input_rsp_valid                             ), //o
    .io_input_rsp_ready                        (system_fabric_iBus_bmb_rsp_ready                                              ), //i
    .io_input_rsp_payload_last                 (system_fabric_iBus_bmb_decoder_io_input_rsp_payload_last                      ), //o
    .io_input_rsp_payload_fragment_source      (system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_source           ), //o
    .io_input_rsp_payload_fragment_opcode      (system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_opcode           ), //o
    .io_input_rsp_payload_fragment_data        (system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_data[63:0]       ), //o
    .io_outputs_0_cmd_valid                    (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_valid                         ), //o
    .io_outputs_0_cmd_ready                    (system_bridge_bmb_arbiter_io_inputs_1_cmd_ready                               ), //i
    .io_outputs_0_cmd_payload_last             (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_last                  ), //o
    .io_outputs_0_cmd_payload_fragment_source  (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_source       ), //o
    .io_outputs_0_cmd_payload_fragment_opcode  (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode       ), //o
    .io_outputs_0_cmd_payload_fragment_address (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_address[31:0]), //o
    .io_outputs_0_cmd_payload_fragment_length  (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_length[5:0]  ), //o
    .io_outputs_0_rsp_valid                    (system_bridge_bmb_arbiter_io_inputs_1_rsp_valid                               ), //i
    .io_outputs_0_rsp_ready                    (system_fabric_iBus_bmb_decoder_io_outputs_0_rsp_ready                         ), //o
    .io_outputs_0_rsp_payload_last             (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_last                        ), //i
    .io_outputs_0_rsp_payload_fragment_source  (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_source             ), //i
    .io_outputs_0_rsp_payload_fragment_opcode  (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode             ), //i
    .io_outputs_0_rsp_payload_fragment_data    (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data[63:0]         )  //i
  );
  BmbArbiter_2 system_bridge_bmb_arbiter (
    .io_inputs_0_cmd_valid                    (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid                         ), //i
    .io_inputs_0_cmd_ready                    (system_bridge_bmb_arbiter_io_inputs_0_cmd_ready                                                  ), //o
    .io_inputs_0_cmd_payload_last             (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last                  ), //i
    .io_inputs_0_cmd_payload_fragment_source  (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_source       ), //i
    .io_inputs_0_cmd_payload_fragment_opcode  (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode       ), //i
    .io_inputs_0_cmd_payload_fragment_address (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address[31:0]), //i
    .io_inputs_0_cmd_payload_fragment_length  (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length[5:0]  ), //i
    .io_inputs_0_cmd_payload_fragment_data    (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_data[63:0]   ), //i
    .io_inputs_0_cmd_payload_fragment_mask    (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_mask[7:0]    ), //i
    .io_inputs_0_cmd_payload_fragment_context (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_context[43:0]), //i
    .io_inputs_0_rsp_valid                    (system_bridge_bmb_arbiter_io_inputs_0_rsp_valid                                                  ), //o
    .io_inputs_0_rsp_ready                    (system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready                         ), //i
    .io_inputs_0_rsp_payload_last             (system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_last                                           ), //o
    .io_inputs_0_rsp_payload_fragment_source  (system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_source                                ), //o
    .io_inputs_0_rsp_payload_fragment_opcode  (system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode                                ), //o
    .io_inputs_0_rsp_payload_fragment_data    (system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data[63:0]                            ), //o
    .io_inputs_0_rsp_payload_fragment_context (system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_context[43:0]                         ), //o
    .io_inputs_1_cmd_valid                    (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_valid                                            ), //i
    .io_inputs_1_cmd_ready                    (system_bridge_bmb_arbiter_io_inputs_1_cmd_ready                                                  ), //o
    .io_inputs_1_cmd_payload_last             (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_last                                     ), //i
    .io_inputs_1_cmd_payload_fragment_source  (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_source                          ), //i
    .io_inputs_1_cmd_payload_fragment_opcode  (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode                          ), //i
    .io_inputs_1_cmd_payload_fragment_address (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_address[31:0]                   ), //i
    .io_inputs_1_cmd_payload_fragment_length  (system_fabric_iBus_bmb_decoder_io_outputs_0_cmd_payload_fragment_length[5:0]                     ), //i
    .io_inputs_1_cmd_payload_fragment_data    (64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx                             ), //i
    .io_inputs_1_cmd_payload_fragment_mask    (8'bxxxxxxxx                                                                                      ), //i
    .io_inputs_1_rsp_valid                    (system_bridge_bmb_arbiter_io_inputs_1_rsp_valid                                                  ), //o
    .io_inputs_1_rsp_ready                    (system_fabric_iBus_bmb_decoder_io_outputs_0_rsp_ready                                            ), //i
    .io_inputs_1_rsp_payload_last             (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_last                                           ), //o
    .io_inputs_1_rsp_payload_fragment_source  (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_source                                ), //o
    .io_inputs_1_rsp_payload_fragment_opcode  (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode                                ), //o
    .io_inputs_1_rsp_payload_fragment_data    (system_bridge_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data[63:0]                            ), //o
    .io_output_cmd_valid                      (system_bridge_bmb_arbiter_io_output_cmd_valid                                                    ), //o
    .io_output_cmd_ready                      (system_bridge_bmb_cmd_ready                                                                      ), //i
    .io_output_cmd_payload_last               (system_bridge_bmb_arbiter_io_output_cmd_payload_last                                             ), //o
    .io_output_cmd_payload_fragment_source    (system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_source[1:0]                             ), //o
    .io_output_cmd_payload_fragment_opcode    (system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_opcode                                  ), //o
    .io_output_cmd_payload_fragment_address   (system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_address[31:0]                           ), //o
    .io_output_cmd_payload_fragment_length    (system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_length[5:0]                             ), //o
    .io_output_cmd_payload_fragment_data      (system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_data[63:0]                              ), //o
    .io_output_cmd_payload_fragment_mask      (system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_mask[7:0]                               ), //o
    .io_output_cmd_payload_fragment_context   (system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_context[43:0]                           ), //o
    .io_output_rsp_valid                      (system_bridge_bmb_rsp_valid                                                                      ), //i
    .io_output_rsp_ready                      (system_bridge_bmb_arbiter_io_output_rsp_ready                                                    ), //o
    .io_output_rsp_payload_last               (system_bridge_bmb_rsp_payload_last                                                               ), //i
    .io_output_rsp_payload_fragment_source    (system_bridge_bmb_rsp_payload_fragment_source[1:0]                                               ), //i
    .io_output_rsp_payload_fragment_opcode    (system_bridge_bmb_rsp_payload_fragment_opcode                                                    ), //i
    .io_output_rsp_payload_fragment_data      (system_bridge_bmb_rsp_payload_fragment_data[63:0]                                                ), //i
    .io_output_rsp_payload_fragment_context   (system_bridge_bmb_rsp_payload_fragment_context[43:0]                                             ), //i
    .io_systemClk                             (io_systemClk                                                                                     ), //i
    .systemCd_logic_outputReset               (systemCd_logic_outputReset                                                                       )  //i
  );
  BmbToAxi4SharedBridge system_ddr_ddrLogic_bmbToAxiBridge (
    .io_input_cmd_valid                    (io_output_cmd_m2sPipe_valid                                                   ), //i
    .io_input_cmd_ready                    (system_ddr_ddrLogic_bmbToAxiBridge_io_input_cmd_ready                         ), //o
    .io_input_cmd_payload_last             (io_output_cmd_m2sPipe_payload_last                                            ), //i
    .io_input_cmd_payload_fragment_source  (io_output_cmd_m2sPipe_payload_fragment_source[1:0]                            ), //i
    .io_input_cmd_payload_fragment_opcode  (io_output_cmd_m2sPipe_payload_fragment_opcode                                 ), //i
    .io_input_cmd_payload_fragment_address (io_output_cmd_m2sPipe_payload_fragment_address[31:0]                          ), //i
    .io_input_cmd_payload_fragment_length  (io_output_cmd_m2sPipe_payload_fragment_length[5:0]                            ), //i
    .io_input_cmd_payload_fragment_data    (io_output_cmd_m2sPipe_payload_fragment_data[127:0]                            ), //i
    .io_input_cmd_payload_fragment_mask    (io_output_cmd_m2sPipe_payload_fragment_mask[15:0]                             ), //i
    .io_input_cmd_payload_fragment_context (io_output_cmd_m2sPipe_payload_fragment_context[45:0]                          ), //i
    .io_input_rsp_valid                    (system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_valid                         ), //o
    .io_input_rsp_ready                    (_zz_io_input_rsp_ready_1                                                      ), //i
    .io_input_rsp_payload_last             (system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_last                  ), //o
    .io_input_rsp_payload_fragment_source  (system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_source[1:0]  ), //o
    .io_input_rsp_payload_fragment_opcode  (system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_opcode       ), //o
    .io_input_rsp_payload_fragment_data    (system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_data[127:0]  ), //o
    .io_input_rsp_payload_fragment_context (system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_context[45:0]), //o
    .io_output_arw_valid                   (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_valid                        ), //o
    .io_output_arw_ready                   (io_output_arw_rValidN                                                         ), //i
    .io_output_arw_payload_addr            (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_addr[31:0]           ), //o
    .io_output_arw_payload_len             (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_len[7:0]             ), //o
    .io_output_arw_payload_size            (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_size[2:0]            ), //o
    .io_output_arw_payload_cache           (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_cache[3:0]           ), //o
    .io_output_arw_payload_prot            (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_prot[2:0]            ), //o
    .io_output_arw_payload_write           (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_write                ), //o
    .io_output_w_valid                     (system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_valid                          ), //o
    .io_output_w_ready                     (io_output_w_rValidN                                                           ), //i
    .io_output_w_payload_data              (system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_data[127:0]            ), //o
    .io_output_w_payload_strb              (system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_strb[15:0]             ), //o
    .io_output_w_payload_last              (system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_last                   ), //o
    .io_output_b_valid                     (system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_valid                         ), //i
    .io_output_b_ready                     (system_ddr_ddrLogic_bmbToAxiBridge_io_output_b_ready                          ), //o
    .io_output_b_payload_resp              (system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_payload_resp[1:0]             ), //i
    .io_output_r_valid                     (system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_valid                         ), //i
    .io_output_r_ready                     (system_ddr_ddrLogic_bmbToAxiBridge_io_output_r_ready                          ), //o
    .io_output_r_payload_data              (system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_data[127:0]           ), //i
    .io_output_r_payload_resp              (system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_resp[1:0]             ), //i
    .io_output_r_payload_last              (system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_last                  ), //i
    .io_memoryClk                          (io_memoryClk                                                                  ), //i
    .ddrCd_logic_outputReset               (ddrCd_logic_outputReset                                                       )  //i
  );
  BmbCcFifo system_ddr_ddrLogic_cc_fifo (
    .io_input_cmd_valid                     (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid                         ), //i
    .io_input_cmd_ready                     (system_ddr_ddrLogic_cc_fifo_io_input_cmd_ready                                                          ), //o
    .io_input_cmd_payload_last              (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last                  ), //i
    .io_input_cmd_payload_fragment_source   (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source[1:0]  ), //i
    .io_input_cmd_payload_fragment_opcode   (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address  (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address[31:0]), //i
    .io_input_cmd_payload_fragment_length   (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length[5:0]  ), //i
    .io_input_cmd_payload_fragment_data     (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data[127:0]  ), //i
    .io_input_cmd_payload_fragment_mask     (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask[15:0]   ), //i
    .io_input_cmd_payload_fragment_context  (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context[45:0]), //i
    .io_input_rsp_valid                     (system_ddr_ddrLogic_cc_fifo_io_input_rsp_valid                                                          ), //o
    .io_input_rsp_ready                     (_zz_io_input_rsp_ready_2                                                                                ), //i
    .io_input_rsp_payload_last              (system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_last                                                   ), //o
    .io_input_rsp_payload_fragment_source   (system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_source[1:0]                                   ), //o
    .io_input_rsp_payload_fragment_opcode   (system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_opcode                                        ), //o
    .io_input_rsp_payload_fragment_data     (system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_data[127:0]                                   ), //o
    .io_input_rsp_payload_fragment_context  (system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_context[45:0]                                 ), //o
    .io_output_cmd_valid                    (system_ddr_ddrLogic_cc_fifo_io_output_cmd_valid                                                         ), //o
    .io_output_cmd_ready                    (system_ddr_ddrLogic_cc_fifo_io_output_cmd_ready                                                         ), //i
    .io_output_cmd_payload_last             (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_last                                                  ), //o
    .io_output_cmd_payload_fragment_source  (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_source[1:0]                                  ), //o
    .io_output_cmd_payload_fragment_opcode  (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_opcode                                       ), //o
    .io_output_cmd_payload_fragment_address (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_address[31:0]                                ), //o
    .io_output_cmd_payload_fragment_length  (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_length[5:0]                                  ), //o
    .io_output_cmd_payload_fragment_data    (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_data[127:0]                                  ), //o
    .io_output_cmd_payload_fragment_mask    (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_mask[15:0]                                   ), //o
    .io_output_cmd_payload_fragment_context (system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_context[45:0]                                ), //o
    .io_output_rsp_valid                    (_zz_when_Stream_l375_2                                                                                  ), //i
    .io_output_rsp_ready                    (system_ddr_ddrLogic_cc_fifo_io_output_rsp_ready                                                         ), //o
    .io_output_rsp_payload_last             (_zz_io_output_rsp_payload_last_1                                                                        ), //i
    .io_output_rsp_payload_fragment_source  (_zz_io_output_rsp_payload_fragment_source_1[1:0]                                                        ), //i
    .io_output_rsp_payload_fragment_opcode  (_zz_io_output_rsp_payload_fragment_opcode_1                                                             ), //i
    .io_output_rsp_payload_fragment_data    (_zz_io_output_rsp_payload_fragment_data_1[127:0]                                                        ), //i
    .io_output_rsp_payload_fragment_context (_zz_io_output_rsp_payload_fragment_context_1[45:0]                                                      ), //i
    .io_systemClk                           (io_systemClk                                                                                            ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                                                              ), //i
    .io_memoryClk                           (io_memoryClk                                                                                            ), //i
    .ddrCd_logic_outputReset                (ddrCd_logic_outputReset                                                                                 )  //i
  );
  Axi4ReadOnlyArbiter system_ddr_ddrLogic_arbiterAxi4Read (
    .io_inputs_0_ar_valid          (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_ar_valid              ), //i
    .io_inputs_0_ar_ready          (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_ar_ready              ), //o
    .io_inputs_0_ar_payload_addr   (system_ddr_ddrLogic_cpuAccess_arw_payload_addr[31:0]                  ), //i
    .io_inputs_0_ar_payload_id     (6'h0                                                                  ), //i
    .io_inputs_0_ar_payload_region (_zz_io_inputs_0_ar_payload_region[3:0]                                ), //i
    .io_inputs_0_ar_payload_len    (system_ddr_ddrLogic_cpuAccess_arw_payload_len[7:0]                    ), //i
    .io_inputs_0_ar_payload_size   (system_ddr_ddrLogic_cpuAccess_arw_payload_size[2:0]                   ), //i
    .io_inputs_0_ar_payload_burst  (2'b01                                                                 ), //i
    .io_inputs_0_ar_payload_lock   (1'b0                                                                  ), //i
    .io_inputs_0_ar_payload_cache  (system_ddr_ddrLogic_cpuAccess_arw_payload_cache[3:0]                  ), //i
    .io_inputs_0_ar_payload_qos    (4'b0000                                                               ), //i
    .io_inputs_0_ar_payload_prot   (system_ddr_ddrLogic_cpuAccess_arw_payload_prot[2:0]                   ), //i
    .io_inputs_0_r_valid           (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_valid               ), //o
    .io_inputs_0_r_ready           (system_ddr_ddrLogic_cpuAccess_r_ready                                 ), //i
    .io_inputs_0_r_payload_data    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_data[127:0] ), //o
    .io_inputs_0_r_payload_id      (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_id[5:0]     ), //o
    .io_inputs_0_r_payload_resp    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_resp[1:0]   ), //o
    .io_inputs_0_r_payload_last    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_last        ), //o
    .io_inputs_1_ar_valid          (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_valid              ), //i
    .io_inputs_1_ar_ready          (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_ar_ready              ), //o
    .io_inputs_1_ar_payload_addr   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_addr[31:0] ), //i
    .io_inputs_1_ar_payload_id     (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_ar_payload_id[5:0]    ), //i
    .io_inputs_1_ar_payload_region (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_region[3:0]), //i
    .io_inputs_1_ar_payload_len    (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_len[7:0]   ), //i
    .io_inputs_1_ar_payload_size   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_size[2:0]  ), //i
    .io_inputs_1_ar_payload_burst  (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_burst[1:0] ), //i
    .io_inputs_1_ar_payload_lock   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_lock       ), //i
    .io_inputs_1_ar_payload_cache  (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_cache[3:0] ), //i
    .io_inputs_1_ar_payload_qos    (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_qos[3:0]   ), //i
    .io_inputs_1_ar_payload_prot   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_prot[2:0]  ), //i
    .io_inputs_1_r_valid           (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_valid               ), //o
    .io_inputs_1_r_ready           (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_ready               ), //i
    .io_inputs_1_r_payload_data    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_data[127:0] ), //o
    .io_inputs_1_r_payload_id      (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_id[5:0]     ), //o
    .io_inputs_1_r_payload_resp    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_resp[1:0]   ), //o
    .io_inputs_1_r_payload_last    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_last        ), //o
    .io_inputs_2_ar_valid          (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_valid              ), //i
    .io_inputs_2_ar_ready          (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_ar_ready              ), //o
    .io_inputs_2_ar_payload_addr   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_addr[31:0] ), //i
    .io_inputs_2_ar_payload_id     (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_ar_payload_id[5:0]    ), //i
    .io_inputs_2_ar_payload_region (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_region[3:0]), //i
    .io_inputs_2_ar_payload_len    (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_len[7:0]   ), //i
    .io_inputs_2_ar_payload_size   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_size[2:0]  ), //i
    .io_inputs_2_ar_payload_burst  (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_burst[1:0] ), //i
    .io_inputs_2_ar_payload_lock   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_lock       ), //i
    .io_inputs_2_ar_payload_cache  (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_cache[3:0] ), //i
    .io_inputs_2_ar_payload_qos    (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_qos[3:0]   ), //i
    .io_inputs_2_ar_payload_prot   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_prot[2:0]  ), //i
    .io_inputs_2_r_valid           (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_valid               ), //o
    .io_inputs_2_r_ready           (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_ready               ), //i
    .io_inputs_2_r_payload_data    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_data[127:0] ), //o
    .io_inputs_2_r_payload_id      (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_id[5:0]     ), //o
    .io_inputs_2_r_payload_resp    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_resp[1:0]   ), //o
    .io_inputs_2_r_payload_last    (system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_last        ), //o
    .io_output_ar_valid            (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_valid                ), //o
    .io_output_ar_ready            (io_output_ar_rValidN                                                  ), //i
    .io_output_ar_payload_addr     (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_addr[31:0]   ), //o
    .io_output_ar_payload_id       (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_id[7:0]      ), //o
    .io_output_ar_payload_region   (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_region[3:0]  ), //o
    .io_output_ar_payload_len      (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_len[7:0]     ), //o
    .io_output_ar_payload_size     (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_size[2:0]    ), //o
    .io_output_ar_payload_burst    (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_burst[1:0]   ), //o
    .io_output_ar_payload_lock     (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_lock         ), //o
    .io_output_ar_payload_cache    (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_cache[3:0]   ), //o
    .io_output_ar_payload_qos      (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_qos[3:0]     ), //o
    .io_output_ar_payload_prot     (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_prot[2:0]    ), //o
    .io_output_r_valid             (system_ddr_ddrLogic_ddrAAxi4_r_valid                                  ), //i
    .io_output_r_ready             (system_ddr_ddrLogic_arbiterAxi4Read_io_output_r_ready                 ), //o
    .io_output_r_payload_data      (system_ddr_ddrLogic_ddrAAxi4_r_payload_data[127:0]                    ), //i
    .io_output_r_payload_id        (system_ddr_ddrLogic_ddrAAxi4_r_payload_id[7:0]                        ), //i
    .io_output_r_payload_resp      (system_ddr_ddrLogic_ddrAAxi4_r_payload_resp[1:0]                      ), //i
    .io_output_r_payload_last      (system_ddr_ddrLogic_ddrAAxi4_r_payload_last                           ), //i
    .io_memoryClk                  (io_memoryClk                                                          ), //i
    .ddrCd_logic_outputReset       (ddrCd_logic_outputReset                                               )  //i
  );
  Axi4WriteOnlyArbiter system_ddr_ddrLogic_arbiterAxi4Write (
    .io_inputs_0_aw_valid          (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_aw_valid             ), //i
    .io_inputs_0_aw_ready          (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_aw_ready             ), //o
    .io_inputs_0_aw_payload_addr   (system_ddr_ddrLogic_cpuAccess_arw_payload_addr[31:0]                  ), //i
    .io_inputs_0_aw_payload_id     (6'h0                                                                  ), //i
    .io_inputs_0_aw_payload_region (_zz_io_inputs_0_aw_payload_region[3:0]                                ), //i
    .io_inputs_0_aw_payload_len    (system_ddr_ddrLogic_cpuAccess_arw_payload_len[7:0]                    ), //i
    .io_inputs_0_aw_payload_size   (system_ddr_ddrLogic_cpuAccess_arw_payload_size[2:0]                   ), //i
    .io_inputs_0_aw_payload_burst  (2'b01                                                                 ), //i
    .io_inputs_0_aw_payload_lock   (1'b0                                                                  ), //i
    .io_inputs_0_aw_payload_cache  (system_ddr_ddrLogic_cpuAccess_arw_payload_cache[3:0]                  ), //i
    .io_inputs_0_aw_payload_qos    (4'b0000                                                               ), //i
    .io_inputs_0_aw_payload_prot   (system_ddr_ddrLogic_cpuAccess_arw_payload_prot[2:0]                   ), //i
    .io_inputs_0_w_valid           (system_ddr_ddrLogic_cpuAccess_w_valid                                 ), //i
    .io_inputs_0_w_ready           (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_w_ready              ), //o
    .io_inputs_0_w_payload_data    (system_ddr_ddrLogic_cpuAccess_w_payload_data[127:0]                   ), //i
    .io_inputs_0_w_payload_strb    (system_ddr_ddrLogic_cpuAccess_w_payload_strb[15:0]                    ), //i
    .io_inputs_0_w_payload_last    (system_ddr_ddrLogic_cpuAccess_w_payload_last                          ), //i
    .io_inputs_0_b_valid           (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_valid              ), //o
    .io_inputs_0_b_ready           (system_ddr_ddrLogic_cpuAccess_b_ready                                 ), //i
    .io_inputs_0_b_payload_id      (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_payload_id[5:0]    ), //o
    .io_inputs_0_b_payload_resp    (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_payload_resp[1:0]  ), //o
    .io_inputs_1_aw_valid          (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_valid              ), //i
    .io_inputs_1_aw_ready          (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_aw_ready             ), //o
    .io_inputs_1_aw_payload_addr   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_addr[31:0] ), //i
    .io_inputs_1_aw_payload_id     (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_aw_payload_id[5:0]   ), //i
    .io_inputs_1_aw_payload_region (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_region[3:0]), //i
    .io_inputs_1_aw_payload_len    (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_len[7:0]   ), //i
    .io_inputs_1_aw_payload_size   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_size[2:0]  ), //i
    .io_inputs_1_aw_payload_burst  (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_burst[1:0] ), //i
    .io_inputs_1_aw_payload_lock   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_lock       ), //i
    .io_inputs_1_aw_payload_cache  (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_cache[3:0] ), //i
    .io_inputs_1_aw_payload_qos    (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_qos[3:0]   ), //i
    .io_inputs_1_aw_payload_prot   (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_prot[2:0]  ), //i
    .io_inputs_1_w_valid           (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_valid               ), //i
    .io_inputs_1_w_ready           (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_w_ready              ), //o
    .io_inputs_1_w_payload_data    (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_data[127:0] ), //i
    .io_inputs_1_w_payload_strb    (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_strb[15:0]  ), //i
    .io_inputs_1_w_payload_last    (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_last        ), //i
    .io_inputs_1_b_valid           (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_valid              ), //o
    .io_inputs_1_b_ready           (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_ready               ), //i
    .io_inputs_1_b_payload_id      (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_payload_id[5:0]    ), //o
    .io_inputs_1_b_payload_resp    (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_payload_resp[1:0]  ), //o
    .io_inputs_2_aw_valid          (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_valid              ), //i
    .io_inputs_2_aw_ready          (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_aw_ready             ), //o
    .io_inputs_2_aw_payload_addr   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_addr[31:0] ), //i
    .io_inputs_2_aw_payload_id     (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_aw_payload_id[5:0]   ), //i
    .io_inputs_2_aw_payload_region (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_region[3:0]), //i
    .io_inputs_2_aw_payload_len    (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_len[7:0]   ), //i
    .io_inputs_2_aw_payload_size   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_size[2:0]  ), //i
    .io_inputs_2_aw_payload_burst  (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_burst[1:0] ), //i
    .io_inputs_2_aw_payload_lock   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_lock       ), //i
    .io_inputs_2_aw_payload_cache  (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_cache[3:0] ), //i
    .io_inputs_2_aw_payload_qos    (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_qos[3:0]   ), //i
    .io_inputs_2_aw_payload_prot   (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_prot[2:0]  ), //i
    .io_inputs_2_w_valid           (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_valid               ), //i
    .io_inputs_2_w_ready           (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_w_ready              ), //o
    .io_inputs_2_w_payload_data    (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_data[127:0] ), //i
    .io_inputs_2_w_payload_strb    (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_strb[15:0]  ), //i
    .io_inputs_2_w_payload_last    (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_last        ), //i
    .io_inputs_2_b_valid           (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_valid              ), //o
    .io_inputs_2_b_ready           (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_ready               ), //i
    .io_inputs_2_b_payload_id      (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_payload_id[5:0]    ), //o
    .io_inputs_2_b_payload_resp    (system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_payload_resp[1:0]  ), //o
    .io_output_aw_valid            (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_valid               ), //o
    .io_output_aw_ready            (io_output_aw_rValidN                                                  ), //i
    .io_output_aw_payload_addr     (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_addr[31:0]  ), //o
    .io_output_aw_payload_id       (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_id[7:0]     ), //o
    .io_output_aw_payload_region   (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_region[3:0] ), //o
    .io_output_aw_payload_len      (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_len[7:0]    ), //o
    .io_output_aw_payload_size     (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_size[2:0]   ), //o
    .io_output_aw_payload_burst    (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_burst[1:0]  ), //o
    .io_output_aw_payload_lock     (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_lock        ), //o
    .io_output_aw_payload_cache    (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_cache[3:0]  ), //o
    .io_output_aw_payload_qos      (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_qos[3:0]    ), //o
    .io_output_aw_payload_prot     (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_prot[2:0]   ), //o
    .io_output_w_valid             (system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_valid                ), //o
    .io_output_w_ready             (system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_ready                ), //i
    .io_output_w_payload_data      (system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_data[127:0]  ), //o
    .io_output_w_payload_strb      (system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_strb[15:0]   ), //o
    .io_output_w_payload_last      (system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_last         ), //o
    .io_output_b_valid             (system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_valid                  ), //i
    .io_output_b_ready             (system_ddr_ddrLogic_arbiterAxi4Write_io_output_b_ready                ), //o
    .io_output_b_payload_id        (system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_payload_id[7:0]        ), //i
    .io_output_b_payload_resp      (system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_payload_resp[1:0]      ), //i
    .io_memoryClk                  (io_memoryClk                                                          ), //i
    .ddrCd_logic_outputReset       (ddrCd_logic_outputReset                                               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_66 ddrCd_logic_outputReset_buffercc (
    .io_dataIn             (ddrCd_logic_outputReset                    ), //i
    .io_dataOut            (ddrCd_logic_outputReset_buffercc_io_dataOut), //o
    .io_ddrMasters_1_clk   (io_ddrMasters_1_clk                        ), //i
    .io_ddrMasters_1_reset (io_ddrMasters_1_reset_read_buffer          )  //i
  );
  Axi4CC system_ddr_ddrLogic_userAdapters_0_bridge (
    .io_input_aw_valid           (io_ddrMasters_1_aw_s2mPipe_m2sPipe_valid                                      ), //i
    .io_input_aw_ready           (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_aw_ready                   ), //o
    .io_input_aw_payload_addr    (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_addr[31:0]                         ), //i
    .io_input_aw_payload_id      (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_id[3:0]                            ), //i
    .io_input_aw_payload_region  (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_region[3:0]                        ), //i
    .io_input_aw_payload_len     (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_len[7:0]                           ), //i
    .io_input_aw_payload_size    (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_size[2:0]                          ), //i
    .io_input_aw_payload_burst   (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_burst[1:0]                         ), //i
    .io_input_aw_payload_lock    (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_lock                               ), //i
    .io_input_aw_payload_cache   (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_cache[3:0]                         ), //i
    .io_input_aw_payload_qos     (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_qos[3:0]                           ), //i
    .io_input_aw_payload_prot    (io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_prot[2:0]                          ), //i
    .io_input_w_valid            (io_ddrMasters_1_w_s2mPipe_m2sPipe_valid                                       ), //i
    .io_input_w_ready            (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_w_ready                    ), //o
    .io_input_w_payload_data     (io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_data[31:0]                          ), //i
    .io_input_w_payload_strb     (io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_strb[3:0]                           ), //i
    .io_input_w_payload_last     (io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_last                                ), //i
    .io_input_b_valid            (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_valid                    ), //o
    .io_input_b_ready            (io_input_b_rValidN                                                            ), //i
    .io_input_b_payload_id       (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_id[3:0]          ), //o
    .io_input_b_payload_resp     (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_resp[1:0]        ), //o
    .io_input_ar_valid           (io_ddrMasters_1_ar_halfPipe_valid                                             ), //i
    .io_input_ar_ready           (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_ar_ready                   ), //o
    .io_input_ar_payload_addr    (io_ddrMasters_1_ar_halfPipe_payload_addr[31:0]                                ), //i
    .io_input_ar_payload_id      (io_ddrMasters_1_ar_halfPipe_payload_id[3:0]                                   ), //i
    .io_input_ar_payload_region  (io_ddrMasters_1_ar_halfPipe_payload_region[3:0]                               ), //i
    .io_input_ar_payload_len     (io_ddrMasters_1_ar_halfPipe_payload_len[7:0]                                  ), //i
    .io_input_ar_payload_size    (io_ddrMasters_1_ar_halfPipe_payload_size[2:0]                                 ), //i
    .io_input_ar_payload_burst   (io_ddrMasters_1_ar_halfPipe_payload_burst[1:0]                                ), //i
    .io_input_ar_payload_lock    (io_ddrMasters_1_ar_halfPipe_payload_lock                                      ), //i
    .io_input_ar_payload_cache   (io_ddrMasters_1_ar_halfPipe_payload_cache[3:0]                                ), //i
    .io_input_ar_payload_qos     (io_ddrMasters_1_ar_halfPipe_payload_qos[3:0]                                  ), //i
    .io_input_ar_payload_prot    (io_ddrMasters_1_ar_halfPipe_payload_prot[2:0]                                 ), //i
    .io_input_r_valid            (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_valid                    ), //o
    .io_input_r_ready            (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_ready                    ), //i
    .io_input_r_payload_data     (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_data[31:0]       ), //o
    .io_input_r_payload_id       (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_id[3:0]          ), //o
    .io_input_r_payload_resp     (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_resp[1:0]        ), //o
    .io_input_r_payload_last     (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_last             ), //o
    .io_output_aw_valid          (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_valid                  ), //o
    .io_output_aw_ready          (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_aw_ready            ), //i
    .io_output_aw_payload_addr   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_addr[31:0]     ), //o
    .io_output_aw_payload_id     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_id[3:0]        ), //o
    .io_output_aw_payload_region (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_region[3:0]    ), //o
    .io_output_aw_payload_len    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_len[7:0]       ), //o
    .io_output_aw_payload_size   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_size[2:0]      ), //o
    .io_output_aw_payload_burst  (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_burst[1:0]     ), //o
    .io_output_aw_payload_lock   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_lock           ), //o
    .io_output_aw_payload_cache  (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_cache[3:0]     ), //o
    .io_output_aw_payload_qos    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_qos[3:0]       ), //o
    .io_output_aw_payload_prot   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_prot[2:0]      ), //o
    .io_output_w_valid           (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_valid                   ), //o
    .io_output_w_ready           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_w_ready             ), //i
    .io_output_w_payload_data    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_data[31:0]      ), //o
    .io_output_w_payload_strb    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_strb[3:0]       ), //o
    .io_output_w_payload_last    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_last            ), //o
    .io_output_b_valid           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_valid             ), //i
    .io_output_b_ready           (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_b_ready                   ), //o
    .io_output_b_payload_id      (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_payload_id[3:0]   ), //i
    .io_output_b_payload_resp    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_payload_resp[1:0] ), //i
    .io_output_ar_valid          (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_valid                  ), //o
    .io_output_ar_ready          (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_ar_ready            ), //i
    .io_output_ar_payload_addr   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_addr[31:0]     ), //o
    .io_output_ar_payload_id     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_id[3:0]        ), //o
    .io_output_ar_payload_region (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_region[3:0]    ), //o
    .io_output_ar_payload_len    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_len[7:0]       ), //o
    .io_output_ar_payload_size   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_size[2:0]      ), //o
    .io_output_ar_payload_burst  (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_burst[1:0]     ), //o
    .io_output_ar_payload_lock   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_lock           ), //o
    .io_output_ar_payload_cache  (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_cache[3:0]     ), //o
    .io_output_ar_payload_qos    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_qos[3:0]       ), //o
    .io_output_ar_payload_prot   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_prot[2:0]      ), //o
    .io_output_r_valid           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_valid             ), //i
    .io_output_r_ready           (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_r_ready                   ), //o
    .io_output_r_payload_data    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_data[31:0]), //i
    .io_output_r_payload_id      (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_id[3:0]   ), //i
    .io_output_r_payload_resp    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_resp[1:0] ), //i
    .io_output_r_payload_last    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_last      ), //i
    .io_ddrMasters_1_clk         (io_ddrMasters_1_clk                                                           ), //i
    .io_ddrMasters_1_reset       (io_ddrMasters_1_reset_read_buffer                                             ), //i
    .io_memoryClk                (io_memoryClk                                                                  ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                                                       )  //i
  );
  Axi4Upsizer system_ddr_ddrLogic_userAdapters_0_upsizer_logic (
    .io_input_aw_valid           (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_valid                     ), //i
    .io_input_aw_ready           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_aw_ready               ), //o
    .io_input_aw_payload_addr    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_addr[31:0]        ), //i
    .io_input_aw_payload_id      (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_id[3:0]           ), //i
    .io_input_aw_payload_region  (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_region[3:0]       ), //i
    .io_input_aw_payload_len     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_len[7:0]          ), //i
    .io_input_aw_payload_size    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_size[2:0]         ), //i
    .io_input_aw_payload_burst   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_burst[1:0]        ), //i
    .io_input_aw_payload_lock    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_lock              ), //i
    .io_input_aw_payload_cache   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_cache[3:0]        ), //i
    .io_input_aw_payload_qos     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_qos[3:0]          ), //i
    .io_input_aw_payload_prot    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_aw_payload_prot[2:0]         ), //i
    .io_input_w_valid            (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_valid                      ), //i
    .io_input_w_ready            (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_w_ready                ), //o
    .io_input_w_payload_data     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_data[31:0]         ), //i
    .io_input_w_payload_strb     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_strb[3:0]          ), //i
    .io_input_w_payload_last     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_w_payload_last               ), //i
    .io_input_b_valid            (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_valid                ), //o
    .io_input_b_ready            (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_b_ready                      ), //i
    .io_input_b_payload_id       (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_payload_id[3:0]      ), //o
    .io_input_b_payload_resp     (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_b_payload_resp[1:0]    ), //o
    .io_input_ar_valid           (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_valid                     ), //i
    .io_input_ar_ready           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_ar_ready               ), //o
    .io_input_ar_payload_addr    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_addr[31:0]        ), //i
    .io_input_ar_payload_id      (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_id[3:0]           ), //i
    .io_input_ar_payload_region  (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_region[3:0]       ), //i
    .io_input_ar_payload_len     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_len[7:0]          ), //i
    .io_input_ar_payload_size    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_size[2:0]         ), //i
    .io_input_ar_payload_burst   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_burst[1:0]        ), //i
    .io_input_ar_payload_lock    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_lock              ), //i
    .io_input_ar_payload_cache   (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_cache[3:0]        ), //i
    .io_input_ar_payload_qos     (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_qos[3:0]          ), //i
    .io_input_ar_payload_prot    (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_ar_payload_prot[2:0]         ), //i
    .io_input_r_valid            (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_valid                ), //o
    .io_input_r_ready            (system_ddr_ddrLogic_userAdapters_0_bridge_io_output_r_ready                      ), //i
    .io_input_r_payload_data     (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_data[31:0]   ), //o
    .io_input_r_payload_id       (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_id[3:0]      ), //o
    .io_input_r_payload_resp     (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_resp[1:0]    ), //o
    .io_input_r_payload_last     (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_input_r_payload_last         ), //o
    .io_output_aw_valid          (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_valid              ), //o
    .io_output_aw_ready          (system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_ready                             ), //i
    .io_output_aw_payload_addr   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_addr[31:0] ), //o
    .io_output_aw_payload_id     (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_id[3:0]    ), //o
    .io_output_aw_payload_region (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_region[3:0]), //o
    .io_output_aw_payload_len    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_len[7:0]   ), //o
    .io_output_aw_payload_size   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_size[2:0]  ), //o
    .io_output_aw_payload_burst  (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_burst[1:0] ), //o
    .io_output_aw_payload_lock   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_lock       ), //o
    .io_output_aw_payload_cache  (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_cache[3:0] ), //o
    .io_output_aw_payload_qos    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_qos[3:0]   ), //o
    .io_output_aw_payload_prot   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_prot[2:0]  ), //o
    .io_output_w_valid           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_valid               ), //o
    .io_output_w_ready           (system_ddr_ddrLogic_userAdapters_0_userAxi4_w_ready                              ), //i
    .io_output_w_payload_data    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_data[127:0] ), //o
    .io_output_w_payload_strb    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_strb[15:0]  ), //o
    .io_output_w_payload_last    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_last        ), //o
    .io_output_b_valid           (system_ddr_ddrLogic_userAdapters_0_userAxi4_b_valid                              ), //i
    .io_output_b_ready           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_b_ready               ), //o
    .io_output_b_payload_id      (system_ddr_ddrLogic_userAdapters_0_userAxi4_b_payload_id[3:0]                    ), //i
    .io_output_b_payload_resp    (system_ddr_ddrLogic_userAdapters_0_userAxi4_b_payload_resp[1:0]                  ), //i
    .io_output_ar_valid          (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_valid              ), //o
    .io_output_ar_ready          (system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_ready                             ), //i
    .io_output_ar_payload_addr   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_addr[31:0] ), //o
    .io_output_ar_payload_id     (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_id[3:0]    ), //o
    .io_output_ar_payload_region (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_region[3:0]), //o
    .io_output_ar_payload_len    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_len[7:0]   ), //o
    .io_output_ar_payload_size   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_size[2:0]  ), //o
    .io_output_ar_payload_burst  (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_burst[1:0] ), //o
    .io_output_ar_payload_lock   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_lock       ), //o
    .io_output_ar_payload_cache  (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_cache[3:0] ), //o
    .io_output_ar_payload_qos    (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_qos[3:0]   ), //o
    .io_output_ar_payload_prot   (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_prot[2:0]  ), //o
    .io_output_r_valid           (system_ddr_ddrLogic_userAdapters_0_userAxi4_r_valid                              ), //i
    .io_output_r_ready           (system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_r_ready               ), //o
    .io_output_r_payload_data    (system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_data[127:0]                ), //i
    .io_output_r_payload_id      (system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_id[3:0]                    ), //i
    .io_output_r_payload_resp    (system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_resp[1:0]                  ), //i
    .io_output_r_payload_last    (system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_last                       ), //i
    .io_memoryClk                (io_memoryClk                                                                     ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                                                          )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_67 ddrCd_logic_outputReset_buffercc_1 (
    .io_dataIn             (ddrCd_logic_outputReset                      ), //i
    .io_dataOut            (ddrCd_logic_outputReset_buffercc_1_io_dataOut), //o
    .io_ddrMasters_0_clk   (io_ddrMasters_0_clk                          ), //i
    .io_ddrMasters_0_reset (io_ddrMasters_0_reset_read_buffer            )  //i
  );
  Axi4CC_1 system_ddr_ddrLogic_userAdapters_1_bridge (
    .io_input_aw_valid           (io_ddrMasters_0_aw_s2mPipe_m2sPipe_valid                                      ), //i
    .io_input_aw_ready           (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_aw_ready                   ), //o
    .io_input_aw_payload_addr    (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_addr[31:0]                         ), //i
    .io_input_aw_payload_id      (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_id[3:0]                            ), //i
    .io_input_aw_payload_region  (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_region[3:0]                        ), //i
    .io_input_aw_payload_len     (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_len[7:0]                           ), //i
    .io_input_aw_payload_size    (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_size[2:0]                          ), //i
    .io_input_aw_payload_burst   (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_burst[1:0]                         ), //i
    .io_input_aw_payload_lock    (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_lock                               ), //i
    .io_input_aw_payload_cache   (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_cache[3:0]                         ), //i
    .io_input_aw_payload_qos     (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_qos[3:0]                           ), //i
    .io_input_aw_payload_prot    (io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_prot[2:0]                          ), //i
    .io_input_w_valid            (io_ddrMasters_0_w_s2mPipe_m2sPipe_valid                                       ), //i
    .io_input_w_ready            (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_w_ready                    ), //o
    .io_input_w_payload_data     (io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_data[63:0]                          ), //i
    .io_input_w_payload_strb     (io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_strb[7:0]                           ), //i
    .io_input_w_payload_last     (io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_last                                ), //i
    .io_input_b_valid            (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_valid                    ), //o
    .io_input_b_ready            (io_input_b_rValidN_1                                                          ), //i
    .io_input_b_payload_id       (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_id[3:0]          ), //o
    .io_input_b_payload_resp     (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_resp[1:0]        ), //o
    .io_input_ar_valid           (io_ddrMasters_0_ar_halfPipe_valid                                             ), //i
    .io_input_ar_ready           (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_ar_ready                   ), //o
    .io_input_ar_payload_addr    (io_ddrMasters_0_ar_halfPipe_payload_addr[31:0]                                ), //i
    .io_input_ar_payload_id      (io_ddrMasters_0_ar_halfPipe_payload_id[3:0]                                   ), //i
    .io_input_ar_payload_region  (io_ddrMasters_0_ar_halfPipe_payload_region[3:0]                               ), //i
    .io_input_ar_payload_len     (io_ddrMasters_0_ar_halfPipe_payload_len[7:0]                                  ), //i
    .io_input_ar_payload_size    (io_ddrMasters_0_ar_halfPipe_payload_size[2:0]                                 ), //i
    .io_input_ar_payload_burst   (io_ddrMasters_0_ar_halfPipe_payload_burst[1:0]                                ), //i
    .io_input_ar_payload_lock    (io_ddrMasters_0_ar_halfPipe_payload_lock                                      ), //i
    .io_input_ar_payload_cache   (io_ddrMasters_0_ar_halfPipe_payload_cache[3:0]                                ), //i
    .io_input_ar_payload_qos     (io_ddrMasters_0_ar_halfPipe_payload_qos[3:0]                                  ), //i
    .io_input_ar_payload_prot    (io_ddrMasters_0_ar_halfPipe_payload_prot[2:0]                                 ), //i
    .io_input_r_valid            (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_valid                    ), //o
    .io_input_r_ready            (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_ready                    ), //i
    .io_input_r_payload_data     (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_data[63:0]       ), //o
    .io_input_r_payload_id       (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_id[3:0]          ), //o
    .io_input_r_payload_resp     (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_resp[1:0]        ), //o
    .io_input_r_payload_last     (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_last             ), //o
    .io_output_aw_valid          (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_valid                  ), //o
    .io_output_aw_ready          (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_aw_ready            ), //i
    .io_output_aw_payload_addr   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_addr[31:0]     ), //o
    .io_output_aw_payload_id     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_id[3:0]        ), //o
    .io_output_aw_payload_region (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_region[3:0]    ), //o
    .io_output_aw_payload_len    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_len[7:0]       ), //o
    .io_output_aw_payload_size   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_size[2:0]      ), //o
    .io_output_aw_payload_burst  (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_burst[1:0]     ), //o
    .io_output_aw_payload_lock   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_lock           ), //o
    .io_output_aw_payload_cache  (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_cache[3:0]     ), //o
    .io_output_aw_payload_qos    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_qos[3:0]       ), //o
    .io_output_aw_payload_prot   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_prot[2:0]      ), //o
    .io_output_w_valid           (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_valid                   ), //o
    .io_output_w_ready           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_w_ready             ), //i
    .io_output_w_payload_data    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_data[63:0]      ), //o
    .io_output_w_payload_strb    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_strb[7:0]       ), //o
    .io_output_w_payload_last    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_last            ), //o
    .io_output_b_valid           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_valid             ), //i
    .io_output_b_ready           (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_b_ready                   ), //o
    .io_output_b_payload_id      (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_payload_id[3:0]   ), //i
    .io_output_b_payload_resp    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_payload_resp[1:0] ), //i
    .io_output_ar_valid          (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_valid                  ), //o
    .io_output_ar_ready          (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_ar_ready            ), //i
    .io_output_ar_payload_addr   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_addr[31:0]     ), //o
    .io_output_ar_payload_id     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_id[3:0]        ), //o
    .io_output_ar_payload_region (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_region[3:0]    ), //o
    .io_output_ar_payload_len    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_len[7:0]       ), //o
    .io_output_ar_payload_size   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_size[2:0]      ), //o
    .io_output_ar_payload_burst  (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_burst[1:0]     ), //o
    .io_output_ar_payload_lock   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_lock           ), //o
    .io_output_ar_payload_cache  (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_cache[3:0]     ), //o
    .io_output_ar_payload_qos    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_qos[3:0]       ), //o
    .io_output_ar_payload_prot   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_prot[2:0]      ), //o
    .io_output_r_valid           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_valid             ), //i
    .io_output_r_ready           (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_r_ready                   ), //o
    .io_output_r_payload_data    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_data[63:0]), //i
    .io_output_r_payload_id      (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_id[3:0]   ), //i
    .io_output_r_payload_resp    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_resp[1:0] ), //i
    .io_output_r_payload_last    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_last      ), //i
    .io_ddrMasters_0_clk         (io_ddrMasters_0_clk                                                           ), //i
    .io_ddrMasters_0_reset       (io_ddrMasters_0_reset_read_buffer                                             ), //i
    .io_memoryClk                (io_memoryClk                                                                  ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                                                       )  //i
  );
  Axi4Upsizer_1 system_ddr_ddrLogic_userAdapters_1_upsizer_logic (
    .io_input_aw_valid           (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_valid                     ), //i
    .io_input_aw_ready           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_aw_ready               ), //o
    .io_input_aw_payload_addr    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_addr[31:0]        ), //i
    .io_input_aw_payload_id      (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_id[3:0]           ), //i
    .io_input_aw_payload_region  (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_region[3:0]       ), //i
    .io_input_aw_payload_len     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_len[7:0]          ), //i
    .io_input_aw_payload_size    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_size[2:0]         ), //i
    .io_input_aw_payload_burst   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_burst[1:0]        ), //i
    .io_input_aw_payload_lock    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_lock              ), //i
    .io_input_aw_payload_cache   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_cache[3:0]        ), //i
    .io_input_aw_payload_qos     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_qos[3:0]          ), //i
    .io_input_aw_payload_prot    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_aw_payload_prot[2:0]         ), //i
    .io_input_w_valid            (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_valid                      ), //i
    .io_input_w_ready            (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_w_ready                ), //o
    .io_input_w_payload_data     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_data[63:0]         ), //i
    .io_input_w_payload_strb     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_strb[7:0]          ), //i
    .io_input_w_payload_last     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_w_payload_last               ), //i
    .io_input_b_valid            (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_valid                ), //o
    .io_input_b_ready            (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_b_ready                      ), //i
    .io_input_b_payload_id       (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_payload_id[3:0]      ), //o
    .io_input_b_payload_resp     (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_b_payload_resp[1:0]    ), //o
    .io_input_ar_valid           (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_valid                     ), //i
    .io_input_ar_ready           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_ar_ready               ), //o
    .io_input_ar_payload_addr    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_addr[31:0]        ), //i
    .io_input_ar_payload_id      (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_id[3:0]           ), //i
    .io_input_ar_payload_region  (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_region[3:0]       ), //i
    .io_input_ar_payload_len     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_len[7:0]          ), //i
    .io_input_ar_payload_size    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_size[2:0]         ), //i
    .io_input_ar_payload_burst   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_burst[1:0]        ), //i
    .io_input_ar_payload_lock    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_lock              ), //i
    .io_input_ar_payload_cache   (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_cache[3:0]        ), //i
    .io_input_ar_payload_qos     (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_qos[3:0]          ), //i
    .io_input_ar_payload_prot    (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_ar_payload_prot[2:0]         ), //i
    .io_input_r_valid            (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_valid                ), //o
    .io_input_r_ready            (system_ddr_ddrLogic_userAdapters_1_bridge_io_output_r_ready                      ), //i
    .io_input_r_payload_data     (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_data[63:0]   ), //o
    .io_input_r_payload_id       (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_id[3:0]      ), //o
    .io_input_r_payload_resp     (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_resp[1:0]    ), //o
    .io_input_r_payload_last     (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_input_r_payload_last         ), //o
    .io_output_aw_valid          (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_valid              ), //o
    .io_output_aw_ready          (system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_ready                             ), //i
    .io_output_aw_payload_addr   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_addr[31:0] ), //o
    .io_output_aw_payload_id     (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_id[3:0]    ), //o
    .io_output_aw_payload_region (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_region[3:0]), //o
    .io_output_aw_payload_len    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_len[7:0]   ), //o
    .io_output_aw_payload_size   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_size[2:0]  ), //o
    .io_output_aw_payload_burst  (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_burst[1:0] ), //o
    .io_output_aw_payload_lock   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_lock       ), //o
    .io_output_aw_payload_cache  (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_cache[3:0] ), //o
    .io_output_aw_payload_qos    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_qos[3:0]   ), //o
    .io_output_aw_payload_prot   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_prot[2:0]  ), //o
    .io_output_w_valid           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_valid               ), //o
    .io_output_w_ready           (system_ddr_ddrLogic_userAdapters_1_userAxi4_w_ready                              ), //i
    .io_output_w_payload_data    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_data[127:0] ), //o
    .io_output_w_payload_strb    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_strb[15:0]  ), //o
    .io_output_w_payload_last    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_last        ), //o
    .io_output_b_valid           (system_ddr_ddrLogic_userAdapters_1_userAxi4_b_valid                              ), //i
    .io_output_b_ready           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_b_ready               ), //o
    .io_output_b_payload_id      (system_ddr_ddrLogic_userAdapters_1_userAxi4_b_payload_id[3:0]                    ), //i
    .io_output_b_payload_resp    (system_ddr_ddrLogic_userAdapters_1_userAxi4_b_payload_resp[1:0]                  ), //i
    .io_output_ar_valid          (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_valid              ), //o
    .io_output_ar_ready          (system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_ready                             ), //i
    .io_output_ar_payload_addr   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_addr[31:0] ), //o
    .io_output_ar_payload_id     (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_id[3:0]    ), //o
    .io_output_ar_payload_region (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_region[3:0]), //o
    .io_output_ar_payload_len    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_len[7:0]   ), //o
    .io_output_ar_payload_size   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_size[2:0]  ), //o
    .io_output_ar_payload_burst  (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_burst[1:0] ), //o
    .io_output_ar_payload_lock   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_lock       ), //o
    .io_output_ar_payload_cache  (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_cache[3:0] ), //o
    .io_output_ar_payload_qos    (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_qos[3:0]   ), //o
    .io_output_ar_payload_prot   (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_prot[2:0]  ), //o
    .io_output_r_valid           (system_ddr_ddrLogic_userAdapters_1_userAxi4_r_valid                              ), //i
    .io_output_r_ready           (system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_r_ready               ), //o
    .io_output_r_payload_data    (system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_data[127:0]                ), //i
    .io_output_r_payload_id      (system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_id[3:0]                    ), //i
    .io_output_r_payload_resp    (system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_resp[1:0]                  ), //i
    .io_output_r_payload_last    (system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_last                       ), //i
    .io_memoryClk                (io_memoryClk                                                                     ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                                                          )  //i
  );
  StreamFifoLowLatency_1 system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo (
    .io_push_valid                       (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_valid                       ), //i
    .io_push_ready                       (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_push_ready          ), //o
    .io_push_payload_len                 (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_payload_len[7:0]            ), //i
    .io_pop_valid                        (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_valid           ), //o
    .io_pop_ready                        (io_pop_rValidN_2                                                              ), //i
    .io_pop_payload_len                  (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_payload_len[7:0]), //o
    .io_flush                            (1'b0                                                                          ), //i
    .io_occupancy                        (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_occupancy[2:0]      ), //o
    .io_availability                     (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_availability[2:0]   ), //o
    .io_memoryClk                        (io_memoryClk                                                                  ), //i
    .system_ddr_ddrLogic_ddrAReset_reset (system_ddr_ddrLogic_ddrAReset_reset                                           )  //i
  );
  BmbToAxi4SharedBridge_1 system_axiA_logic_bmbToAxiBridge (
    .io_input_cmd_valid                    (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid                         ), //i
    .io_input_cmd_ready                    (system_axiA_logic_bmbToAxiBridge_io_input_cmd_ready                                                      ), //o
    .io_input_cmd_payload_last             (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last                  ), //i
    .io_input_cmd_payload_fragment_source  (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source[1:0]  ), //i
    .io_input_cmd_payload_fragment_opcode  (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address[31:0]), //i
    .io_input_cmd_payload_fragment_length  (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length[5:0]  ), //i
    .io_input_cmd_payload_fragment_data    (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data[31:0]   ), //i
    .io_input_cmd_payload_fragment_mask    (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask[3:0]    ), //i
    .io_input_cmd_payload_fragment_context (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context[44:0]), //i
    .io_input_rsp_valid                    (system_axiA_logic_bmbToAxiBridge_io_input_rsp_valid                                                      ), //o
    .io_input_rsp_ready                    (_zz_io_input_rsp_ready_3                                                                                 ), //i
    .io_input_rsp_payload_last             (system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_last                                               ), //o
    .io_input_rsp_payload_fragment_source  (system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_source[1:0]                               ), //o
    .io_input_rsp_payload_fragment_opcode  (system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_opcode                                    ), //o
    .io_input_rsp_payload_fragment_data    (system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_data[31:0]                                ), //o
    .io_input_rsp_payload_fragment_context (system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_context[44:0]                             ), //o
    .io_output_arw_valid                   (system_axiA_logic_bmbToAxiBridge_io_output_arw_valid                                                     ), //o
    .io_output_arw_ready                   (system_axiA_logic_bmbToAxiBridge_io_output_arw_ready                                                     ), //i
    .io_output_arw_payload_addr            (system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_addr[31:0]                                        ), //o
    .io_output_arw_payload_len             (system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_len[7:0]                                          ), //o
    .io_output_arw_payload_size            (system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_size[2:0]                                         ), //o
    .io_output_arw_payload_cache           (system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_cache[3:0]                                        ), //o
    .io_output_arw_payload_prot            (system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_prot[2:0]                                         ), //o
    .io_output_arw_payload_write           (system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_write                                             ), //o
    .io_output_w_valid                     (system_axiA_logic_bmbToAxiBridge_io_output_w_valid                                                       ), //o
    .io_output_w_ready                     (system_axiA_logic_axiAAdapted_w_ready                                                                    ), //i
    .io_output_w_payload_data              (system_axiA_logic_bmbToAxiBridge_io_output_w_payload_data[31:0]                                          ), //o
    .io_output_w_payload_strb              (system_axiA_logic_bmbToAxiBridge_io_output_w_payload_strb[3:0]                                           ), //o
    .io_output_w_payload_last              (system_axiA_logic_bmbToAxiBridge_io_output_w_payload_last                                                ), //o
    .io_output_b_valid                     (system_axiA_logic_axiAAdapted_b_valid                                                                    ), //i
    .io_output_b_ready                     (system_axiA_logic_bmbToAxiBridge_io_output_b_ready                                                       ), //o
    .io_output_b_payload_resp              (system_axiA_logic_axiAAdapted_b_payload_resp[1:0]                                                        ), //i
    .io_output_r_valid                     (system_axiA_logic_axiAAdapted_r_valid                                                                    ), //i
    .io_output_r_ready                     (system_axiA_logic_bmbToAxiBridge_io_output_r_ready                                                       ), //o
    .io_output_r_payload_data              (system_axiA_logic_axiAAdapted_r_payload_data[31:0]                                                       ), //i
    .io_output_r_payload_resp              (system_axiA_logic_axiAAdapted_r_payload_resp[1:0]                                                        ), //i
    .io_output_r_payload_last              (system_axiA_logic_axiAAdapted_r_payload_last                                                             ), //i
    .io_peripheralClk                      (io_peripheralClk                                                                                         ), //i
    .peripheralCd_logic_outputReset        (peripheralCd_logic_outputReset                                                                           )  //i
  );
  BmbDecoderPerSource system_bridge_bmb_decoder (
    .io_input_cmd_valid                        (system_bridge_bmb_cmd_s2mPipe_m2sPipe_valid                               ), //i
    .io_input_cmd_ready                        (system_bridge_bmb_decoder_io_input_cmd_ready                              ), //o
    .io_input_cmd_payload_last                 (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_last                        ), //i
    .io_input_cmd_payload_fragment_source      (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_source[1:0]        ), //i
    .io_input_cmd_payload_fragment_opcode      (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_opcode             ), //i
    .io_input_cmd_payload_fragment_address     (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_address[31:0]      ), //i
    .io_input_cmd_payload_fragment_length      (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_length[5:0]        ), //i
    .io_input_cmd_payload_fragment_data        (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_data[63:0]         ), //i
    .io_input_cmd_payload_fragment_mask        (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_mask[7:0]          ), //i
    .io_input_cmd_payload_fragment_context     (system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_context[43:0]      ), //i
    .io_input_rsp_valid                        (system_bridge_bmb_decoder_io_input_rsp_valid                              ), //o
    .io_input_rsp_ready                        (system_bridge_bmb_rsp_ready                                               ), //i
    .io_input_rsp_payload_last                 (system_bridge_bmb_decoder_io_input_rsp_payload_last                       ), //o
    .io_input_rsp_payload_fragment_source      (system_bridge_bmb_decoder_io_input_rsp_payload_fragment_source[1:0]       ), //o
    .io_input_rsp_payload_fragment_opcode      (system_bridge_bmb_decoder_io_input_rsp_payload_fragment_opcode            ), //o
    .io_input_rsp_payload_fragment_data        (system_bridge_bmb_decoder_io_input_rsp_payload_fragment_data[63:0]        ), //o
    .io_input_rsp_payload_fragment_context     (system_bridge_bmb_decoder_io_input_rsp_payload_fragment_context[43:0]     ), //o
    .io_outputs_0_cmd_valid                    (system_bridge_bmb_decoder_io_outputs_0_cmd_valid                          ), //o
    .io_outputs_0_cmd_ready                    (system_bridge_bmb_unburstify_1_io_input_cmd_ready                         ), //i
    .io_outputs_0_cmd_payload_last             (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_last                   ), //o
    .io_outputs_0_cmd_payload_fragment_source  (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_source[1:0]   ), //o
    .io_outputs_0_cmd_payload_fragment_opcode  (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode        ), //o
    .io_outputs_0_cmd_payload_fragment_address (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_address[31:0] ), //o
    .io_outputs_0_cmd_payload_fragment_length  (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_length[5:0]   ), //o
    .io_outputs_0_cmd_payload_fragment_data    (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_data[63:0]    ), //o
    .io_outputs_0_cmd_payload_fragment_mask    (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_mask[7:0]     ), //o
    .io_outputs_0_cmd_payload_fragment_context (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_context[43:0] ), //o
    .io_outputs_0_rsp_valid                    (system_bridge_bmb_unburstify_1_io_input_rsp_valid                         ), //i
    .io_outputs_0_rsp_ready                    (system_bridge_bmb_decoder_io_outputs_0_rsp_ready                          ), //o
    .io_outputs_0_rsp_payload_last             (system_bridge_bmb_unburstify_1_io_input_rsp_payload_last                  ), //i
    .io_outputs_0_rsp_payload_fragment_source  (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_source[1:0]  ), //i
    .io_outputs_0_rsp_payload_fragment_opcode  (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_opcode       ), //i
    .io_outputs_0_rsp_payload_fragment_data    (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_data[63:0]   ), //i
    .io_outputs_0_rsp_payload_fragment_context (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_context[43:0]), //i
    .io_outputs_1_cmd_valid                    (system_bridge_bmb_decoder_io_outputs_1_cmd_valid                          ), //o
    .io_outputs_1_cmd_ready                    (system_bridge_bmb_downSizer_1_io_input_cmd_ready                          ), //i
    .io_outputs_1_cmd_payload_last             (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_last                   ), //o
    .io_outputs_1_cmd_payload_fragment_source  (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_source[1:0]   ), //o
    .io_outputs_1_cmd_payload_fragment_opcode  (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_opcode        ), //o
    .io_outputs_1_cmd_payload_fragment_address (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_address[31:0] ), //o
    .io_outputs_1_cmd_payload_fragment_length  (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_length[5:0]   ), //o
    .io_outputs_1_cmd_payload_fragment_data    (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_data[63:0]    ), //o
    .io_outputs_1_cmd_payload_fragment_mask    (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_mask[7:0]     ), //o
    .io_outputs_1_cmd_payload_fragment_context (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_context[43:0] ), //o
    .io_outputs_1_rsp_valid                    (system_bridge_bmb_downSizer_1_io_input_rsp_valid                          ), //i
    .io_outputs_1_rsp_ready                    (system_bridge_bmb_decoder_io_outputs_1_rsp_ready                          ), //o
    .io_outputs_1_rsp_payload_last             (system_bridge_bmb_downSizer_1_io_input_rsp_payload_last                   ), //i
    .io_outputs_1_rsp_payload_fragment_source  (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_source[1:0]   ), //i
    .io_outputs_1_rsp_payload_fragment_opcode  (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_opcode        ), //i
    .io_outputs_1_rsp_payload_fragment_data    (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_data[63:0]    ), //i
    .io_outputs_1_rsp_payload_fragment_context (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_context[43:0] ), //i
    .io_outputs_2_cmd_valid                    (system_bridge_bmb_decoder_io_outputs_2_cmd_valid                          ), //o
    .io_outputs_2_cmd_ready                    (system_bridge_bmb_upSizer_io_input_cmd_ready                              ), //i
    .io_outputs_2_cmd_payload_last             (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_last                   ), //o
    .io_outputs_2_cmd_payload_fragment_source  (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_source[1:0]   ), //o
    .io_outputs_2_cmd_payload_fragment_opcode  (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_opcode        ), //o
    .io_outputs_2_cmd_payload_fragment_address (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_address[31:0] ), //o
    .io_outputs_2_cmd_payload_fragment_length  (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_length[5:0]   ), //o
    .io_outputs_2_cmd_payload_fragment_data    (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_data[63:0]    ), //o
    .io_outputs_2_cmd_payload_fragment_mask    (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_mask[7:0]     ), //o
    .io_outputs_2_cmd_payload_fragment_context (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_context[43:0] ), //o
    .io_outputs_2_rsp_valid                    (system_bridge_bmb_upSizer_io_input_rsp_valid                              ), //i
    .io_outputs_2_rsp_ready                    (system_bridge_bmb_decoder_io_outputs_2_rsp_ready                          ), //o
    .io_outputs_2_rsp_payload_last             (system_bridge_bmb_upSizer_io_input_rsp_payload_last                       ), //i
    .io_outputs_2_rsp_payload_fragment_source  (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_source[1:0]       ), //i
    .io_outputs_2_rsp_payload_fragment_opcode  (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_opcode            ), //i
    .io_outputs_2_rsp_payload_fragment_data    (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_data[63:0]        ), //i
    .io_outputs_2_rsp_payload_fragment_context (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_context[43:0]     ), //i
    .io_outputs_3_cmd_valid                    (system_bridge_bmb_decoder_io_outputs_3_cmd_valid                          ), //o
    .io_outputs_3_cmd_ready                    (system_bridge_bmb_downSizer_io_input_cmd_ready                            ), //i
    .io_outputs_3_cmd_payload_last             (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_last                   ), //o
    .io_outputs_3_cmd_payload_fragment_source  (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_source[1:0]   ), //o
    .io_outputs_3_cmd_payload_fragment_opcode  (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_opcode        ), //o
    .io_outputs_3_cmd_payload_fragment_address (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_address[31:0] ), //o
    .io_outputs_3_cmd_payload_fragment_length  (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_length[5:0]   ), //o
    .io_outputs_3_cmd_payload_fragment_data    (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_data[63:0]    ), //o
    .io_outputs_3_cmd_payload_fragment_mask    (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_mask[7:0]     ), //o
    .io_outputs_3_cmd_payload_fragment_context (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_context[43:0] ), //o
    .io_outputs_3_rsp_valid                    (system_bridge_bmb_downSizer_io_input_rsp_valid                            ), //i
    .io_outputs_3_rsp_ready                    (system_bridge_bmb_decoder_io_outputs_3_rsp_ready                          ), //o
    .io_outputs_3_rsp_payload_last             (system_bridge_bmb_downSizer_io_input_rsp_payload_last                     ), //i
    .io_outputs_3_rsp_payload_fragment_source  (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_source[1:0]     ), //i
    .io_outputs_3_rsp_payload_fragment_opcode  (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_opcode          ), //i
    .io_outputs_3_rsp_payload_fragment_data    (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_data[63:0]      ), //i
    .io_outputs_3_rsp_payload_fragment_context (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_context[43:0]   ), //i
    .io_systemClk                              (io_systemClk                                                              ), //i
    .systemCd_logic_outputReset                (systemCd_logic_outputReset                                                )  //i
  );
  BmbUpSizerBridge system_bridge_bmb_upSizer (
    .io_input_cmd_valid                     (system_bridge_bmb_decoder_io_outputs_2_cmd_valid                                        ), //i
    .io_input_cmd_ready                     (system_bridge_bmb_upSizer_io_input_cmd_ready                                            ), //o
    .io_input_cmd_payload_last              (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_last                                 ), //i
    .io_input_cmd_payload_fragment_source   (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_source[1:0]                 ), //i
    .io_input_cmd_payload_fragment_opcode   (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_opcode                      ), //i
    .io_input_cmd_payload_fragment_address  (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_address[31:0]               ), //i
    .io_input_cmd_payload_fragment_length   (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_length[5:0]                 ), //i
    .io_input_cmd_payload_fragment_data     (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_data[63:0]                  ), //i
    .io_input_cmd_payload_fragment_mask     (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_mask[7:0]                   ), //i
    .io_input_cmd_payload_fragment_context  (system_bridge_bmb_decoder_io_outputs_2_cmd_payload_fragment_context[43:0]               ), //i
    .io_input_rsp_valid                     (system_bridge_bmb_upSizer_io_input_rsp_valid                                            ), //o
    .io_input_rsp_ready                     (system_bridge_bmb_decoder_io_outputs_2_rsp_ready                                        ), //i
    .io_input_rsp_payload_last              (system_bridge_bmb_upSizer_io_input_rsp_payload_last                                     ), //o
    .io_input_rsp_payload_fragment_source   (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_source[1:0]                     ), //o
    .io_input_rsp_payload_fragment_opcode   (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_opcode                          ), //o
    .io_input_rsp_payload_fragment_data     (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_data[63:0]                      ), //o
    .io_input_rsp_payload_fragment_context  (system_bridge_bmb_upSizer_io_input_rsp_payload_fragment_context[43:0]                   ), //o
    .io_output_cmd_valid                    (system_bridge_bmb_upSizer_io_output_cmd_valid                                           ), //o
    .io_output_cmd_ready                    (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready                         ), //i
    .io_output_cmd_payload_last             (system_bridge_bmb_upSizer_io_output_cmd_payload_last                                    ), //o
    .io_output_cmd_payload_fragment_source  (system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_source[1:0]                    ), //o
    .io_output_cmd_payload_fragment_opcode  (system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_opcode                         ), //o
    .io_output_cmd_payload_fragment_address (system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_address[31:0]                  ), //o
    .io_output_cmd_payload_fragment_length  (system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_length[5:0]                    ), //o
    .io_output_cmd_payload_fragment_data    (system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_data[127:0]                    ), //o
    .io_output_cmd_payload_fragment_mask    (system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_mask[15:0]                     ), //o
    .io_output_cmd_payload_fragment_context (system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_context[45:0]                  ), //o
    .io_output_rsp_valid                    (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid                         ), //i
    .io_output_rsp_ready                    (system_bridge_bmb_upSizer_io_output_rsp_ready                                           ), //o
    .io_output_rsp_payload_last             (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last                  ), //i
    .io_output_rsp_payload_fragment_source  (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source[1:0]  ), //i
    .io_output_rsp_payload_fragment_opcode  (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode       ), //i
    .io_output_rsp_payload_fragment_data    (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data[127:0]  ), //i
    .io_output_rsp_payload_fragment_context (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context[45:0]), //i
    .io_systemClk                           (io_systemClk                                                                            ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                                              )  //i
  );
  BmbDownSizerBridge system_bridge_bmb_downSizer (
    .io_input_cmd_valid                     (system_bridge_bmb_decoder_io_outputs_3_cmd_valid                         ), //i
    .io_input_cmd_ready                     (system_bridge_bmb_downSizer_io_input_cmd_ready                           ), //o
    .io_input_cmd_payload_last              (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_source   (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_source[1:0]  ), //i
    .io_input_cmd_payload_fragment_opcode   (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address  (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_address[31:0]), //i
    .io_input_cmd_payload_fragment_length   (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_length[5:0]  ), //i
    .io_input_cmd_payload_fragment_data     (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_data[63:0]   ), //i
    .io_input_cmd_payload_fragment_mask     (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_mask[7:0]    ), //i
    .io_input_cmd_payload_fragment_context  (system_bridge_bmb_decoder_io_outputs_3_cmd_payload_fragment_context[43:0]), //i
    .io_input_rsp_valid                     (system_bridge_bmb_downSizer_io_input_rsp_valid                           ), //o
    .io_input_rsp_ready                     (system_bridge_bmb_decoder_io_outputs_3_rsp_ready                         ), //i
    .io_input_rsp_payload_last              (system_bridge_bmb_downSizer_io_input_rsp_payload_last                    ), //o
    .io_input_rsp_payload_fragment_source   (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_source[1:0]    ), //o
    .io_input_rsp_payload_fragment_opcode   (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_opcode         ), //o
    .io_input_rsp_payload_fragment_data     (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_data[63:0]     ), //o
    .io_input_rsp_payload_fragment_context  (system_bridge_bmb_downSizer_io_input_rsp_payload_fragment_context[43:0]  ), //o
    .io_output_cmd_valid                    (system_bridge_bmb_downSizer_io_output_cmd_valid                          ), //o
    .io_output_cmd_ready                    (system_bridge_bmb_crossClock_io_input_cmd_ready                          ), //i
    .io_output_cmd_payload_last             (system_bridge_bmb_downSizer_io_output_cmd_payload_last                   ), //o
    .io_output_cmd_payload_fragment_source  (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_source[1:0]   ), //o
    .io_output_cmd_payload_fragment_opcode  (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_opcode        ), //o
    .io_output_cmd_payload_fragment_address (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_address[31:0] ), //o
    .io_output_cmd_payload_fragment_length  (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_length[5:0]   ), //o
    .io_output_cmd_payload_fragment_data    (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_data[31:0]    ), //o
    .io_output_cmd_payload_fragment_mask    (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_mask[3:0]     ), //o
    .io_output_cmd_payload_fragment_context (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_context[44:0] ), //o
    .io_output_rsp_valid                    (system_bridge_bmb_crossClock_io_input_rsp_valid                          ), //i
    .io_output_rsp_ready                    (system_bridge_bmb_downSizer_io_output_rsp_ready                          ), //o
    .io_output_rsp_payload_last             (system_bridge_bmb_crossClock_io_input_rsp_payload_last                   ), //i
    .io_output_rsp_payload_fragment_source  (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_source[1:0]   ), //i
    .io_output_rsp_payload_fragment_opcode  (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_opcode        ), //i
    .io_output_rsp_payload_fragment_data    (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_data[31:0]    ), //i
    .io_output_rsp_payload_fragment_context (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_context[44:0] ), //i
    .io_systemClk                           (io_systemClk                                                             ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                               )  //i
  );
  BmbCcFifo_1 system_bridge_bmb_crossClock (
    .io_input_cmd_valid                                                                  (system_bridge_bmb_downSizer_io_output_cmd_valid                                                                 ), //i
    .io_input_cmd_ready                                                                  (system_bridge_bmb_crossClock_io_input_cmd_ready                                                                 ), //o
    .io_input_cmd_payload_last                                                           (system_bridge_bmb_downSizer_io_output_cmd_payload_last                                                          ), //i
    .io_input_cmd_payload_fragment_source                                                (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_source[1:0]                                          ), //i
    .io_input_cmd_payload_fragment_opcode                                                (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_opcode                                               ), //i
    .io_input_cmd_payload_fragment_address                                               (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_address[31:0]                                        ), //i
    .io_input_cmd_payload_fragment_length                                                (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_length[5:0]                                          ), //i
    .io_input_cmd_payload_fragment_data                                                  (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_data[31:0]                                           ), //i
    .io_input_cmd_payload_fragment_mask                                                  (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_mask[3:0]                                            ), //i
    .io_input_cmd_payload_fragment_context                                               (system_bridge_bmb_downSizer_io_output_cmd_payload_fragment_context[44:0]                                        ), //i
    .io_input_rsp_valid                                                                  (system_bridge_bmb_crossClock_io_input_rsp_valid                                                                 ), //o
    .io_input_rsp_ready                                                                  (system_bridge_bmb_downSizer_io_output_rsp_ready                                                                 ), //i
    .io_input_rsp_payload_last                                                           (system_bridge_bmb_crossClock_io_input_rsp_payload_last                                                          ), //o
    .io_input_rsp_payload_fragment_source                                                (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_source[1:0]                                          ), //o
    .io_input_rsp_payload_fragment_opcode                                                (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_opcode                                               ), //o
    .io_input_rsp_payload_fragment_data                                                  (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_data[31:0]                                           ), //o
    .io_input_rsp_payload_fragment_context                                               (system_bridge_bmb_crossClock_io_input_rsp_payload_fragment_context[44:0]                                        ), //o
    .io_output_cmd_valid                                                                 (system_bridge_bmb_crossClock_io_output_cmd_valid                                                                ), //o
    .io_output_cmd_ready                                                                 (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready                                                ), //i
    .io_output_cmd_payload_last                                                          (system_bridge_bmb_crossClock_io_output_cmd_payload_last                                                         ), //o
    .io_output_cmd_payload_fragment_source                                               (system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_source[1:0]                                         ), //o
    .io_output_cmd_payload_fragment_opcode                                               (system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_opcode                                              ), //o
    .io_output_cmd_payload_fragment_address                                              (system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_address[31:0]                                       ), //o
    .io_output_cmd_payload_fragment_length                                               (system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_length[5:0]                                         ), //o
    .io_output_cmd_payload_fragment_data                                                 (system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_data[31:0]                                          ), //o
    .io_output_cmd_payload_fragment_mask                                                 (system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_mask[3:0]                                           ), //o
    .io_output_cmd_payload_fragment_context                                              (system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_context[44:0]                                       ), //o
    .io_output_rsp_valid                                                                 (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid                                                ), //i
    .io_output_rsp_ready                                                                 (system_bridge_bmb_crossClock_io_output_rsp_ready                                                                ), //o
    .io_output_rsp_payload_last                                                          (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last                                         ), //i
    .io_output_rsp_payload_fragment_source                                               (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source[1:0]                         ), //i
    .io_output_rsp_payload_fragment_opcode                                               (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode                              ), //i
    .io_output_rsp_payload_fragment_data                                                 (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data[31:0]                          ), //i
    .io_output_rsp_payload_fragment_context                                              (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context[44:0]                       ), //i
    .io_systemClk                                                                        (io_systemClk                                                                                                    ), //i
    .systemCd_logic_outputReset                                                          (systemCd_logic_outputReset                                                                                      ), //i
    .io_peripheralClk                                                                    (io_peripheralClk                                                                                                ), //i
    .peripheralCd_logic_outputReset                                                      (peripheralCd_logic_outputReset                                                                                  ), //i
    .system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1     (system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1    ), //o
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //o
  );
  BmbOnChipRam system_ramA_logic (
    .io_bus_cmd_valid                    (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_valid                         ), //i
    .io_bus_cmd_ready                    (system_ramA_logic_io_bus_cmd_ready                                                                  ), //o
    .io_bus_cmd_payload_last             (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_last                  ), //i
    .io_bus_cmd_payload_fragment_opcode  (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_opcode       ), //i
    .io_bus_cmd_payload_fragment_address (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_address[10:0]), //i
    .io_bus_cmd_payload_fragment_length  (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_length[2:0]  ), //i
    .io_bus_cmd_payload_fragment_data    (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_data[63:0]   ), //i
    .io_bus_cmd_payload_fragment_mask    (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_mask[7:0]    ), //i
    .io_bus_cmd_payload_fragment_context (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_context[47:0]), //i
    .io_bus_rsp_valid                    (system_ramA_logic_io_bus_rsp_valid                                                                  ), //o
    .io_bus_rsp_ready                    (_zz_io_bus_rsp_ready                                                                                ), //i
    .io_bus_rsp_payload_last             (system_ramA_logic_io_bus_rsp_payload_last                                                           ), //o
    .io_bus_rsp_payload_fragment_opcode  (system_ramA_logic_io_bus_rsp_payload_fragment_opcode                                                ), //o
    .io_bus_rsp_payload_fragment_data    (system_ramA_logic_io_bus_rsp_payload_fragment_data[63:0]                                            ), //o
    .io_bus_rsp_payload_fragment_context (system_ramA_logic_io_bus_rsp_payload_fragment_context[47:0]                                         ), //o
    .io_systemClk                        (io_systemClk                                                                                        ), //i
    .systemCd_logic_outputReset          (systemCd_logic_outputReset                                                                          )  //i
  );
  BmbDownSizerBridge system_bridge_bmb_downSizer_1 (
    .io_input_cmd_valid                     (system_bridge_bmb_decoder_io_outputs_1_cmd_valid                          ), //i
    .io_input_cmd_ready                     (system_bridge_bmb_downSizer_1_io_input_cmd_ready                          ), //o
    .io_input_cmd_payload_last              (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_last                   ), //i
    .io_input_cmd_payload_fragment_source   (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_source[1:0]   ), //i
    .io_input_cmd_payload_fragment_opcode   (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_opcode        ), //i
    .io_input_cmd_payload_fragment_address  (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_address[31:0] ), //i
    .io_input_cmd_payload_fragment_length   (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_length[5:0]   ), //i
    .io_input_cmd_payload_fragment_data     (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_data[63:0]    ), //i
    .io_input_cmd_payload_fragment_mask     (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_mask[7:0]     ), //i
    .io_input_cmd_payload_fragment_context  (system_bridge_bmb_decoder_io_outputs_1_cmd_payload_fragment_context[43:0] ), //i
    .io_input_rsp_valid                     (system_bridge_bmb_downSizer_1_io_input_rsp_valid                          ), //o
    .io_input_rsp_ready                     (system_bridge_bmb_decoder_io_outputs_1_rsp_ready                          ), //i
    .io_input_rsp_payload_last              (system_bridge_bmb_downSizer_1_io_input_rsp_payload_last                   ), //o
    .io_input_rsp_payload_fragment_source   (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_source[1:0]   ), //o
    .io_input_rsp_payload_fragment_opcode   (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_opcode        ), //o
    .io_input_rsp_payload_fragment_data     (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_data[63:0]    ), //o
    .io_input_rsp_payload_fragment_context  (system_bridge_bmb_downSizer_1_io_input_rsp_payload_fragment_context[43:0] ), //o
    .io_output_cmd_valid                    (system_bridge_bmb_downSizer_1_io_output_cmd_valid                         ), //o
    .io_output_cmd_ready                    (system_bridge_bmb_unburstify_io_input_cmd_ready                           ), //i
    .io_output_cmd_payload_last             (system_bridge_bmb_downSizer_1_io_output_cmd_payload_last                  ), //o
    .io_output_cmd_payload_fragment_source  (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_source[1:0]  ), //o
    .io_output_cmd_payload_fragment_opcode  (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_opcode       ), //o
    .io_output_cmd_payload_fragment_address (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_address[31:0]), //o
    .io_output_cmd_payload_fragment_length  (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_length[5:0]  ), //o
    .io_output_cmd_payload_fragment_data    (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_data[31:0]   ), //o
    .io_output_cmd_payload_fragment_mask    (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_mask[3:0]    ), //o
    .io_output_cmd_payload_fragment_context (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_context[44:0]), //o
    .io_output_rsp_valid                    (system_bridge_bmb_unburstify_io_input_rsp_valid                           ), //i
    .io_output_rsp_ready                    (system_bridge_bmb_downSizer_1_io_output_rsp_ready                         ), //o
    .io_output_rsp_payload_last             (system_bridge_bmb_unburstify_io_input_rsp_payload_last                    ), //i
    .io_output_rsp_payload_fragment_source  (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_source[1:0]    ), //i
    .io_output_rsp_payload_fragment_opcode  (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_opcode         ), //i
    .io_output_rsp_payload_fragment_data    (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_data[31:0]     ), //i
    .io_output_rsp_payload_fragment_context (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_context[44:0]  ), //i
    .io_systemClk                           (io_systemClk                                                              ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                                )  //i
  );
  BmbUnburstify system_bridge_bmb_unburstify (
    .io_input_cmd_valid                     (system_bridge_bmb_downSizer_1_io_output_cmd_valid                         ), //i
    .io_input_cmd_ready                     (system_bridge_bmb_unburstify_io_input_cmd_ready                           ), //o
    .io_input_cmd_payload_last              (system_bridge_bmb_downSizer_1_io_output_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_source   (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_source[1:0]  ), //i
    .io_input_cmd_payload_fragment_opcode   (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address  (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_address[31:0]), //i
    .io_input_cmd_payload_fragment_length   (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_length[5:0]  ), //i
    .io_input_cmd_payload_fragment_data     (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_data[31:0]   ), //i
    .io_input_cmd_payload_fragment_mask     (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_mask[3:0]    ), //i
    .io_input_cmd_payload_fragment_context  (system_bridge_bmb_downSizer_1_io_output_cmd_payload_fragment_context[44:0]), //i
    .io_input_rsp_valid                     (system_bridge_bmb_unburstify_io_input_rsp_valid                           ), //o
    .io_input_rsp_ready                     (system_bridge_bmb_downSizer_1_io_output_rsp_ready                         ), //i
    .io_input_rsp_payload_last              (system_bridge_bmb_unburstify_io_input_rsp_payload_last                    ), //o
    .io_input_rsp_payload_fragment_source   (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_source[1:0]    ), //o
    .io_input_rsp_payload_fragment_opcode   (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_opcode         ), //o
    .io_input_rsp_payload_fragment_data     (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_data[31:0]     ), //o
    .io_input_rsp_payload_fragment_context  (system_bridge_bmb_unburstify_io_input_rsp_payload_fragment_context[44:0]  ), //o
    .io_output_cmd_valid                    (system_bridge_bmb_unburstify_io_output_cmd_valid                          ), //o
    .io_output_cmd_ready                    (system_bridge_bmb_crossClock_1_io_input_cmd_ready                         ), //i
    .io_output_cmd_payload_last             (system_bridge_bmb_unburstify_io_output_cmd_payload_last                   ), //o
    .io_output_cmd_payload_fragment_opcode  (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_opcode        ), //o
    .io_output_cmd_payload_fragment_address (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_address[31:0] ), //o
    .io_output_cmd_payload_fragment_length  (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_length[1:0]   ), //o
    .io_output_cmd_payload_fragment_data    (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_data[31:0]    ), //o
    .io_output_cmd_payload_fragment_mask    (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_mask[3:0]     ), //o
    .io_output_cmd_payload_fragment_context (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_context[48:0] ), //o
    .io_output_rsp_valid                    (system_bridge_bmb_crossClock_1_io_input_rsp_valid                         ), //i
    .io_output_rsp_ready                    (system_bridge_bmb_unburstify_io_output_rsp_ready                          ), //o
    .io_output_rsp_payload_last             (system_bridge_bmb_crossClock_1_io_input_rsp_payload_last                  ), //i
    .io_output_rsp_payload_fragment_opcode  (system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_opcode       ), //i
    .io_output_rsp_payload_fragment_data    (system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_data[31:0]   ), //i
    .io_output_rsp_payload_fragment_context (system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_context[48:0]), //i
    .io_systemClk                           (io_systemClk                                                              ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                                )  //i
  );
  BmbCcToggle system_bridge_bmb_crossClock_1 (
    .io_input_cmd_valid                                                                  (system_bridge_bmb_unburstify_io_output_cmd_valid                                                                ), //i
    .io_input_cmd_ready                                                                  (system_bridge_bmb_crossClock_1_io_input_cmd_ready                                                               ), //o
    .io_input_cmd_payload_last                                                           (system_bridge_bmb_unburstify_io_output_cmd_payload_last                                                         ), //i
    .io_input_cmd_payload_fragment_opcode                                                (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_opcode                                              ), //i
    .io_input_cmd_payload_fragment_address                                               (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_address[31:0]                                       ), //i
    .io_input_cmd_payload_fragment_length                                                (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_length[1:0]                                         ), //i
    .io_input_cmd_payload_fragment_data                                                  (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_data[31:0]                                          ), //i
    .io_input_cmd_payload_fragment_mask                                                  (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_mask[3:0]                                           ), //i
    .io_input_cmd_payload_fragment_context                                               (system_bridge_bmb_unburstify_io_output_cmd_payload_fragment_context[48:0]                                       ), //i
    .io_input_rsp_valid                                                                  (system_bridge_bmb_crossClock_1_io_input_rsp_valid                                                               ), //o
    .io_input_rsp_ready                                                                  (system_bridge_bmb_unburstify_io_output_rsp_ready                                                                ), //i
    .io_input_rsp_payload_last                                                           (system_bridge_bmb_crossClock_1_io_input_rsp_payload_last                                                        ), //o
    .io_input_rsp_payload_fragment_opcode                                                (system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_opcode                                             ), //o
    .io_input_rsp_payload_fragment_data                                                  (system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_data[31:0]                                         ), //o
    .io_input_rsp_payload_fragment_context                                               (system_bridge_bmb_crossClock_1_io_input_rsp_payload_fragment_context[48:0]                                      ), //o
    .io_output_cmd_valid                                                                 (system_bridge_bmb_crossClock_1_io_output_cmd_valid                                                              ), //o
    .io_output_cmd_ready                                                                 (system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready                                       ), //i
    .io_output_cmd_payload_last                                                          (system_bridge_bmb_crossClock_1_io_output_cmd_payload_last                                                       ), //o
    .io_output_cmd_payload_fragment_opcode                                               (system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_opcode                                            ), //o
    .io_output_cmd_payload_fragment_address                                              (system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_address[31:0]                                     ), //o
    .io_output_cmd_payload_fragment_length                                               (system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_length[1:0]                                       ), //o
    .io_output_cmd_payload_fragment_data                                                 (system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_data[31:0]                                        ), //o
    .io_output_cmd_payload_fragment_mask                                                 (system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_mask[3:0]                                         ), //o
    .io_output_cmd_payload_fragment_context                                              (system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_context[48:0]                                     ), //o
    .io_output_rsp_valid                                                                 (system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid                                       ), //i
    .io_output_rsp_ready                                                                 (system_bridge_bmb_crossClock_1_io_output_rsp_ready                                                              ), //o
    .io_output_rsp_payload_last                                                          (system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last                                ), //i
    .io_output_rsp_payload_fragment_opcode                                               (system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode                     ), //i
    .io_output_rsp_payload_fragment_data                                                 (system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data[31:0]                 ), //i
    .io_output_rsp_payload_fragment_context                                              (system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context[48:0]              ), //i
    .io_systemClk                                                                        (io_systemClk                                                                                                    ), //i
    .systemCd_logic_outputReset                                                          (systemCd_logic_outputReset                                                                                      ), //i
    .io_peripheralClk                                                                    (io_peripheralClk                                                                                                ), //i
    .system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1     (system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1    ), //i
    .peripheralCd_logic_outputReset                                                      (peripheralCd_logic_outputReset                                                                                  ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //i
  );
  BmbUnburstify_1 system_bridge_bmb_unburstify_1 (
    .io_input_cmd_valid                     (system_bridge_bmb_decoder_io_outputs_0_cmd_valid                                          ), //i
    .io_input_cmd_ready                     (system_bridge_bmb_unburstify_1_io_input_cmd_ready                                         ), //o
    .io_input_cmd_payload_last              (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_last                                   ), //i
    .io_input_cmd_payload_fragment_source   (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_source[1:0]                   ), //i
    .io_input_cmd_payload_fragment_opcode   (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode                        ), //i
    .io_input_cmd_payload_fragment_address  (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_address[31:0]                 ), //i
    .io_input_cmd_payload_fragment_length   (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_length[5:0]                   ), //i
    .io_input_cmd_payload_fragment_data     (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_data[63:0]                    ), //i
    .io_input_cmd_payload_fragment_mask     (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_mask[7:0]                     ), //i
    .io_input_cmd_payload_fragment_context  (system_bridge_bmb_decoder_io_outputs_0_cmd_payload_fragment_context[43:0]                 ), //i
    .io_input_rsp_valid                     (system_bridge_bmb_unburstify_1_io_input_rsp_valid                                         ), //o
    .io_input_rsp_ready                     (system_bridge_bmb_decoder_io_outputs_0_rsp_ready                                          ), //i
    .io_input_rsp_payload_last              (system_bridge_bmb_unburstify_1_io_input_rsp_payload_last                                  ), //o
    .io_input_rsp_payload_fragment_source   (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_source[1:0]                  ), //o
    .io_input_rsp_payload_fragment_opcode   (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_opcode                       ), //o
    .io_input_rsp_payload_fragment_data     (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_data[63:0]                   ), //o
    .io_input_rsp_payload_fragment_context  (system_bridge_bmb_unburstify_1_io_input_rsp_payload_fragment_context[43:0]                ), //o
    .io_output_cmd_valid                    (system_bridge_bmb_unburstify_1_io_output_cmd_valid                                        ), //o
    .io_output_cmd_ready                    (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready                         ), //i
    .io_output_cmd_payload_last             (system_bridge_bmb_unburstify_1_io_output_cmd_payload_last                                 ), //o
    .io_output_cmd_payload_fragment_opcode  (system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_opcode                      ), //o
    .io_output_cmd_payload_fragment_address (system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_address[31:0]               ), //o
    .io_output_cmd_payload_fragment_length  (system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_length[2:0]                 ), //o
    .io_output_cmd_payload_fragment_data    (system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_data[63:0]                  ), //o
    .io_output_cmd_payload_fragment_mask    (system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_mask[7:0]                   ), //o
    .io_output_cmd_payload_fragment_context (system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_context[47:0]               ), //o
    .io_output_rsp_valid                    (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid                         ), //i
    .io_output_rsp_ready                    (system_bridge_bmb_unburstify_1_io_output_rsp_ready                                        ), //o
    .io_output_rsp_payload_last             (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last                  ), //i
    .io_output_rsp_payload_fragment_opcode  (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode       ), //i
    .io_output_rsp_payload_fragment_data    (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data[63:0]   ), //i
    .io_output_rsp_payload_fragment_context (system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context[47:0]), //i
    .io_systemClk                           (io_systemClk                                                                              ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                                                )  //i
  );
  BmbDecoder_1 system_bmbPeripheral_bmb_decoder (
    .io_input_cmd_valid                         (system_bmbPeripheral_bmb_cmd_combStage_valid                                     ), //i
    .io_input_cmd_ready                         (system_bmbPeripheral_bmb_decoder_io_input_cmd_ready                              ), //o
    .io_input_cmd_payload_last                  (system_bmbPeripheral_bmb_cmd_combStage_payload_last                              ), //i
    .io_input_cmd_payload_fragment_opcode       (system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_opcode                   ), //i
    .io_input_cmd_payload_fragment_address      (system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_address[23:0]            ), //i
    .io_input_cmd_payload_fragment_length       (system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_length[1:0]              ), //i
    .io_input_cmd_payload_fragment_data         (system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_data[31:0]               ), //i
    .io_input_cmd_payload_fragment_mask         (system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_mask[3:0]                ), //i
    .io_input_cmd_payload_fragment_context      (system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_context[48:0]            ), //i
    .io_input_rsp_valid                         (system_bmbPeripheral_bmb_decoder_io_input_rsp_valid                              ), //o
    .io_input_rsp_ready                         (_zz_io_input_rsp_ready_4                                                         ), //i
    .io_input_rsp_payload_last                  (system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_last                       ), //o
    .io_input_rsp_payload_fragment_opcode       (system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_opcode            ), //o
    .io_input_rsp_payload_fragment_data         (system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_data[31:0]        ), //o
    .io_input_rsp_payload_fragment_context      (system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_context[48:0]     ), //o
    .io_outputs_0_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_valid                          ), //o
    .io_outputs_0_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_16                                ), //i
    .io_outputs_0_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_last                   ), //o
    .io_outputs_0_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode        ), //o
    .io_outputs_0_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_0_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_0_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_0_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_0_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_0_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_16                                ), //i
    .io_outputs_0_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_0_rsp_ready                          ), //o
    .io_outputs_0_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_16                         ), //i
    .io_outputs_0_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_16              ), //i
    .io_outputs_0_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_16[31:0]          ), //i
    .io_outputs_0_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_16[48:0]       ), //i
    .io_outputs_1_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_valid                          ), //o
    .io_outputs_1_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready                                   ), //i
    .io_outputs_1_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_last                   ), //o
    .io_outputs_1_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_opcode        ), //o
    .io_outputs_1_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_1_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_1_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_1_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_1_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_1_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid                                   ), //i
    .io_outputs_1_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_1_rsp_ready                          ), //o
    .io_outputs_1_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last                            ), //i
    .io_outputs_1_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode                 ), //i
    .io_outputs_1_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data[31:0]             ), //i
    .io_outputs_1_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context[48:0]          ), //i
    .io_outputs_2_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_valid                          ), //o
    .io_outputs_2_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_1                                 ), //i
    .io_outputs_2_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_last                   ), //o
    .io_outputs_2_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_opcode        ), //o
    .io_outputs_2_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_2_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_2_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_2_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_2_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_2_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_1                                 ), //i
    .io_outputs_2_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_2_rsp_ready                          ), //o
    .io_outputs_2_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_1                          ), //i
    .io_outputs_2_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_1               ), //i
    .io_outputs_2_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_1[31:0]           ), //i
    .io_outputs_2_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_1[48:0]        ), //i
    .io_outputs_3_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_valid                          ), //o
    .io_outputs_3_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_2                                 ), //i
    .io_outputs_3_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_last                   ), //o
    .io_outputs_3_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_opcode        ), //o
    .io_outputs_3_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_3_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_3_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_3_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_3_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_3_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_2                                 ), //i
    .io_outputs_3_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_3_rsp_ready                          ), //o
    .io_outputs_3_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_2                          ), //i
    .io_outputs_3_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_2               ), //i
    .io_outputs_3_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_2[31:0]           ), //i
    .io_outputs_3_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_2[48:0]        ), //i
    .io_outputs_4_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_valid                          ), //o
    .io_outputs_4_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_3                                 ), //i
    .io_outputs_4_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_last                   ), //o
    .io_outputs_4_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_opcode        ), //o
    .io_outputs_4_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_4_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_4_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_4_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_4_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_4_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_3                                 ), //i
    .io_outputs_4_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_4_rsp_ready                          ), //o
    .io_outputs_4_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_3                          ), //i
    .io_outputs_4_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_3               ), //i
    .io_outputs_4_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_3[31:0]           ), //i
    .io_outputs_4_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_3[48:0]        ), //i
    .io_outputs_5_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_valid                          ), //o
    .io_outputs_5_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_4                                 ), //i
    .io_outputs_5_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_last                   ), //o
    .io_outputs_5_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_opcode        ), //o
    .io_outputs_5_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_5_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_5_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_5_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_5_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_5_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_4                                 ), //i
    .io_outputs_5_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_5_rsp_ready                          ), //o
    .io_outputs_5_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_4                          ), //i
    .io_outputs_5_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_4               ), //i
    .io_outputs_5_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_4[31:0]           ), //i
    .io_outputs_5_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_4[48:0]        ), //i
    .io_outputs_6_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_valid                          ), //o
    .io_outputs_6_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_5                                 ), //i
    .io_outputs_6_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_last                   ), //o
    .io_outputs_6_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_opcode        ), //o
    .io_outputs_6_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_6_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_6_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_6_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_6_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_6_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_5                                 ), //i
    .io_outputs_6_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_6_rsp_ready                          ), //o
    .io_outputs_6_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_5                          ), //i
    .io_outputs_6_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_5               ), //i
    .io_outputs_6_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_5[31:0]           ), //i
    .io_outputs_6_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_5[48:0]        ), //i
    .io_outputs_7_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_valid                          ), //o
    .io_outputs_7_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_6                                 ), //i
    .io_outputs_7_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_last                   ), //o
    .io_outputs_7_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_opcode        ), //o
    .io_outputs_7_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_7_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_7_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_7_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_7_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_7_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_6                                 ), //i
    .io_outputs_7_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_7_rsp_ready                          ), //o
    .io_outputs_7_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_6                          ), //i
    .io_outputs_7_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_6               ), //i
    .io_outputs_7_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_6[31:0]           ), //i
    .io_outputs_7_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_6[48:0]        ), //i
    .io_outputs_8_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_valid                          ), //o
    .io_outputs_8_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_7                                 ), //i
    .io_outputs_8_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_last                   ), //o
    .io_outputs_8_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_opcode        ), //o
    .io_outputs_8_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_8_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_8_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_8_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_8_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_8_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_7                                 ), //i
    .io_outputs_8_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_8_rsp_ready                          ), //o
    .io_outputs_8_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_7                          ), //i
    .io_outputs_8_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_7               ), //i
    .io_outputs_8_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_7[31:0]           ), //i
    .io_outputs_8_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_7[48:0]        ), //i
    .io_outputs_9_cmd_valid                     (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_valid                          ), //o
    .io_outputs_9_cmd_ready                     (system_bmbPeripheral_bmb_withoutMask_cmd_ready_8                                 ), //i
    .io_outputs_9_cmd_payload_last              (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_last                   ), //o
    .io_outputs_9_cmd_payload_fragment_opcode   (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_opcode        ), //o
    .io_outputs_9_cmd_payload_fragment_address  (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_address[23:0] ), //o
    .io_outputs_9_cmd_payload_fragment_length   (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_length[1:0]   ), //o
    .io_outputs_9_cmd_payload_fragment_data     (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_data[31:0]    ), //o
    .io_outputs_9_cmd_payload_fragment_mask     (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_mask[3:0]     ), //o
    .io_outputs_9_cmd_payload_fragment_context  (system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_context[48:0] ), //o
    .io_outputs_9_rsp_valid                     (system_bmbPeripheral_bmb_withoutMask_rsp_valid_8                                 ), //i
    .io_outputs_9_rsp_ready                     (system_bmbPeripheral_bmb_decoder_io_outputs_9_rsp_ready                          ), //o
    .io_outputs_9_rsp_payload_last              (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_8                          ), //i
    .io_outputs_9_rsp_payload_fragment_opcode   (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_8               ), //i
    .io_outputs_9_rsp_payload_fragment_data     (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_8[31:0]           ), //i
    .io_outputs_9_rsp_payload_fragment_context  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_8[48:0]        ), //i
    .io_outputs_10_cmd_valid                    (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_valid                         ), //o
    .io_outputs_10_cmd_ready                    (system_bmbPeripheral_bmb_withoutMask_cmd_ready_9                                 ), //i
    .io_outputs_10_cmd_payload_last             (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_last                  ), //o
    .io_outputs_10_cmd_payload_fragment_opcode  (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_opcode       ), //o
    .io_outputs_10_cmd_payload_fragment_address (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_address[23:0]), //o
    .io_outputs_10_cmd_payload_fragment_length  (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_length[1:0]  ), //o
    .io_outputs_10_cmd_payload_fragment_data    (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_data[31:0]   ), //o
    .io_outputs_10_cmd_payload_fragment_mask    (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_mask[3:0]    ), //o
    .io_outputs_10_cmd_payload_fragment_context (system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_context[48:0]), //o
    .io_outputs_10_rsp_valid                    (system_bmbPeripheral_bmb_withoutMask_rsp_valid_9                                 ), //i
    .io_outputs_10_rsp_ready                    (system_bmbPeripheral_bmb_decoder_io_outputs_10_rsp_ready                         ), //o
    .io_outputs_10_rsp_payload_last             (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_9                          ), //i
    .io_outputs_10_rsp_payload_fragment_opcode  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_9               ), //i
    .io_outputs_10_rsp_payload_fragment_data    (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_9[31:0]           ), //i
    .io_outputs_10_rsp_payload_fragment_context (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_9[48:0]        ), //i
    .io_outputs_11_cmd_valid                    (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_valid                         ), //o
    .io_outputs_11_cmd_ready                    (system_bmbPeripheral_bmb_withoutMask_cmd_ready_10                                ), //i
    .io_outputs_11_cmd_payload_last             (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_last                  ), //o
    .io_outputs_11_cmd_payload_fragment_opcode  (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_opcode       ), //o
    .io_outputs_11_cmd_payload_fragment_address (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_address[23:0]), //o
    .io_outputs_11_cmd_payload_fragment_length  (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_length[1:0]  ), //o
    .io_outputs_11_cmd_payload_fragment_data    (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_data[31:0]   ), //o
    .io_outputs_11_cmd_payload_fragment_mask    (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_mask[3:0]    ), //o
    .io_outputs_11_cmd_payload_fragment_context (system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_context[48:0]), //o
    .io_outputs_11_rsp_valid                    (system_bmbPeripheral_bmb_withoutMask_rsp_valid_10                                ), //i
    .io_outputs_11_rsp_ready                    (system_bmbPeripheral_bmb_decoder_io_outputs_11_rsp_ready                         ), //o
    .io_outputs_11_rsp_payload_last             (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_10                         ), //i
    .io_outputs_11_rsp_payload_fragment_opcode  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_10              ), //i
    .io_outputs_11_rsp_payload_fragment_data    (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_10[31:0]          ), //i
    .io_outputs_11_rsp_payload_fragment_context (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_10[48:0]       ), //i
    .io_outputs_12_cmd_valid                    (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_valid                         ), //o
    .io_outputs_12_cmd_ready                    (system_bmbPeripheral_bmb_withoutMask_cmd_ready_11                                ), //i
    .io_outputs_12_cmd_payload_last             (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_last                  ), //o
    .io_outputs_12_cmd_payload_fragment_opcode  (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_opcode       ), //o
    .io_outputs_12_cmd_payload_fragment_address (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_address[23:0]), //o
    .io_outputs_12_cmd_payload_fragment_length  (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_length[1:0]  ), //o
    .io_outputs_12_cmd_payload_fragment_data    (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_data[31:0]   ), //o
    .io_outputs_12_cmd_payload_fragment_mask    (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_mask[3:0]    ), //o
    .io_outputs_12_cmd_payload_fragment_context (system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_context[48:0]), //o
    .io_outputs_12_rsp_valid                    (system_bmbPeripheral_bmb_withoutMask_rsp_valid_11                                ), //i
    .io_outputs_12_rsp_ready                    (system_bmbPeripheral_bmb_decoder_io_outputs_12_rsp_ready                         ), //o
    .io_outputs_12_rsp_payload_last             (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_11                         ), //i
    .io_outputs_12_rsp_payload_fragment_opcode  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_11              ), //i
    .io_outputs_12_rsp_payload_fragment_data    (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_11[31:0]          ), //i
    .io_outputs_12_rsp_payload_fragment_context (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_11[48:0]       ), //i
    .io_outputs_13_cmd_valid                    (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_valid                         ), //o
    .io_outputs_13_cmd_ready                    (system_bmbPeripheral_bmb_withoutMask_cmd_ready_12                                ), //i
    .io_outputs_13_cmd_payload_last             (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_last                  ), //o
    .io_outputs_13_cmd_payload_fragment_opcode  (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_opcode       ), //o
    .io_outputs_13_cmd_payload_fragment_address (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_address[23:0]), //o
    .io_outputs_13_cmd_payload_fragment_length  (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_length[1:0]  ), //o
    .io_outputs_13_cmd_payload_fragment_data    (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_data[31:0]   ), //o
    .io_outputs_13_cmd_payload_fragment_mask    (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_mask[3:0]    ), //o
    .io_outputs_13_cmd_payload_fragment_context (system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_context[48:0]), //o
    .io_outputs_13_rsp_valid                    (system_bmbPeripheral_bmb_withoutMask_rsp_valid_12                                ), //i
    .io_outputs_13_rsp_ready                    (system_bmbPeripheral_bmb_decoder_io_outputs_13_rsp_ready                         ), //o
    .io_outputs_13_rsp_payload_last             (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_12                         ), //i
    .io_outputs_13_rsp_payload_fragment_opcode  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_12              ), //i
    .io_outputs_13_rsp_payload_fragment_data    (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_12[31:0]          ), //i
    .io_outputs_13_rsp_payload_fragment_context (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_12[48:0]       ), //i
    .io_outputs_14_cmd_valid                    (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_valid                         ), //o
    .io_outputs_14_cmd_ready                    (system_bmbPeripheral_bmb_withoutMask_cmd_ready_13                                ), //i
    .io_outputs_14_cmd_payload_last             (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_last                  ), //o
    .io_outputs_14_cmd_payload_fragment_opcode  (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_opcode       ), //o
    .io_outputs_14_cmd_payload_fragment_address (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_address[23:0]), //o
    .io_outputs_14_cmd_payload_fragment_length  (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_length[1:0]  ), //o
    .io_outputs_14_cmd_payload_fragment_data    (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_data[31:0]   ), //o
    .io_outputs_14_cmd_payload_fragment_mask    (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_mask[3:0]    ), //o
    .io_outputs_14_cmd_payload_fragment_context (system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_context[48:0]), //o
    .io_outputs_14_rsp_valid                    (system_bmbPeripheral_bmb_withoutMask_rsp_valid_13                                ), //i
    .io_outputs_14_rsp_ready                    (system_bmbPeripheral_bmb_decoder_io_outputs_14_rsp_ready                         ), //o
    .io_outputs_14_rsp_payload_last             (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_13                         ), //i
    .io_outputs_14_rsp_payload_fragment_opcode  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_13              ), //i
    .io_outputs_14_rsp_payload_fragment_data    (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_13[31:0]          ), //i
    .io_outputs_14_rsp_payload_fragment_context (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_13[48:0]       ), //i
    .io_outputs_15_cmd_valid                    (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_valid                         ), //o
    .io_outputs_15_cmd_ready                    (system_bmbPeripheral_bmb_withoutMask_cmd_ready_14                                ), //i
    .io_outputs_15_cmd_payload_last             (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_last                  ), //o
    .io_outputs_15_cmd_payload_fragment_opcode  (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_opcode       ), //o
    .io_outputs_15_cmd_payload_fragment_address (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_address[23:0]), //o
    .io_outputs_15_cmd_payload_fragment_length  (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_length[1:0]  ), //o
    .io_outputs_15_cmd_payload_fragment_data    (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_data[31:0]   ), //o
    .io_outputs_15_cmd_payload_fragment_mask    (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_mask[3:0]    ), //o
    .io_outputs_15_cmd_payload_fragment_context (system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_context[48:0]), //o
    .io_outputs_15_rsp_valid                    (system_bmbPeripheral_bmb_withoutMask_rsp_valid_14                                ), //i
    .io_outputs_15_rsp_ready                    (system_bmbPeripheral_bmb_decoder_io_outputs_15_rsp_ready                         ), //o
    .io_outputs_15_rsp_payload_last             (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_14                         ), //i
    .io_outputs_15_rsp_payload_fragment_opcode  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_14              ), //i
    .io_outputs_15_rsp_payload_fragment_data    (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_14[31:0]          ), //i
    .io_outputs_15_rsp_payload_fragment_context (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_14[48:0]       ), //i
    .io_outputs_16_cmd_valid                    (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_valid                         ), //o
    .io_outputs_16_cmd_ready                    (system_bmbPeripheral_bmb_withoutMask_cmd_ready_15                                ), //i
    .io_outputs_16_cmd_payload_last             (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_last                  ), //o
    .io_outputs_16_cmd_payload_fragment_opcode  (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_opcode       ), //o
    .io_outputs_16_cmd_payload_fragment_address (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_address[23:0]), //o
    .io_outputs_16_cmd_payload_fragment_length  (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_length[1:0]  ), //o
    .io_outputs_16_cmd_payload_fragment_data    (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_data[31:0]   ), //o
    .io_outputs_16_cmd_payload_fragment_mask    (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_mask[3:0]    ), //o
    .io_outputs_16_cmd_payload_fragment_context (system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_context[48:0]), //o
    .io_outputs_16_rsp_valid                    (system_bmbPeripheral_bmb_withoutMask_rsp_valid_15                                ), //i
    .io_outputs_16_rsp_ready                    (system_bmbPeripheral_bmb_decoder_io_outputs_16_rsp_ready                         ), //o
    .io_outputs_16_rsp_payload_last             (system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_15                         ), //i
    .io_outputs_16_rsp_payload_fragment_opcode  (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_15              ), //i
    .io_outputs_16_rsp_payload_fragment_data    (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_15[31:0]          ), //i
    .io_outputs_16_rsp_payload_fragment_context (system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_15[48:0]       ), //i
    .io_peripheralClk                           (io_peripheralClk                                                                 ), //i
    .peripheralCd_logic_outputReset             (peripheralCd_logic_outputReset                                                   )  //i
  );
  BmbClint system_clint_logic (
    .io_bus_cmd_valid                    (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_bus_cmd_ready                    (system_clint_logic_io_bus_cmd_ready                                                        ), //o
    .io_bus_cmd_payload_last             (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_bus_cmd_payload_fragment_opcode  (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_bus_cmd_payload_fragment_address (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[15:0]), //i
    .io_bus_cmd_payload_fragment_length  (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_bus_cmd_payload_fragment_data    (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_bus_cmd_payload_fragment_context (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_bus_rsp_valid                    (system_clint_logic_io_bus_rsp_valid                                                        ), //o
    .io_bus_rsp_ready                    (system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_bus_rsp_payload_last             (system_clint_logic_io_bus_rsp_payload_last                                                 ), //o
    .io_bus_rsp_payload_fragment_opcode  (system_clint_logic_io_bus_rsp_payload_fragment_opcode                                      ), //o
    .io_bus_rsp_payload_fragment_data    (system_clint_logic_io_bus_rsp_payload_fragment_data[31:0]                                  ), //o
    .io_bus_rsp_payload_fragment_context (system_clint_logic_io_bus_rsp_payload_fragment_context[48:0]                               ), //o
    .io_timerInterrupt                   (system_clint_logic_io_timerInterrupt[1:0]                                                  ), //o
    .io_softwareInterrupt                (system_clint_logic_io_softwareInterrupt[1:0]                                               ), //o
    .io_time                             (system_clint_logic_io_time[63:0]                                                           ), //o
    .io_stop                             (system_peripheralStopTime                                                                  ), //i
    .io_peripheralClk                    (io_peripheralClk                                                                           ), //i
    .peripheralCd_logic_outputReset      (peripheralCd_logic_outputReset                                                             )  //i
  );
  BmbUartCtrl system_uart_0_io_logic (
    .io_bus_cmd_valid                    (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_bus_cmd_ready                    (system_uart_0_io_logic_io_bus_cmd_ready                                                                 ), //o
    .io_bus_cmd_payload_last             (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_bus_cmd_payload_fragment_opcode  (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_bus_cmd_payload_fragment_address (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[5:0] ), //i
    .io_bus_cmd_payload_fragment_length  (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_bus_cmd_payload_fragment_data    (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_bus_cmd_payload_fragment_context (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_bus_rsp_valid                    (system_uart_0_io_logic_io_bus_rsp_valid                                                                 ), //o
    .io_bus_rsp_ready                    (_zz_io_bus_rsp_ready_1                                                                                  ), //i
    .io_bus_rsp_payload_last             (system_uart_0_io_logic_io_bus_rsp_payload_last                                                          ), //o
    .io_bus_rsp_payload_fragment_opcode  (system_uart_0_io_logic_io_bus_rsp_payload_fragment_opcode                                               ), //o
    .io_bus_rsp_payload_fragment_data    (system_uart_0_io_logic_io_bus_rsp_payload_fragment_data[31:0]                                           ), //o
    .io_bus_rsp_payload_fragment_context (system_uart_0_io_logic_io_bus_rsp_payload_fragment_context[48:0]                                        ), //o
    .io_uart_txd                         (system_uart_0_io_logic_io_uart_txd                                                                      ), //o
    .io_uart_rxd                         (system_uart_0_io_rxd                                                                                    ), //i
    .io_interrupt                        (system_uart_0_io_logic_io_interrupt                                                                     ), //o
    .io_peripheralClk                    (io_peripheralClk                                                                                        ), //i
    .peripheralCd_logic_outputReset      (peripheralCd_logic_outputReset                                                                          )  //i
  );
  BmbSpiXdrMasterCtrl system_spi_0_io_logic (
    .io_ctrl_cmd_valid                    (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_ctrl_cmd_ready                    (system_spi_0_io_logic_io_ctrl_cmd_ready                                                                ), //o
    .io_ctrl_cmd_payload_last             (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_ctrl_cmd_payload_fragment_address (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[11:0]), //i
    .io_ctrl_cmd_payload_fragment_length  (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_ctrl_cmd_payload_fragment_data    (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_ctrl_cmd_payload_fragment_context (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_ctrl_rsp_valid                    (system_spi_0_io_logic_io_ctrl_rsp_valid                                                                ), //o
    .io_ctrl_rsp_ready                    (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                                  ), //i
    .io_ctrl_rsp_payload_last             (system_spi_0_io_logic_io_ctrl_rsp_payload_last                                                         ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_opcode                                              ), //o
    .io_ctrl_rsp_payload_fragment_data    (system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_data[31:0]                                          ), //o
    .io_ctrl_rsp_payload_fragment_context (system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_context[48:0]                                       ), //o
    .io_spi_sclk_write                    (system_spi_0_io_logic_io_spi_sclk_write                                                                ), //o
    .io_spi_data_0_writeEnable            (system_spi_0_io_logic_io_spi_data_0_writeEnable                                                        ), //o
    .io_spi_data_0_read                   (system_spi_0_io_data_0_read                                                                            ), //i
    .io_spi_data_0_write                  (system_spi_0_io_logic_io_spi_data_0_write                                                              ), //o
    .io_spi_data_1_writeEnable            (system_spi_0_io_logic_io_spi_data_1_writeEnable                                                        ), //o
    .io_spi_data_1_read                   (system_spi_0_io_data_1_read                                                                            ), //i
    .io_spi_data_1_write                  (system_spi_0_io_logic_io_spi_data_1_write                                                              ), //o
    .io_spi_data_2_writeEnable            (system_spi_0_io_logic_io_spi_data_2_writeEnable                                                        ), //o
    .io_spi_data_2_read                   (system_spi_0_io_data_2_read                                                                            ), //i
    .io_spi_data_2_write                  (system_spi_0_io_logic_io_spi_data_2_write                                                              ), //o
    .io_spi_data_3_writeEnable            (system_spi_0_io_logic_io_spi_data_3_writeEnable                                                        ), //o
    .io_spi_data_3_read                   (system_spi_0_io_data_3_read                                                                            ), //i
    .io_spi_data_3_write                  (system_spi_0_io_logic_io_spi_data_3_write                                                              ), //o
    .io_spi_ss                            (system_spi_0_io_logic_io_spi_ss                                                                        ), //o
    .io_interrupt                         (system_spi_0_io_logic_io_interrupt                                                                     ), //o
    .io_peripheralClk                     (io_peripheralClk                                                                                       ), //i
    .peripheralCd_logic_outputReset       (peripheralCd_logic_outputReset                                                                         )  //i
  );
  BmbSpiXdrMasterCtrl system_spi_1_io_logic (
    .io_ctrl_cmd_valid                    (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_ctrl_cmd_ready                    (system_spi_1_io_logic_io_ctrl_cmd_ready                                                                ), //o
    .io_ctrl_cmd_payload_last             (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_ctrl_cmd_payload_fragment_address (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[11:0]), //i
    .io_ctrl_cmd_payload_fragment_length  (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_ctrl_cmd_payload_fragment_data    (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_ctrl_cmd_payload_fragment_context (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_ctrl_rsp_valid                    (system_spi_1_io_logic_io_ctrl_rsp_valid                                                                ), //o
    .io_ctrl_rsp_ready                    (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                                  ), //i
    .io_ctrl_rsp_payload_last             (system_spi_1_io_logic_io_ctrl_rsp_payload_last                                                         ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_opcode                                              ), //o
    .io_ctrl_rsp_payload_fragment_data    (system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_data[31:0]                                          ), //o
    .io_ctrl_rsp_payload_fragment_context (system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_context[48:0]                                       ), //o
    .io_spi_sclk_write                    (system_spi_1_io_logic_io_spi_sclk_write                                                                ), //o
    .io_spi_data_0_writeEnable            (system_spi_1_io_logic_io_spi_data_0_writeEnable                                                        ), //o
    .io_spi_data_0_read                   (system_spi_1_io_data_0_read                                                                            ), //i
    .io_spi_data_0_write                  (system_spi_1_io_logic_io_spi_data_0_write                                                              ), //o
    .io_spi_data_1_writeEnable            (system_spi_1_io_logic_io_spi_data_1_writeEnable                                                        ), //o
    .io_spi_data_1_read                   (system_spi_1_io_data_1_read                                                                            ), //i
    .io_spi_data_1_write                  (system_spi_1_io_logic_io_spi_data_1_write                                                              ), //o
    .io_spi_data_2_writeEnable            (system_spi_1_io_logic_io_spi_data_2_writeEnable                                                        ), //o
    .io_spi_data_2_read                   (system_spi_1_io_data_2_read                                                                            ), //i
    .io_spi_data_2_write                  (system_spi_1_io_logic_io_spi_data_2_write                                                              ), //o
    .io_spi_data_3_writeEnable            (system_spi_1_io_logic_io_spi_data_3_writeEnable                                                        ), //o
    .io_spi_data_3_read                   (system_spi_1_io_data_3_read                                                                            ), //i
    .io_spi_data_3_write                  (system_spi_1_io_logic_io_spi_data_3_write                                                              ), //o
    .io_spi_ss                            (system_spi_1_io_logic_io_spi_ss                                                                        ), //o
    .io_interrupt                         (system_spi_1_io_logic_io_interrupt                                                                     ), //o
    .io_peripheralClk                     (io_peripheralClk                                                                                       ), //i
    .peripheralCd_logic_outputReset       (peripheralCd_logic_outputReset                                                                         )  //i
  );
  BmbI2cCtrl system_i2c_0_io_logic (
    .io_ctrl_cmd_valid                    (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_ctrl_cmd_ready                    (system_i2c_0_io_logic_io_ctrl_cmd_ready                                                                ), //o
    .io_ctrl_cmd_payload_last             (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_ctrl_cmd_payload_fragment_address (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[7:0] ), //i
    .io_ctrl_cmd_payload_fragment_length  (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_ctrl_cmd_payload_fragment_data    (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_ctrl_cmd_payload_fragment_context (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_ctrl_rsp_valid                    (system_i2c_0_io_logic_io_ctrl_rsp_valid                                                                ), //o
    .io_ctrl_rsp_ready                    (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                                  ), //i
    .io_ctrl_rsp_payload_last             (system_i2c_0_io_logic_io_ctrl_rsp_payload_last                                                         ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_opcode                                              ), //o
    .io_ctrl_rsp_payload_fragment_data    (system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_data[31:0]                                          ), //o
    .io_ctrl_rsp_payload_fragment_context (system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_context[48:0]                                       ), //o
    .io_i2c_sda_write                     (system_i2c_0_io_logic_io_i2c_sda_write                                                                 ), //o
    .io_i2c_sda_read                      (system_i2c_0_io_sda_read                                                                               ), //i
    .io_i2c_scl_write                     (system_i2c_0_io_logic_io_i2c_scl_write                                                                 ), //o
    .io_i2c_scl_read                      (system_i2c_0_io_scl_read                                                                               ), //i
    .io_interrupt                         (system_i2c_0_io_logic_io_interrupt                                                                     ), //o
    .io_peripheralClk                     (io_peripheralClk                                                                                       ), //i
    .peripheralCd_logic_outputReset       (peripheralCd_logic_outputReset                                                                         )  //i
  );
  BmbI2cCtrl system_i2c_2_io_logic (
    .io_ctrl_cmd_valid                    (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_ctrl_cmd_ready                    (system_i2c_2_io_logic_io_ctrl_cmd_ready                                                                ), //o
    .io_ctrl_cmd_payload_last             (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_ctrl_cmd_payload_fragment_address (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[7:0] ), //i
    .io_ctrl_cmd_payload_fragment_length  (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_ctrl_cmd_payload_fragment_data    (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_ctrl_cmd_payload_fragment_context (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_ctrl_rsp_valid                    (system_i2c_2_io_logic_io_ctrl_rsp_valid                                                                ), //o
    .io_ctrl_rsp_ready                    (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                                  ), //i
    .io_ctrl_rsp_payload_last             (system_i2c_2_io_logic_io_ctrl_rsp_payload_last                                                         ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_opcode                                              ), //o
    .io_ctrl_rsp_payload_fragment_data    (system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_data[31:0]                                          ), //o
    .io_ctrl_rsp_payload_fragment_context (system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_context[48:0]                                       ), //o
    .io_i2c_sda_write                     (system_i2c_2_io_logic_io_i2c_sda_write                                                                 ), //o
    .io_i2c_sda_read                      (system_i2c_2_io_sda_read                                                                               ), //i
    .io_i2c_scl_write                     (system_i2c_2_io_logic_io_i2c_scl_write                                                                 ), //o
    .io_i2c_scl_read                      (system_i2c_2_io_scl_read                                                                               ), //i
    .io_interrupt                         (system_i2c_2_io_logic_io_interrupt                                                                     ), //o
    .io_peripheralClk                     (io_peripheralClk                                                                                       ), //i
    .peripheralCd_logic_outputReset       (peripheralCd_logic_outputReset                                                                         )  //i
  );
  BmbI2cCtrl system_i2c_1_io_logic (
    .io_ctrl_cmd_valid                    (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_ctrl_cmd_ready                    (system_i2c_1_io_logic_io_ctrl_cmd_ready                                                                ), //o
    .io_ctrl_cmd_payload_last             (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_ctrl_cmd_payload_fragment_address (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[7:0] ), //i
    .io_ctrl_cmd_payload_fragment_length  (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_ctrl_cmd_payload_fragment_data    (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_ctrl_cmd_payload_fragment_context (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_ctrl_rsp_valid                    (system_i2c_1_io_logic_io_ctrl_rsp_valid                                                                ), //o
    .io_ctrl_rsp_ready                    (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                                  ), //i
    .io_ctrl_rsp_payload_last             (system_i2c_1_io_logic_io_ctrl_rsp_payload_last                                                         ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_opcode                                              ), //o
    .io_ctrl_rsp_payload_fragment_data    (system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_data[31:0]                                          ), //o
    .io_ctrl_rsp_payload_fragment_context (system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_context[48:0]                                       ), //o
    .io_i2c_sda_write                     (system_i2c_1_io_logic_io_i2c_sda_write                                                                 ), //o
    .io_i2c_sda_read                      (system_i2c_1_io_sda_read                                                                               ), //i
    .io_i2c_scl_write                     (system_i2c_1_io_logic_io_i2c_scl_write                                                                 ), //o
    .io_i2c_scl_read                      (system_i2c_1_io_scl_read                                                                               ), //i
    .io_interrupt                         (system_i2c_1_io_logic_io_interrupt                                                                     ), //o
    .io_peripheralClk                     (io_peripheralClk                                                                                       ), //i
    .peripheralCd_logic_outputReset       (peripheralCd_logic_outputReset                                                                         )  //i
  );
  EfxTimerCtrl system_userTimer_1_logic (
    .io_ctrl_cmd_valid                    (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_ctrl_cmd_ready                    (system_userTimer_1_logic_io_ctrl_cmd_ready                                                                ), //o
    .io_ctrl_cmd_payload_last             (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_ctrl_cmd_payload_fragment_address (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[7:0] ), //i
    .io_ctrl_cmd_payload_fragment_length  (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_ctrl_cmd_payload_fragment_data    (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_ctrl_cmd_payload_fragment_context (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_ctrl_rsp_valid                    (system_userTimer_1_logic_io_ctrl_rsp_valid                                                                ), //o
    .io_ctrl_rsp_ready                    (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                                  ), //i
    .io_ctrl_rsp_payload_last             (system_userTimer_1_logic_io_ctrl_rsp_payload_last                                                         ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_opcode                                              ), //o
    .io_ctrl_rsp_payload_fragment_data    (system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_data[31:0]                                          ), //o
    .io_ctrl_rsp_payload_fragment_context (system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_context[48:0]                                       ), //o
    .io_interrupts                        (system_userTimer_1_logic_io_interrupts                                                                    ), //o
    .io_peripheralClk                     (io_peripheralClk                                                                                          ), //i
    .peripheralCd_logic_outputReset       (peripheralCd_logic_outputReset                                                                            )  //i
  );
  EfxTimerCtrl system_userTimer_0_logic (
    .io_ctrl_cmd_valid                    (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid                         ), //i
    .io_ctrl_cmd_ready                    (system_userTimer_0_logic_io_ctrl_cmd_ready                                                                ), //o
    .io_ctrl_cmd_payload_last             (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last                  ), //i
    .io_ctrl_cmd_payload_fragment_opcode  (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode       ), //i
    .io_ctrl_cmd_payload_fragment_address (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address[7:0] ), //i
    .io_ctrl_cmd_payload_fragment_length  (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length[1:0]  ), //i
    .io_ctrl_cmd_payload_fragment_data    (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data[31:0]   ), //i
    .io_ctrl_cmd_payload_fragment_context (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context[48:0]), //i
    .io_ctrl_rsp_valid                    (system_userTimer_0_logic_io_ctrl_rsp_valid                                                                ), //o
    .io_ctrl_rsp_ready                    (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                                  ), //i
    .io_ctrl_rsp_payload_last             (system_userTimer_0_logic_io_ctrl_rsp_payload_last                                                         ), //o
    .io_ctrl_rsp_payload_fragment_opcode  (system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_opcode                                              ), //o
    .io_ctrl_rsp_payload_fragment_data    (system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_data[31:0]                                          ), //o
    .io_ctrl_rsp_payload_fragment_context (system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_context[48:0]                                       ), //o
    .io_interrupts                        (system_userTimer_0_logic_io_interrupts                                                                    ), //o
    .io_peripheralClk                     (io_peripheralClk                                                                                          ), //i
    .peripheralCd_logic_outputReset       (peripheralCd_logic_outputReset                                                                            )  //i
  );
  BmbGpio2 system_gpio_0_io_logic (
    .io_gpio_read                        (system_gpio_0_io_read[3:0]                                                                     ), //i
    .io_gpio_write                       (system_gpio_0_io_logic_io_gpio_write[3:0]                                                      ), //o
    .io_gpio_writeEnable                 (system_gpio_0_io_logic_io_gpio_writeEnable[3:0]                                                ), //o
    .io_bus_cmd_valid                    (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_bus_cmd_ready                    (system_gpio_0_io_logic_io_bus_cmd_ready                                                        ), //o
    .io_bus_cmd_payload_last             (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_bus_cmd_payload_fragment_opcode  (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_bus_cmd_payload_fragment_address (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[7:0] ), //i
    .io_bus_cmd_payload_fragment_length  (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_bus_cmd_payload_fragment_data    (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_bus_cmd_payload_fragment_context (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_bus_rsp_valid                    (system_gpio_0_io_logic_io_bus_rsp_valid                                                        ), //o
    .io_bus_rsp_ready                    (system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_bus_rsp_payload_last             (system_gpio_0_io_logic_io_bus_rsp_payload_last                                                 ), //o
    .io_bus_rsp_payload_fragment_opcode  (system_gpio_0_io_logic_io_bus_rsp_payload_fragment_opcode                                      ), //o
    .io_bus_rsp_payload_fragment_data    (system_gpio_0_io_logic_io_bus_rsp_payload_fragment_data[31:0]                                  ), //o
    .io_bus_rsp_payload_fragment_context (system_gpio_0_io_logic_io_bus_rsp_payload_fragment_context[48:0]                               ), //o
    .io_interrupt                        (system_gpio_0_io_logic_io_interrupt[3:0]                                                       ), //o
    .io_peripheralClk                    (io_peripheralClk                                                                               ), //i
    .peripheralCd_logic_outputReset      (peripheralCd_logic_outputReset                                                                 )  //i
  );
  BmbWatchdog system_watchdog_logic_logic (
    .io_bus_cmd_valid                    (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_bus_cmd_ready                    (system_watchdog_logic_logic_io_bus_cmd_ready                                                        ), //o
    .io_bus_cmd_payload_last             (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_bus_cmd_payload_fragment_opcode  (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_bus_cmd_payload_fragment_address (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[7:0] ), //i
    .io_bus_cmd_payload_fragment_length  (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_bus_cmd_payload_fragment_data    (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_bus_cmd_payload_fragment_context (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_bus_rsp_valid                    (system_watchdog_logic_logic_io_bus_rsp_valid                                                        ), //o
    .io_bus_rsp_ready                    (system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_bus_rsp_payload_last             (system_watchdog_logic_logic_io_bus_rsp_payload_last                                                 ), //o
    .io_bus_rsp_payload_fragment_opcode  (system_watchdog_logic_logic_io_bus_rsp_payload_fragment_opcode                                      ), //o
    .io_bus_rsp_payload_fragment_data    (system_watchdog_logic_logic_io_bus_rsp_payload_fragment_data[31:0]                                  ), //o
    .io_bus_rsp_payload_fragment_context (system_watchdog_logic_logic_io_bus_rsp_payload_fragment_context[48:0]                               ), //o
    .io_panics                           (system_watchdog_logic_logic_io_panics[1:0]                                                          ), //o
    .io_heartBeat                        (system_peripheralStopTime                                                                           ), //i
    .io_peripheralClk                    (io_peripheralClk                                                                                    ), //i
    .peripheralCd_logic_outputReset      (peripheralCd_logic_outputReset                                                                      )  //i
  );
  BmbToApb3Bridge io_apbSlave_2_logic (
    .io_input_cmd_valid                    (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_input_cmd_ready                    (io_apbSlave_2_logic_io_input_cmd_ready                                                       ), //o
    .io_input_cmd_payload_last             (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_opcode  (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[15:0]), //i
    .io_input_cmd_payload_fragment_length  (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_input_cmd_payload_fragment_data    (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_input_cmd_payload_fragment_context (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_input_rsp_valid                    (io_apbSlave_2_logic_io_input_rsp_valid                                                       ), //o
    .io_input_rsp_ready                    (io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_input_rsp_payload_last             (io_apbSlave_2_logic_io_input_rsp_payload_last                                                ), //o
    .io_input_rsp_payload_fragment_opcode  (io_apbSlave_2_logic_io_input_rsp_payload_fragment_opcode                                     ), //o
    .io_input_rsp_payload_fragment_data    (io_apbSlave_2_logic_io_input_rsp_payload_fragment_data[31:0]                                 ), //o
    .io_input_rsp_payload_fragment_context (io_apbSlave_2_logic_io_input_rsp_payload_fragment_context[48:0]                              ), //o
    .io_output_PADDR                       (io_apbSlave_2_logic_io_output_PADDR[15:0]                                                    ), //o
    .io_output_PSEL                        (io_apbSlave_2_logic_io_output_PSEL                                                           ), //o
    .io_output_PENABLE                     (io_apbSlave_2_logic_io_output_PENABLE                                                        ), //o
    .io_output_PREADY                      (io_apbSlave_2_PREADY                                                                         ), //i
    .io_output_PWRITE                      (io_apbSlave_2_logic_io_output_PWRITE                                                         ), //o
    .io_output_PWDATA                      (io_apbSlave_2_logic_io_output_PWDATA[31:0]                                                   ), //o
    .io_output_PRDATA                      (io_apbSlave_2_PRDATA[31:0]                                                                   ), //i
    .io_output_PSLVERROR                   (io_apbSlave_2_PSLVERROR                                                                      ), //i
    .io_peripheralClk                      (io_peripheralClk                                                                             ), //i
    .peripheralCd_logic_outputReset        (peripheralCd_logic_outputReset                                                               )  //i
  );
  BmbToApb3Bridge io_apbSlave_1_logic (
    .io_input_cmd_valid                    (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_input_cmd_ready                    (io_apbSlave_1_logic_io_input_cmd_ready                                                       ), //o
    .io_input_cmd_payload_last             (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_opcode  (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[15:0]), //i
    .io_input_cmd_payload_fragment_length  (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_input_cmd_payload_fragment_data    (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_input_cmd_payload_fragment_context (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_input_rsp_valid                    (io_apbSlave_1_logic_io_input_rsp_valid                                                       ), //o
    .io_input_rsp_ready                    (io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_input_rsp_payload_last             (io_apbSlave_1_logic_io_input_rsp_payload_last                                                ), //o
    .io_input_rsp_payload_fragment_opcode  (io_apbSlave_1_logic_io_input_rsp_payload_fragment_opcode                                     ), //o
    .io_input_rsp_payload_fragment_data    (io_apbSlave_1_logic_io_input_rsp_payload_fragment_data[31:0]                                 ), //o
    .io_input_rsp_payload_fragment_context (io_apbSlave_1_logic_io_input_rsp_payload_fragment_context[48:0]                              ), //o
    .io_output_PADDR                       (io_apbSlave_1_logic_io_output_PADDR[15:0]                                                    ), //o
    .io_output_PSEL                        (io_apbSlave_1_logic_io_output_PSEL                                                           ), //o
    .io_output_PENABLE                     (io_apbSlave_1_logic_io_output_PENABLE                                                        ), //o
    .io_output_PREADY                      (io_apbSlave_1_PREADY                                                                         ), //i
    .io_output_PWRITE                      (io_apbSlave_1_logic_io_output_PWRITE                                                         ), //o
    .io_output_PWDATA                      (io_apbSlave_1_logic_io_output_PWDATA[31:0]                                                   ), //o
    .io_output_PRDATA                      (io_apbSlave_1_PRDATA[31:0]                                                                   ), //i
    .io_output_PSLVERROR                   (io_apbSlave_1_PSLVERROR                                                                      ), //i
    .io_peripheralClk                      (io_peripheralClk                                                                             ), //i
    .peripheralCd_logic_outputReset        (peripheralCd_logic_outputReset                                                               )  //i
  );
  BmbToApb3Bridge io_apbSlave_4_logic (
    .io_input_cmd_valid                    (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_input_cmd_ready                    (io_apbSlave_4_logic_io_input_cmd_ready                                                       ), //o
    .io_input_cmd_payload_last             (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_opcode  (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[15:0]), //i
    .io_input_cmd_payload_fragment_length  (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_input_cmd_payload_fragment_data    (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_input_cmd_payload_fragment_context (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_input_rsp_valid                    (io_apbSlave_4_logic_io_input_rsp_valid                                                       ), //o
    .io_input_rsp_ready                    (io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_input_rsp_payload_last             (io_apbSlave_4_logic_io_input_rsp_payload_last                                                ), //o
    .io_input_rsp_payload_fragment_opcode  (io_apbSlave_4_logic_io_input_rsp_payload_fragment_opcode                                     ), //o
    .io_input_rsp_payload_fragment_data    (io_apbSlave_4_logic_io_input_rsp_payload_fragment_data[31:0]                                 ), //o
    .io_input_rsp_payload_fragment_context (io_apbSlave_4_logic_io_input_rsp_payload_fragment_context[48:0]                              ), //o
    .io_output_PADDR                       (io_apbSlave_4_logic_io_output_PADDR[15:0]                                                    ), //o
    .io_output_PSEL                        (io_apbSlave_4_logic_io_output_PSEL                                                           ), //o
    .io_output_PENABLE                     (io_apbSlave_4_logic_io_output_PENABLE                                                        ), //o
    .io_output_PREADY                      (io_apbSlave_4_PREADY                                                                         ), //i
    .io_output_PWRITE                      (io_apbSlave_4_logic_io_output_PWRITE                                                         ), //o
    .io_output_PWDATA                      (io_apbSlave_4_logic_io_output_PWDATA[31:0]                                                   ), //o
    .io_output_PRDATA                      (io_apbSlave_4_PRDATA[31:0]                                                                   ), //i
    .io_output_PSLVERROR                   (io_apbSlave_4_PSLVERROR                                                                      ), //i
    .io_peripheralClk                      (io_peripheralClk                                                                             ), //i
    .peripheralCd_logic_outputReset        (peripheralCd_logic_outputReset                                                               )  //i
  );
  BmbToApb3Bridge io_apbSlave_0_logic (
    .io_input_cmd_valid                    (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_input_cmd_ready                    (io_apbSlave_0_logic_io_input_cmd_ready                                                       ), //o
    .io_input_cmd_payload_last             (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_opcode  (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[15:0]), //i
    .io_input_cmd_payload_fragment_length  (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_input_cmd_payload_fragment_data    (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_input_cmd_payload_fragment_context (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_input_rsp_valid                    (io_apbSlave_0_logic_io_input_rsp_valid                                                       ), //o
    .io_input_rsp_ready                    (io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_input_rsp_payload_last             (io_apbSlave_0_logic_io_input_rsp_payload_last                                                ), //o
    .io_input_rsp_payload_fragment_opcode  (io_apbSlave_0_logic_io_input_rsp_payload_fragment_opcode                                     ), //o
    .io_input_rsp_payload_fragment_data    (io_apbSlave_0_logic_io_input_rsp_payload_fragment_data[31:0]                                 ), //o
    .io_input_rsp_payload_fragment_context (io_apbSlave_0_logic_io_input_rsp_payload_fragment_context[48:0]                              ), //o
    .io_output_PADDR                       (io_apbSlave_0_logic_io_output_PADDR[15:0]                                                    ), //o
    .io_output_PSEL                        (io_apbSlave_0_logic_io_output_PSEL                                                           ), //o
    .io_output_PENABLE                     (io_apbSlave_0_logic_io_output_PENABLE                                                        ), //o
    .io_output_PREADY                      (io_apbSlave_0_PREADY                                                                         ), //i
    .io_output_PWRITE                      (io_apbSlave_0_logic_io_output_PWRITE                                                         ), //o
    .io_output_PWDATA                      (io_apbSlave_0_logic_io_output_PWDATA[31:0]                                                   ), //o
    .io_output_PRDATA                      (io_apbSlave_0_PRDATA[31:0]                                                                   ), //i
    .io_output_PSLVERROR                   (io_apbSlave_0_PSLVERROR                                                                      ), //i
    .io_peripheralClk                      (io_peripheralClk                                                                             ), //i
    .peripheralCd_logic_outputReset        (peripheralCd_logic_outputReset                                                               )  //i
  );
  BmbToApb3Bridge io_apbSlave_3_logic (
    .io_input_cmd_valid                    (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid                         ), //i
    .io_input_cmd_ready                    (io_apbSlave_3_logic_io_input_cmd_ready                                                       ), //o
    .io_input_cmd_payload_last             (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last                  ), //i
    .io_input_cmd_payload_fragment_opcode  (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode       ), //i
    .io_input_cmd_payload_fragment_address (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address[15:0]), //i
    .io_input_cmd_payload_fragment_length  (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length[1:0]  ), //i
    .io_input_cmd_payload_fragment_data    (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data[31:0]   ), //i
    .io_input_cmd_payload_fragment_context (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context[48:0]), //i
    .io_input_rsp_valid                    (io_apbSlave_3_logic_io_input_rsp_valid                                                       ), //o
    .io_input_rsp_ready                    (io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready                         ), //i
    .io_input_rsp_payload_last             (io_apbSlave_3_logic_io_input_rsp_payload_last                                                ), //o
    .io_input_rsp_payload_fragment_opcode  (io_apbSlave_3_logic_io_input_rsp_payload_fragment_opcode                                     ), //o
    .io_input_rsp_payload_fragment_data    (io_apbSlave_3_logic_io_input_rsp_payload_fragment_data[31:0]                                 ), //o
    .io_input_rsp_payload_fragment_context (io_apbSlave_3_logic_io_input_rsp_payload_fragment_context[48:0]                              ), //o
    .io_output_PADDR                       (io_apbSlave_3_logic_io_output_PADDR[15:0]                                                    ), //o
    .io_output_PSEL                        (io_apbSlave_3_logic_io_output_PSEL                                                           ), //o
    .io_output_PENABLE                     (io_apbSlave_3_logic_io_output_PENABLE                                                        ), //o
    .io_output_PREADY                      (io_apbSlave_3_PREADY                                                                         ), //i
    .io_output_PWRITE                      (io_apbSlave_3_logic_io_output_PWRITE                                                         ), //o
    .io_output_PWDATA                      (io_apbSlave_3_logic_io_output_PWDATA[31:0]                                                   ), //o
    .io_output_PRDATA                      (io_apbSlave_3_PRDATA[31:0]                                                                   ), //i
    .io_output_PSLVERROR                   (io_apbSlave_3_PSLVERROR                                                                      ), //i
    .io_peripheralClk                      (io_peripheralClk                                                                             ), //i
    .peripheralCd_logic_outputReset        (peripheralCd_logic_outputReset                                                               )  //i
  );
  StreamCCByToggle_2 io_time_sync_cc (
    .io_input_valid                                                                      (1'b1                                                                                                            ), //i
    .io_input_ready                                                                      (io_time_sync_cc_io_input_ready                                                                                  ), //o
    .io_input_payload                                                                    (system_clint_logic_io_time[63:0]                                                                                ), //i
    .io_output_valid                                                                     (io_time_sync_cc_io_output_valid                                                                                 ), //o
    .io_output_ready                                                                     (1'b1                                                                                                            ), //i
    .io_output_payload                                                                   (io_time_sync_cc_io_output_payload[63:0]                                                                         ), //o
    .io_peripheralClk                                                                    (io_peripheralClk                                                                                                ), //i
    .peripheralCd_logic_outputReset                                                      (peripheralCd_logic_outputReset                                                                                  ), //i
    .io_systemClk                                                                        (io_systemClk                                                                                                    ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //i
  );
  StreamCCByToggle_2 io_time_sync_cc_1 (
    .io_input_valid                                                                      (1'b1                                                                                                            ), //i
    .io_input_ready                                                                      (io_time_sync_cc_1_io_input_ready                                                                                ), //o
    .io_input_payload                                                                    (system_clint_logic_io_time[63:0]                                                                                ), //i
    .io_output_valid                                                                     (io_time_sync_cc_1_io_output_valid                                                                               ), //o
    .io_output_ready                                                                     (1'b1                                                                                                            ), //i
    .io_output_payload                                                                   (io_time_sync_cc_1_io_output_payload[63:0]                                                                       ), //o
    .io_peripheralClk                                                                    (io_peripheralClk                                                                                                ), //i
    .peripheralCd_logic_outputReset                                                      (peripheralCd_logic_outputReset                                                                                  ), //i
    .io_systemClk                                                                        (io_systemClk                                                                                                    ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC bufferCC_74 (
    .io_dataIn                  (bufferCC_74_io_dataIn     ), //i
    .io_dataOut                 (bufferCC_74_io_dataOut    ), //o
    .io_systemClk               (io_systemClk              ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset)  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC bufferCC_75 (
    .io_dataIn                  (bufferCC_75_io_dataIn     ), //i
    .io_dataOut                 (bufferCC_75_io_dataOut    ), //o
    .io_systemClk               (io_systemClk              ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset)  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC bufferCC_76 (
    .io_dataIn                  (bufferCC_76_io_dataIn     ), //i
    .io_dataOut                 (bufferCC_76_io_dataOut    ), //o
    .io_systemClk               (io_systemClk              ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset)  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC bufferCC_77 (
    .io_dataIn                  (bufferCC_77_io_dataIn     ), //i
    .io_dataOut                 (bufferCC_77_io_dataOut    ), //o
    .io_systemClk               (io_systemClk              ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset)  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC system_cores_0_externalInterrupt_plic_target_iep_regNext_buffercc (
    .io_dataIn                  (system_cores_0_externalInterrupt_plic_target_iep_regNext                    ), //i
    .io_dataOut                 (system_cores_0_externalInterrupt_plic_target_iep_regNext_buffercc_io_dataOut), //o
    .io_systemClk               (io_systemClk                                                                ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                                                  )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC system_cores_1_externalInterrupt_plic_target_iep_regNext_buffercc (
    .io_dataIn                  (system_cores_1_externalInterrupt_plic_target_iep_regNext                    ), //i
    .io_dataOut                 (system_cores_1_externalInterrupt_plic_target_iep_regNext_buffercc_io_dataOut), //o
    .io_systemClk               (io_systemClk                                                                ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                                                  )  //i
  );
  initial begin
    debugCd_logic_holdingLogic_resetCounter = 12'h0;
    debugCd_logic_outputReset = 1'b1;
    system_ddr_ddrLogic_ddrAReset_counter = 5'h0;
    system_ddr_ddrLogic_ddrAReset_reset = 1'b1;
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(system_cores_0_debugRiscv_dmToHart_payload_op)
      DebugDmToHartOp_DATA : system_cores_0_debugRiscv_dmToHart_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : system_cores_0_debugRiscv_dmToHart_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : system_cores_0_debugRiscv_dmToHart_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : system_cores_0_debugRiscv_dmToHart_payload_op_string = "REG_READ ";
      default : system_cores_0_debugRiscv_dmToHart_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(system_cores_1_debugRiscv_dmToHart_payload_op)
      DebugDmToHartOp_DATA : system_cores_1_debugRiscv_dmToHart_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : system_cores_1_debugRiscv_dmToHart_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : system_cores_1_debugRiscv_dmToHart_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : system_cores_1_debugRiscv_dmToHart_payload_op_string = "REG_READ ";
      default : system_cores_1_debugRiscv_dmToHart_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_commit_m2sPipe_payload_opcode)
      FpuOpcode_LOAD : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "FCVT_X_X";
      default : FpuPlugin_port_commit_m2sPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_commit_rData_opcode)
      FpuOpcode_LOAD : FpuPlugin_port_commit_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_commit_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_commit_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_commit_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_commit_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_commit_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_commit_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_commit_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_commit_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_commit_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_commit_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_commit_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_commit_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_commit_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_commit_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_commit_rData_opcode_string = "FCVT_X_X";
      default : FpuPlugin_port_commit_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_commit_m2sPipe_payload_opcode_1)
      FpuOpcode_LOAD : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "FCVT_X_X";
      default : FpuPlugin_port_commit_m2sPipe_payload_opcode_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_commit_rData_opcode_1)
      FpuOpcode_LOAD : FpuPlugin_port_commit_rData_opcode_1_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_commit_rData_opcode_1_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_commit_rData_opcode_1_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_commit_rData_opcode_1_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_commit_rData_opcode_1_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_commit_rData_opcode_1_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_commit_rData_opcode_1_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_commit_rData_opcode_1_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_commit_rData_opcode_1_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_commit_rData_opcode_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_commit_rData_opcode_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_commit_rData_opcode_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_commit_rData_opcode_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_commit_rData_opcode_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_commit_rData_opcode_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_commit_rData_opcode_1_string = "FCVT_X_X";
      default : FpuPlugin_port_commit_rData_opcode_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_harts_0_dmToHart_regNext_payload_op)
      DebugDmToHartOp_DATA : io_harts_0_dmToHart_regNext_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : io_harts_0_dmToHart_regNext_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : io_harts_0_dmToHart_regNext_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : io_harts_0_dmToHart_regNext_payload_op_string = "REG_READ ";
      default : io_harts_0_dmToHart_regNext_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_harts_1_dmToHart_regNext_payload_op)
      DebugDmToHartOp_DATA : io_harts_1_dmToHart_regNext_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : io_harts_1_dmToHart_regNext_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : io_harts_1_dmToHart_regNext_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : io_harts_1_dmToHart_regNext_payload_op_string = "REG_READ ";
      default : io_harts_1_dmToHart_regNext_payload_op_string = "?????????";
    endcase
  end
  `endif

  always @(*) begin
    debugCd_logic_inputResetTrigger = 1'b0;
    if(debugCd_logic_inputResetAdapter_stuff_syncTrigger) begin
      debugCd_logic_inputResetTrigger = 1'b1;
    end
  end

  always @(*) begin
    debugCd_logic_outputResetUnbuffered = 1'b0;
    if(when_ClockDomainGenerator_l222) begin
      debugCd_logic_outputResetUnbuffered = 1'b1;
    end
  end

  assign when_ClockDomainGenerator_l222 = (debugCd_logic_holdingLogic_resetCounter != 12'hfff);
  always @(*) begin
    ddrCd_logic_inputResetTrigger = 1'b0;
    if(debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut) begin
      ddrCd_logic_inputResetTrigger = 1'b1;
    end
    if(system_riscvJtag_debug_systemReset_asyncAssertSyncDeassert_buffercc_io_dataOut) begin
      ddrCd_logic_inputResetTrigger = 1'b1;
    end
  end

  always @(*) begin
    ddrCd_logic_outputResetUnbuffered = 1'b0;
    if(when_ClockDomainGenerator_l222_1) begin
      ddrCd_logic_outputResetUnbuffered = 1'b1;
    end
  end

  assign when_ClockDomainGenerator_l222_1 = (ddrCd_logic_holdingLogic_resetCounter != 6'h3f);
  always @(*) begin
    peripheralCd_logic_inputResetTrigger = 1'b0;
    if(ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut) begin
      peripheralCd_logic_inputResetTrigger = 1'b1;
    end
  end

  always @(*) begin
    peripheralCd_logic_outputResetUnbuffered = 1'b0;
    if(when_ClockDomainGenerator_l222_2) begin
      peripheralCd_logic_outputResetUnbuffered = 1'b1;
    end
  end

  assign when_ClockDomainGenerator_l222_2 = (peripheralCd_logic_holdingLogic_resetCounter != 6'h3f);
  assign io_asyncReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign debugCd_logic_inputResetAdapter_stuff_syncTrigger = io_asyncReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign debugCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  always @(*) begin
    systemCd_logic_inputResetTrigger = 1'b0;
    if(peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut) begin
      systemCd_logic_inputResetTrigger = 1'b1;
    end
  end

  always @(*) begin
    systemCd_logic_outputResetUnbuffered = 1'b0;
    if(when_ClockDomainGenerator_l222_3) begin
      systemCd_logic_outputResetUnbuffered = 1'b1;
    end
  end

  assign when_ClockDomainGenerator_l222_3 = (systemCd_logic_holdingLogic_resetCounter != 6'h3f);
  assign peripheralCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign ddrCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign userInterruptA_interrupt = userInterruptA_buffercc_io_dataOut;
  assign userInterruptD_interrupt = userInterruptD_buffercc_io_dataOut;
  assign userInterruptC_interrupt = userInterruptC_buffercc_io_dataOut;
  assign userInterruptB_interrupt = userInterruptB_buffercc_io_dataOut;
  assign when_PlicGateway_l21 = (! userInterruptA_interrupt_plic_gateway_waitCompletion);
  assign when_PlicGateway_l21_1 = (! userInterruptD_interrupt_plic_gateway_waitCompletion);
  assign when_PlicGateway_l21_2 = (! userInterruptC_interrupt_plic_gateway_waitCompletion);
  assign when_PlicGateway_l21_3 = (! userInterruptB_interrupt_plic_gateway_waitCompletion);
  always @(*) begin
    system_coreStopTime = 1'b0;
    if(_zz_1) begin
      system_coreStopTime = 1'b1;
    end
  end

  assign system_cores_0_iBus_cmd_valid = system_cores_0_logic_cpu_iBus_cmd_valid;
  assign system_cores_0_iBus_cmd_payload_fragment_opcode = 1'b0;
  assign system_cores_0_iBus_cmd_payload_fragment_address = system_cores_0_logic_cpu_iBus_cmd_payload_address;
  assign system_cores_0_iBus_cmd_payload_fragment_length = 6'h3f;
  assign system_cores_0_iBus_cmd_payload_last = 1'b1;
  assign system_cores_0_logic_cpu_iBus_rsp_payload_error = (system_cores_0_iBus_rsp_payload_fragment_opcode == 1'b1);
  assign system_cores_0_iBus_rsp_ready = 1'b1;
  always @(*) begin
    _zz_dBus_cmd_ready = dBus_Bridge_withWriteBuffer_buffer_stream_ready;
    if(when_Stream_l375) begin
      _zz_dBus_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! dBus_Bridge_withWriteBuffer_buffer_stream_valid);
  assign dBus_Bridge_withWriteBuffer_buffer_stream_valid = _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid;
  assign dBus_Bridge_withWriteBuffer_aggregationCounterFull = (dBus_Bridge_withWriteBuffer_aggregationCounter == 4'b1111);
  assign dBus_Bridge_withWriteBuffer_timerFull = dBus_Bridge_withWriteBuffer_timer[5];
  assign dBus_Bridge_withWriteBuffer_hit = (system_cores_0_logic_cpu_dBus_cmd_payload_address[31 : 3] == dBus_Bridge_withWriteBuffer_buffer_address[31 : 3]);
  assign dBus_Bridge_withWriteBuffer_canAggregate = ((((((system_cores_0_logic_cpu_dBus_cmd_valid && system_cores_0_logic_cpu_dBus_cmd_payload_wr) && (! system_cores_0_logic_cpu_dBus_cmd_payload_uncached)) && (! system_cores_0_logic_cpu_dBus_cmd_payload_exclusive)) && (! dBus_Bridge_withWriteBuffer_timerFull)) && (! dBus_Bridge_withWriteBuffer_aggregationCounterFull)) && ((! dBus_Bridge_withWriteBuffer_buffer_stream_valid) || (dBus_Bridge_withWriteBuffer_aggregationEnabled && dBus_Bridge_withWriteBuffer_hit)));
  assign dBus_Bridge_withWriteBuffer_doFlush = ((((system_cores_0_logic_cpu_dBus_cmd_valid && (! dBus_Bridge_withWriteBuffer_canAggregate)) || dBus_Bridge_withWriteBuffer_timerFull) || dBus_Bridge_withWriteBuffer_aggregationCounterFull) || (! dBus_Bridge_withWriteBuffer_aggregationEnabled));
  always @(*) begin
    dBus_Bridge_withWriteBuffer_halt = 1'b0;
    if(when_DataCache_l523) begin
      dBus_Bridge_withWriteBuffer_halt = 1'b1;
    end
  end

  assign dBus_cmd_fire = (system_cores_0_logic_cpu_dBus_cmd_valid && _zz_dBus_cmd_ready);
  assign when_DataCache_l465 = (dBus_Bridge_withWriteBuffer_buffer_stream_valid && (! dBus_Bridge_withWriteBuffer_timerFull));
  assign dBus_Bridge_bus_cmd_fire = (dBus_Bridge_bus_cmd_valid && dBus_Bridge_bus_cmd_ready);
  assign when_DataCache_l468 = (dBus_Bridge_bus_cmd_fire || (! dBus_Bridge_withWriteBuffer_buffer_stream_valid));
  assign dBus_Bridge_withWriteBuffer_buffer_stream_ready = (((dBus_Bridge_bus_cmd_ready && dBus_Bridge_withWriteBuffer_doFlush) || dBus_Bridge_withWriteBuffer_canAggregate) && (! dBus_Bridge_withWriteBuffer_halt));
  assign dBus_Bridge_bus_cmd_valid = ((dBus_Bridge_withWriteBuffer_buffer_stream_valid && dBus_Bridge_withWriteBuffer_doFlush) && (! dBus_Bridge_withWriteBuffer_halt));
  assign dBus_Bridge_bus_cmd_payload_last = 1'b1;
  assign dBus_Bridge_bus_cmd_payload_fragment_opcode = (dBus_Bridge_withWriteBuffer_buffer_write ? 1'b1 : 1'b0);
  assign dBus_Bridge_bus_cmd_payload_fragment_address = dBus_Bridge_withWriteBuffer_buffer_address;
  assign dBus_Bridge_bus_cmd_payload_fragment_length = dBus_Bridge_withWriteBuffer_buffer_length;
  assign dBus_Bridge_bus_cmd_payload_fragment_data = dBus_Bridge_withWriteBuffer_buffer_data;
  assign dBus_Bridge_bus_cmd_payload_fragment_mask = dBus_Bridge_withWriteBuffer_buffer_mask;
  assign dBus_Bridge_bus_cmd_payload_fragment_exclusive = dBus_Bridge_withWriteBuffer_buffer_exclusive;
  assign dBus_Bridge_bus_cmd_payload_fragment_context = dBus_Bridge_withWriteBuffer_busCmdContext_rspCount;
  assign dBus_Bridge_withWriteBuffer_busCmdContext_rspCount = dBus_Bridge_withWriteBuffer_aggregationCounter;
  assign when_DataCache_l493 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[0]);
  assign when_DataCache_l493_1 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[1]);
  assign when_DataCache_l493_2 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[2]);
  assign when_DataCache_l493_3 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[3]);
  assign when_DataCache_l493_4 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[4]);
  assign when_DataCache_l493_5 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[5]);
  assign when_DataCache_l493_6 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[6]);
  assign when_DataCache_l493_7 = (1'b1 && system_cores_0_logic_cpu_dBus_cmd_payload_mask[7]);
  always @(*) begin
    _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'bxxxxxx;
    case(system_cores_0_logic_cpu_dBus_cmd_payload_size)
      3'b000 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'h0;
      end
      3'b001 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'h01;
      end
      3'b010 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'h03;
      end
      3'b011 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'h07;
      end
      3'b100 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'h0f;
      end
      3'b101 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'h1f;
      end
      3'b110 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length = 6'h3f;
      end
      default : begin
      end
    endcase
  end

  assign when_DataCache_l506 = ((system_cores_0_logic_cpu_dBus_cmd_payload_wr && (! system_cores_0_logic_cpu_dBus_cmd_payload_uncached)) && (! system_cores_0_logic_cpu_dBus_cmd_payload_exclusive));
  assign dBus_Bridge_withWriteBuffer_rspCtx_rspCount = dBus_Bridge_bus_rsp_payload_fragment_context[3 : 0];
  assign dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_valid = (dBus_Bridge_bus_cmd_fire && (dBus_Bridge_bus_cmd_payload_fragment_opcode == 1'b1));
  assign dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_payload = dBus_Bridge_withWriteBuffer_aggregationCounter;
  assign when_DataCache_l523 = (! dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_ready);
  assign dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_ready = dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_push_ready;
  assign io_pop_s2mPipe_valid = (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_valid || (! io_pop_rValidN));
  assign io_pop_s2mPipe_payload = (io_pop_rValidN ? dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_payload : io_pop_rData);
  always @(*) begin
    io_pop_s2mPipe_ready = dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_ready;
    if(when_Stream_l375_1) begin
      io_pop_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_valid);
  assign dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_valid = io_pop_s2mPipe_rValid;
  assign dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_payload = io_pop_s2mPipe_rData;
  assign dBus_Bridge_bus_sync_fire = (dBus_Bridge_bus_sync_valid && dBus_Bridge_bus_sync_ready);
  assign dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_ready = dBus_Bridge_bus_sync_fire;
  assign dBus_Bridge_bus_sync_ready = system_cores_0_logic_cpu_dBus_sync_ready;
  assign system_cores_0_logic_cpu_dBus_rsp_payload_error = (dBus_Bridge_bus_rsp_payload_fragment_opcode == 1'b1);
  assign dBus_Bridge_bus_rsp_ready = 1'b1;
  assign system_cores_0_logic_cpu_dBus_inv_payload_fragment_address = (dBus_Bridge_bus_inv_payload_address + _zz_dBus_inv_payload_fragment_address);
  assign system_cores_0_logic_cpu_dBus_inv_payload_last = 1'b1;
  assign dBus_Bridge_bus_inv_ready = (system_cores_0_logic_cpu_dBus_inv_payload_last && system_cores_0_logic_cpu_dBus_inv_ready);
  assign when_Stream_l445 = (! system_cores_0_logic_cpu_dBus_ack_payload_last);
  always @(*) begin
    dBus_ack_thrown_valid = system_cores_0_logic_cpu_dBus_ack_valid;
    if(when_Stream_l445) begin
      dBus_ack_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    system_cores_0_logic_cpu_dBus_ack_ready = dBus_ack_thrown_ready;
    if(when_Stream_l445) begin
      system_cores_0_logic_cpu_dBus_ack_ready = 1'b1;
    end
  end

  assign dBus_ack_thrown_payload_last = system_cores_0_logic_cpu_dBus_ack_payload_last;
  assign dBus_ack_thrown_payload_fragment_hit = system_cores_0_logic_cpu_dBus_ack_payload_fragment_hit;
  assign dBus_Bridge_bus_ack_valid = dBus_ack_thrown_valid;
  assign dBus_ack_thrown_ready = dBus_Bridge_bus_ack_ready;
  assign system_cores_0_debugRiscv_halted = system_cores_0_logic_cpu_debugBus_halted;
  assign system_cores_0_debugRiscv_running = system_cores_0_logic_cpu_debugBus_running;
  assign system_cores_0_debugRiscv_unavailable = system_cores_0_logic_cpu_debugBus_unavailable;
  assign system_cores_0_debugRiscv_exception = system_cores_0_logic_cpu_debugBus_exception;
  assign system_cores_0_debugRiscv_commit = system_cores_0_logic_cpu_debugBus_commit;
  assign system_cores_0_debugRiscv_ebreak = system_cores_0_logic_cpu_debugBus_ebreak;
  assign system_cores_0_debugRiscv_redo = system_cores_0_logic_cpu_debugBus_redo;
  assign system_cores_0_debugRiscv_regSuccess = system_cores_0_logic_cpu_debugBus_regSuccess;
  assign system_cores_0_debugRiscv_haveReset = system_cores_0_logic_cpu_debugBus_haveReset;
  assign system_cores_0_debugRiscv_resume_rsp_valid = system_cores_0_logic_cpu_debugBus_resume_rsp_valid;
  assign system_cores_0_debugRiscv_hartToDm_valid = system_cores_0_logic_cpu_debugBus_hartToDm_valid;
  assign system_cores_0_debugRiscv_hartToDm_payload_address = system_cores_0_logic_cpu_debugBus_hartToDm_payload_address;
  assign system_cores_0_debugRiscv_hartToDm_payload_data = system_cores_0_logic_cpu_debugBus_hartToDm_payload_data;
  assign system_cores_1_iBus_cmd_valid = system_cores_1_logic_cpu_iBus_cmd_valid;
  assign system_cores_1_iBus_cmd_payload_fragment_opcode = 1'b0;
  assign system_cores_1_iBus_cmd_payload_fragment_address = system_cores_1_logic_cpu_iBus_cmd_payload_address;
  assign system_cores_1_iBus_cmd_payload_fragment_length = 6'h3f;
  assign system_cores_1_iBus_cmd_payload_last = 1'b1;
  assign system_cores_1_logic_cpu_iBus_rsp_payload_error = (system_cores_1_iBus_rsp_payload_fragment_opcode == 1'b1);
  assign system_cores_1_iBus_rsp_ready = 1'b1;
  always @(*) begin
    _zz_dBus_cmd_ready_1 = dBus_Bridge_withWriteBuffer_buffer_stream_ready_1;
    if(when_Stream_l375_2) begin
      _zz_dBus_cmd_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_2 = (! dBus_Bridge_withWriteBuffer_buffer_stream_valid_1);
  assign dBus_Bridge_withWriteBuffer_buffer_stream_valid_1 = _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid_1;
  assign dBus_Bridge_withWriteBuffer_aggregationCounterFull_1 = (dBus_Bridge_withWriteBuffer_aggregationCounter_1 == 4'b1111);
  assign dBus_Bridge_withWriteBuffer_timerFull_1 = dBus_Bridge_withWriteBuffer_timer_1[5];
  assign dBus_Bridge_withWriteBuffer_hit_1 = (system_cores_1_logic_cpu_dBus_cmd_payload_address[31 : 3] == dBus_Bridge_withWriteBuffer_buffer_address_1[31 : 3]);
  assign dBus_Bridge_withWriteBuffer_canAggregate_1 = ((((((system_cores_1_logic_cpu_dBus_cmd_valid && system_cores_1_logic_cpu_dBus_cmd_payload_wr) && (! system_cores_1_logic_cpu_dBus_cmd_payload_uncached)) && (! system_cores_1_logic_cpu_dBus_cmd_payload_exclusive)) && (! dBus_Bridge_withWriteBuffer_timerFull_1)) && (! dBus_Bridge_withWriteBuffer_aggregationCounterFull_1)) && ((! dBus_Bridge_withWriteBuffer_buffer_stream_valid_1) || (dBus_Bridge_withWriteBuffer_aggregationEnabled_1 && dBus_Bridge_withWriteBuffer_hit_1)));
  assign dBus_Bridge_withWriteBuffer_doFlush_1 = ((((system_cores_1_logic_cpu_dBus_cmd_valid && (! dBus_Bridge_withWriteBuffer_canAggregate_1)) || dBus_Bridge_withWriteBuffer_timerFull_1) || dBus_Bridge_withWriteBuffer_aggregationCounterFull_1) || (! dBus_Bridge_withWriteBuffer_aggregationEnabled_1));
  always @(*) begin
    dBus_Bridge_withWriteBuffer_halt_1 = 1'b0;
    if(when_DataCache_l523_1) begin
      dBus_Bridge_withWriteBuffer_halt_1 = 1'b1;
    end
  end

  assign dBus_cmd_fire_1 = (system_cores_1_logic_cpu_dBus_cmd_valid && _zz_dBus_cmd_ready_1);
  assign when_DataCache_l465_1 = (dBus_Bridge_withWriteBuffer_buffer_stream_valid_1 && (! dBus_Bridge_withWriteBuffer_timerFull_1));
  assign dBus_Bridge_bus_cmd_fire_1 = (dBus_Bridge_bus_cmd_valid_1 && dBus_Bridge_bus_cmd_ready_1);
  assign when_DataCache_l468_1 = (dBus_Bridge_bus_cmd_fire_1 || (! dBus_Bridge_withWriteBuffer_buffer_stream_valid_1));
  assign dBus_Bridge_withWriteBuffer_buffer_stream_ready_1 = (((dBus_Bridge_bus_cmd_ready_1 && dBus_Bridge_withWriteBuffer_doFlush_1) || dBus_Bridge_withWriteBuffer_canAggregate_1) && (! dBus_Bridge_withWriteBuffer_halt_1));
  assign dBus_Bridge_bus_cmd_valid_1 = ((dBus_Bridge_withWriteBuffer_buffer_stream_valid_1 && dBus_Bridge_withWriteBuffer_doFlush_1) && (! dBus_Bridge_withWriteBuffer_halt_1));
  assign dBus_Bridge_bus_cmd_payload_last_1 = 1'b1;
  assign dBus_Bridge_bus_cmd_payload_fragment_opcode_1 = (dBus_Bridge_withWriteBuffer_buffer_write_1 ? 1'b1 : 1'b0);
  assign dBus_Bridge_bus_cmd_payload_fragment_address_1 = dBus_Bridge_withWriteBuffer_buffer_address_1;
  assign dBus_Bridge_bus_cmd_payload_fragment_length_1 = dBus_Bridge_withWriteBuffer_buffer_length_1;
  assign dBus_Bridge_bus_cmd_payload_fragment_data_1 = dBus_Bridge_withWriteBuffer_buffer_data_1;
  assign dBus_Bridge_bus_cmd_payload_fragment_mask_1 = dBus_Bridge_withWriteBuffer_buffer_mask_1;
  assign dBus_Bridge_bus_cmd_payload_fragment_exclusive_1 = dBus_Bridge_withWriteBuffer_buffer_exclusive_1;
  assign dBus_Bridge_bus_cmd_payload_fragment_context_1 = dBus_Bridge_withWriteBuffer_busCmdContext_rspCount_1;
  assign dBus_Bridge_withWriteBuffer_busCmdContext_rspCount_1 = dBus_Bridge_withWriteBuffer_aggregationCounter_1;
  assign when_DataCache_l493_8 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[0]);
  assign when_DataCache_l493_9 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[1]);
  assign when_DataCache_l493_10 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[2]);
  assign when_DataCache_l493_11 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[3]);
  assign when_DataCache_l493_12 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[4]);
  assign when_DataCache_l493_13 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[5]);
  assign when_DataCache_l493_14 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[6]);
  assign when_DataCache_l493_15 = (1'b1 && system_cores_1_logic_cpu_dBus_cmd_payload_mask[7]);
  always @(*) begin
    _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'bxxxxxx;
    case(system_cores_1_logic_cpu_dBus_cmd_payload_size)
      3'b000 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'h0;
      end
      3'b001 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'h01;
      end
      3'b010 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'h03;
      end
      3'b011 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'h07;
      end
      3'b100 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'h0f;
      end
      3'b101 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'h1f;
      end
      3'b110 : begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_length_1 = 6'h3f;
      end
      default : begin
      end
    endcase
  end

  assign when_DataCache_l506_1 = ((system_cores_1_logic_cpu_dBus_cmd_payload_wr && (! system_cores_1_logic_cpu_dBus_cmd_payload_uncached)) && (! system_cores_1_logic_cpu_dBus_cmd_payload_exclusive));
  assign dBus_Bridge_withWriteBuffer_rspCtx_rspCount_1 = dBus_Bridge_bus_rsp_payload_fragment_context_1[3 : 0];
  assign dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_valid_1 = (dBus_Bridge_bus_cmd_fire_1 && (dBus_Bridge_bus_cmd_payload_fragment_opcode_1 == 1'b1));
  assign dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_payload_1 = dBus_Bridge_withWriteBuffer_aggregationCounter_1;
  assign when_DataCache_l523_1 = (! dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_ready_1);
  assign dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_ready_1 = dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_push_ready;
  assign io_pop_s2mPipe_valid_1 = (dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_valid || (! io_pop_rValidN_1));
  assign io_pop_s2mPipe_payload_1 = (io_pop_rValidN_1 ? dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_payload : io_pop_rData_1);
  always @(*) begin
    io_pop_s2mPipe_ready_1 = dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_ready_1;
    if(when_Stream_l375_3) begin
      io_pop_s2mPipe_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_3 = (! dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_valid_1);
  assign dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_valid_1 = io_pop_s2mPipe_rValid_1;
  assign dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_payload_1 = io_pop_s2mPipe_rData_1;
  assign dBus_Bridge_bus_sync_fire_1 = (dBus_Bridge_bus_sync_valid_1 && dBus_Bridge_bus_sync_ready_1);
  assign dBus_Bridge_withWriteBuffer_syncLogic_syncCtx_ready_1 = dBus_Bridge_bus_sync_fire_1;
  assign dBus_Bridge_bus_sync_ready_1 = system_cores_1_logic_cpu_dBus_sync_ready;
  assign system_cores_1_logic_cpu_dBus_rsp_payload_error = (dBus_Bridge_bus_rsp_payload_fragment_opcode_1 == 1'b1);
  assign dBus_Bridge_bus_rsp_ready_1 = 1'b1;
  assign system_cores_1_logic_cpu_dBus_inv_payload_fragment_address = (dBus_Bridge_bus_inv_payload_address_1 + _zz_dBus_inv_payload_fragment_address_2);
  assign system_cores_1_logic_cpu_dBus_inv_payload_last = 1'b1;
  assign dBus_Bridge_bus_inv_ready_1 = (system_cores_1_logic_cpu_dBus_inv_payload_last && system_cores_1_logic_cpu_dBus_inv_ready);
  assign when_Stream_l445_1 = (! system_cores_1_logic_cpu_dBus_ack_payload_last);
  always @(*) begin
    dBus_ack_thrown_valid_1 = system_cores_1_logic_cpu_dBus_ack_valid;
    if(when_Stream_l445_1) begin
      dBus_ack_thrown_valid_1 = 1'b0;
    end
  end

  always @(*) begin
    system_cores_1_logic_cpu_dBus_ack_ready = dBus_ack_thrown_ready_1;
    if(when_Stream_l445_1) begin
      system_cores_1_logic_cpu_dBus_ack_ready = 1'b1;
    end
  end

  assign dBus_ack_thrown_payload_last_1 = system_cores_1_logic_cpu_dBus_ack_payload_last;
  assign dBus_ack_thrown_payload_fragment_hit_1 = system_cores_1_logic_cpu_dBus_ack_payload_fragment_hit;
  assign dBus_Bridge_bus_ack_valid_1 = dBus_ack_thrown_valid_1;
  assign dBus_ack_thrown_ready_1 = dBus_Bridge_bus_ack_ready_1;
  assign system_cores_1_debugRiscv_halted = system_cores_1_logic_cpu_debugBus_halted;
  assign system_cores_1_debugRiscv_running = system_cores_1_logic_cpu_debugBus_running;
  assign system_cores_1_debugRiscv_unavailable = system_cores_1_logic_cpu_debugBus_unavailable;
  assign system_cores_1_debugRiscv_exception = system_cores_1_logic_cpu_debugBus_exception;
  assign system_cores_1_debugRiscv_commit = system_cores_1_logic_cpu_debugBus_commit;
  assign system_cores_1_debugRiscv_ebreak = system_cores_1_logic_cpu_debugBus_ebreak;
  assign system_cores_1_debugRiscv_redo = system_cores_1_logic_cpu_debugBus_redo;
  assign system_cores_1_debugRiscv_regSuccess = system_cores_1_logic_cpu_debugBus_regSuccess;
  assign system_cores_1_debugRiscv_haveReset = system_cores_1_logic_cpu_debugBus_haveReset;
  assign system_cores_1_debugRiscv_resume_rsp_valid = system_cores_1_logic_cpu_debugBus_resume_rsp_valid;
  assign system_cores_1_debugRiscv_hartToDm_valid = system_cores_1_logic_cpu_debugBus_hartToDm_valid;
  assign system_cores_1_debugRiscv_hartToDm_payload_address = system_cores_1_logic_cpu_debugBus_hartToDm_payload_address;
  assign system_cores_1_debugRiscv_hartToDm_payload_data = system_cores_1_logic_cpu_debugBus_hartToDm_payload_data;
  assign system_cores_0_iBus_cmd_combStage_valid = system_cores_0_iBus_cmd_valid;
  assign system_cores_0_iBus_cmd_ready = system_cores_0_iBus_cmd_combStage_ready;
  assign system_cores_0_iBus_cmd_combStage_payload_last = system_cores_0_iBus_cmd_payload_last;
  assign system_cores_0_iBus_cmd_combStage_payload_fragment_opcode = system_cores_0_iBus_cmd_payload_fragment_opcode;
  assign system_cores_0_iBus_cmd_combStage_payload_fragment_address = system_cores_0_iBus_cmd_payload_fragment_address;
  assign system_cores_0_iBus_cmd_combStage_payload_fragment_length = system_cores_0_iBus_cmd_payload_fragment_length;
  assign system_cores_0_iBus_cmd_combStage_ready = system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_ready;
  always @(*) begin
    _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready = system_cores_0_iBus_rsp_ready;
    if(when_Stream_l375_4) begin
      _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready = 1'b1;
    end
  end

  assign when_Stream_l375_4 = (! _zz_system_cores_0_iBus_rsp_valid);
  assign _zz_system_cores_0_iBus_rsp_valid = _zz_system_cores_0_iBus_rsp_valid_1;
  assign system_cores_0_iBus_rsp_valid = _zz_system_cores_0_iBus_rsp_valid;
  assign system_cores_0_iBus_rsp_payload_last = _zz_system_cores_0_iBus_rsp_payload_last;
  assign system_cores_0_iBus_rsp_payload_fragment_opcode = _zz_system_cores_0_iBus_rsp_payload_fragment_opcode;
  assign system_cores_0_iBus_rsp_payload_fragment_data = _zz_system_cores_0_iBus_rsp_payload_fragment_data;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_valid = system_cores_0_iBus_cmd_combStage_valid;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready = _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_last = system_cores_0_iBus_cmd_combStage_payload_last;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_opcode = system_cores_0_iBus_cmd_combStage_payload_fragment_opcode;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_address = system_cores_0_iBus_cmd_combStage_payload_fragment_address;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_length = system_cores_0_iBus_cmd_combStage_payload_fragment_length;
  assign system_cores_1_iBus_cmd_combStage_valid = system_cores_1_iBus_cmd_valid;
  assign system_cores_1_iBus_cmd_ready = system_cores_1_iBus_cmd_combStage_ready;
  assign system_cores_1_iBus_cmd_combStage_payload_last = system_cores_1_iBus_cmd_payload_last;
  assign system_cores_1_iBus_cmd_combStage_payload_fragment_opcode = system_cores_1_iBus_cmd_payload_fragment_opcode;
  assign system_cores_1_iBus_cmd_combStage_payload_fragment_address = system_cores_1_iBus_cmd_payload_fragment_address;
  assign system_cores_1_iBus_cmd_combStage_payload_fragment_length = system_cores_1_iBus_cmd_payload_fragment_length;
  assign system_cores_1_iBus_cmd_combStage_ready = system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready;
  always @(*) begin
    _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready = system_cores_1_iBus_rsp_ready;
    if(when_Stream_l375_5) begin
      _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready = 1'b1;
    end
  end

  assign when_Stream_l375_5 = (! _zz_system_cores_1_iBus_rsp_valid);
  assign _zz_system_cores_1_iBus_rsp_valid = _zz_system_cores_1_iBus_rsp_valid_1;
  assign system_cores_1_iBus_rsp_valid = _zz_system_cores_1_iBus_rsp_valid;
  assign system_cores_1_iBus_rsp_payload_last = _zz_system_cores_1_iBus_rsp_payload_last;
  assign system_cores_1_iBus_rsp_payload_fragment_opcode = _zz_system_cores_1_iBus_rsp_payload_fragment_opcode;
  assign system_cores_1_iBus_rsp_payload_fragment_data = _zz_system_cores_1_iBus_rsp_payload_fragment_data;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid = system_cores_1_iBus_cmd_combStage_valid;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready = _zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last = system_cores_1_iBus_cmd_combStage_payload_last;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode = system_cores_1_iBus_cmd_combStage_payload_fragment_opcode;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address = system_cores_1_iBus_cmd_combStage_payload_fragment_address;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length = system_cores_1_iBus_cmd_combStage_payload_fragment_length;
  always @(*) begin
    dBus_Bridge_bus_cmd_ready = dBus_Bridge_bus_cmd_m2sPipe_ready;
    if(when_Stream_l375_6) begin
      dBus_Bridge_bus_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l375_6 = (! dBus_Bridge_bus_cmd_m2sPipe_valid);
  assign dBus_Bridge_bus_cmd_m2sPipe_valid = dBus_Bridge_bus_cmd_rValid;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_last = dBus_Bridge_bus_cmd_rData_last;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_opcode = dBus_Bridge_bus_cmd_rData_fragment_opcode;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_exclusive = dBus_Bridge_bus_cmd_rData_fragment_exclusive;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_address = dBus_Bridge_bus_cmd_rData_fragment_address;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_length = dBus_Bridge_bus_cmd_rData_fragment_length;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_data = dBus_Bridge_bus_cmd_rData_fragment_data;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_mask = dBus_Bridge_bus_cmd_rData_fragment_mask;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_context = dBus_Bridge_bus_cmd_rData_fragment_context;
  assign dBus_Bridge_bus_cmd_m2sPipe_ready = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_ready;
  assign dBus_Bridge_bus_rsp_valid = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_valid;
  assign dBus_Bridge_bus_rsp_payload_last = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_last;
  assign dBus_Bridge_bus_rsp_payload_fragment_opcode = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_opcode;
  assign dBus_Bridge_bus_rsp_payload_fragment_exclusive = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_exclusive;
  assign dBus_Bridge_bus_rsp_payload_fragment_data = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_data;
  assign dBus_Bridge_bus_rsp_payload_fragment_context = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_context;
  always @(*) begin
    _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready = dBus_Bridge_bus_inv_ready;
    if(when_Stream_l375_7) begin
      _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready = 1'b1;
    end
  end

  assign when_Stream_l375_7 = (! _zz_dBus_Bridge_bus_inv_valid);
  assign _zz_dBus_Bridge_bus_inv_valid = _zz_dBus_Bridge_bus_inv_valid_1;
  assign dBus_Bridge_bus_inv_valid = _zz_dBus_Bridge_bus_inv_valid;
  assign dBus_Bridge_bus_inv_payload_all = _zz_dBus_Bridge_bus_inv_payload_all;
  assign dBus_Bridge_bus_inv_payload_address = _zz_dBus_Bridge_bus_inv_payload_address;
  assign dBus_Bridge_bus_inv_payload_length = _zz_dBus_Bridge_bus_inv_payload_length;
  always @(*) begin
    dBus_Bridge_bus_ack_ready = dBus_Bridge_bus_ack_m2sPipe_ready;
    if(when_Stream_l375_8) begin
      dBus_Bridge_bus_ack_ready = 1'b1;
    end
  end

  assign when_Stream_l375_8 = (! dBus_Bridge_bus_ack_m2sPipe_valid);
  assign dBus_Bridge_bus_ack_m2sPipe_valid = dBus_Bridge_bus_ack_rValid;
  assign dBus_Bridge_bus_ack_m2sPipe_ready = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_ack_ready;
  always @(*) begin
    _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready = dBus_Bridge_bus_sync_ready;
    if(when_Stream_l375_9) begin
      _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready = 1'b1;
    end
  end

  assign when_Stream_l375_9 = (! _zz_dBus_Bridge_bus_sync_valid);
  assign _zz_dBus_Bridge_bus_sync_valid = _zz_dBus_Bridge_bus_sync_valid_1;
  assign dBus_Bridge_bus_sync_valid = _zz_dBus_Bridge_bus_sync_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_valid = dBus_Bridge_bus_cmd_m2sPipe_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready = dBus_Bridge_bus_rsp_ready;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_last = dBus_Bridge_bus_cmd_m2sPipe_payload_last;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_opcode = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_opcode;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_address = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_address;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_length = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_length;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_data = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_data;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_mask = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_mask;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_context = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_payload_fragment_exclusive = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready = _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_ack_valid = dBus_Bridge_bus_ack_m2sPipe_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready = _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready;
  always @(*) begin
    dBus_Bridge_bus_cmd_ready_1 = dBus_Bridge_bus_cmd_m2sPipe_ready_1;
    if(when_Stream_l375_10) begin
      dBus_Bridge_bus_cmd_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_10 = (! dBus_Bridge_bus_cmd_m2sPipe_valid_1);
  assign dBus_Bridge_bus_cmd_m2sPipe_valid_1 = dBus_Bridge_bus_cmd_rValid_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_last_1 = dBus_Bridge_bus_cmd_rData_last_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_opcode_1 = dBus_Bridge_bus_cmd_rData_fragment_opcode_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_exclusive_1 = dBus_Bridge_bus_cmd_rData_fragment_exclusive_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_address_1 = dBus_Bridge_bus_cmd_rData_fragment_address_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_length_1 = dBus_Bridge_bus_cmd_rData_fragment_length_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_data_1 = dBus_Bridge_bus_cmd_rData_fragment_data_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_mask_1 = dBus_Bridge_bus_cmd_rData_fragment_mask_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_context_1 = dBus_Bridge_bus_cmd_rData_fragment_context_1;
  assign dBus_Bridge_bus_cmd_m2sPipe_ready_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready;
  assign dBus_Bridge_bus_rsp_valid_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid;
  assign dBus_Bridge_bus_rsp_payload_last_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last;
  assign dBus_Bridge_bus_rsp_payload_fragment_opcode_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode;
  assign dBus_Bridge_bus_rsp_payload_fragment_exclusive_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_exclusive;
  assign dBus_Bridge_bus_rsp_payload_fragment_data_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data;
  assign dBus_Bridge_bus_rsp_payload_fragment_context_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_context;
  always @(*) begin
    _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready = dBus_Bridge_bus_inv_ready_1;
    if(when_Stream_l375_11) begin
      _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready = 1'b1;
    end
  end

  assign when_Stream_l375_11 = (! _zz_dBus_Bridge_bus_inv_valid_2);
  assign _zz_dBus_Bridge_bus_inv_valid_2 = _zz_dBus_Bridge_bus_inv_valid_3;
  assign dBus_Bridge_bus_inv_valid_1 = _zz_dBus_Bridge_bus_inv_valid_2;
  assign dBus_Bridge_bus_inv_payload_all_1 = _zz_dBus_Bridge_bus_inv_payload_all_1;
  assign dBus_Bridge_bus_inv_payload_address_1 = _zz_dBus_Bridge_bus_inv_payload_address_1;
  assign dBus_Bridge_bus_inv_payload_length_1 = _zz_dBus_Bridge_bus_inv_payload_length_1;
  always @(*) begin
    dBus_Bridge_bus_ack_ready_1 = dBus_Bridge_bus_ack_m2sPipe_ready_1;
    if(when_Stream_l375_12) begin
      dBus_Bridge_bus_ack_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_12 = (! dBus_Bridge_bus_ack_m2sPipe_valid_1);
  assign dBus_Bridge_bus_ack_m2sPipe_valid_1 = dBus_Bridge_bus_ack_rValid_1;
  assign dBus_Bridge_bus_ack_m2sPipe_ready_1 = system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_ack_ready;
  always @(*) begin
    _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready = dBus_Bridge_bus_sync_ready_1;
    if(when_Stream_l375_13) begin
      _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready = 1'b1;
    end
  end

  assign when_Stream_l375_13 = (! _zz_dBus_Bridge_bus_sync_valid_2);
  assign _zz_dBus_Bridge_bus_sync_valid_2 = _zz_dBus_Bridge_bus_sync_valid_3;
  assign dBus_Bridge_bus_sync_valid_1 = _zz_dBus_Bridge_bus_sync_valid_2;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid = dBus_Bridge_bus_cmd_m2sPipe_valid_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready = dBus_Bridge_bus_rsp_ready_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last = dBus_Bridge_bus_cmd_m2sPipe_payload_last_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_opcode_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_address_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_length_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_data = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_data_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_mask = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_mask_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_context = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_context_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_exclusive = dBus_Bridge_bus_cmd_m2sPipe_payload_fragment_exclusive_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready = _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_ack_valid = dBus_Bridge_bus_ack_m2sPipe_valid_1;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready = _zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready;
  assign system_peripheralStopTime = system_coreStopTime_buffercc_io_dataOut;
  always @(*) begin
    system_cores_0_logic_cpu_FpuPlugin_port_commit_ready = FpuPlugin_port_commit_m2sPipe_ready;
    if(when_Stream_l375_14) begin
      system_cores_0_logic_cpu_FpuPlugin_port_commit_ready = 1'b1;
    end
  end

  assign when_Stream_l375_14 = (! FpuPlugin_port_commit_m2sPipe_valid);
  assign FpuPlugin_port_commit_m2sPipe_valid = FpuPlugin_port_commit_rValid;
  assign FpuPlugin_port_commit_m2sPipe_payload_opcode = FpuPlugin_port_commit_rData_opcode;
  assign FpuPlugin_port_commit_m2sPipe_payload_rd = FpuPlugin_port_commit_rData_rd;
  assign FpuPlugin_port_commit_m2sPipe_payload_write = FpuPlugin_port_commit_rData_write;
  assign FpuPlugin_port_commit_m2sPipe_payload_value = FpuPlugin_port_commit_rData_value;
  assign FpuPlugin_port_commit_m2sPipe_ready = system_fpu_logic_io_port_0_commit_ready;
  assign io_port_0_rsp_s2mPipe_valid = (system_fpu_logic_io_port_0_rsp_valid || (! io_port_0_rsp_rValidN));
  assign io_port_0_rsp_s2mPipe_payload_value = (io_port_0_rsp_rValidN ? system_fpu_logic_io_port_0_rsp_payload_value : io_port_0_rsp_rData_value);
  assign io_port_0_rsp_s2mPipe_payload_NV = (io_port_0_rsp_rValidN ? system_fpu_logic_io_port_0_rsp_payload_NV : io_port_0_rsp_rData_NV);
  assign io_port_0_rsp_s2mPipe_payload_NX = (io_port_0_rsp_rValidN ? system_fpu_logic_io_port_0_rsp_payload_NX : io_port_0_rsp_rData_NX);
  assign io_port_0_rsp_s2mPipe_ready = system_cores_0_logic_cpu_FpuPlugin_port_rsp_ready;
  always @(*) begin
    system_cores_1_logic_cpu_FpuPlugin_port_commit_ready = FpuPlugin_port_commit_m2sPipe_ready_1;
    if(when_Stream_l375_15) begin
      system_cores_1_logic_cpu_FpuPlugin_port_commit_ready = 1'b1;
    end
  end

  assign when_Stream_l375_15 = (! FpuPlugin_port_commit_m2sPipe_valid_1);
  assign FpuPlugin_port_commit_m2sPipe_valid_1 = FpuPlugin_port_commit_rValid_1;
  assign FpuPlugin_port_commit_m2sPipe_payload_opcode_1 = FpuPlugin_port_commit_rData_opcode_1;
  assign FpuPlugin_port_commit_m2sPipe_payload_rd_1 = FpuPlugin_port_commit_rData_rd_1;
  assign FpuPlugin_port_commit_m2sPipe_payload_write_1 = FpuPlugin_port_commit_rData_write_1;
  assign FpuPlugin_port_commit_m2sPipe_payload_value_1 = FpuPlugin_port_commit_rData_value_1;
  assign FpuPlugin_port_commit_m2sPipe_ready_1 = system_fpu_logic_io_port_1_commit_ready;
  assign io_port_1_rsp_s2mPipe_valid = (system_fpu_logic_io_port_1_rsp_valid || (! io_port_1_rsp_rValidN));
  assign io_port_1_rsp_s2mPipe_payload_value = (io_port_1_rsp_rValidN ? system_fpu_logic_io_port_1_rsp_payload_value : io_port_1_rsp_rData_value);
  assign io_port_1_rsp_s2mPipe_payload_NV = (io_port_1_rsp_rValidN ? system_fpu_logic_io_port_1_rsp_payload_NV : io_port_1_rsp_rData_NV);
  assign io_port_1_rsp_s2mPipe_payload_NX = (io_port_1_rsp_rValidN ? system_fpu_logic_io_port_1_rsp_payload_NX : io_port_1_rsp_rData_NX);
  assign io_port_1_rsp_s2mPipe_ready = system_cores_1_logic_cpu_FpuPlugin_port_rsp_ready;
  assign cpu0_customInstruction_cmd_valid = system_cores_0_logic_cpu_CfuPlugin_bus_cmd_valid;
  assign cpu0_customInstruction_function_id = system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_function_id;
  assign cpu0_customInstruction_inputs_0 = system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_0;
  assign cpu0_customInstruction_inputs_1 = system_cores_0_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_1;
  assign cpu0_customInstruction_rsp_ready = system_cores_0_logic_cpu_CfuPlugin_bus_rsp_ready;
  assign cpu1_customInstruction_cmd_valid = system_cores_1_logic_cpu_CfuPlugin_bus_cmd_valid;
  assign cpu1_customInstruction_function_id = system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_function_id;
  assign cpu1_customInstruction_inputs_0 = system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_0;
  assign cpu1_customInstruction_inputs_1 = system_cores_1_logic_cpu_CfuPlugin_bus_cmd_payload_inputs_1;
  assign cpu1_customInstruction_rsp_ready = system_cores_1_logic_cpu_CfuPlugin_bus_rsp_ready;
  assign system_riscvJtag_debug_systemReset = system_riscvJtag_debug_logic_dm_io_ndmreset;
  assign system_cores_0_debugRiscv_ackReset = system_riscvJtag_debug_logic_dm_io_harts_0_ackReset;
  assign system_cores_0_debugRiscv_resume_cmd_valid = system_riscvJtag_debug_logic_dm_io_harts_0_resume_cmd_valid;
  assign system_cores_0_debugRiscv_haltReq = system_riscvJtag_debug_logic_dm_io_harts_0_haltReq;
  assign system_cores_0_debugRiscv_dmToHart_valid = io_harts_0_dmToHart_regNext_valid;
  assign system_cores_0_debugRiscv_dmToHart_payload_op = io_harts_0_dmToHart_regNext_payload_op;
  assign system_cores_0_debugRiscv_dmToHart_payload_address = io_harts_0_dmToHart_regNext_payload_address;
  assign system_cores_0_debugRiscv_dmToHart_payload_data = io_harts_0_dmToHart_regNext_payload_data;
  assign system_cores_0_debugRiscv_dmToHart_payload_size = io_harts_0_dmToHart_regNext_payload_size;
  assign system_cores_1_debugRiscv_ackReset = system_riscvJtag_debug_logic_dm_io_harts_1_ackReset;
  assign system_cores_1_debugRiscv_resume_cmd_valid = system_riscvJtag_debug_logic_dm_io_harts_1_resume_cmd_valid;
  assign system_cores_1_debugRiscv_haltReq = system_riscvJtag_debug_logic_dm_io_harts_1_haltReq;
  assign system_cores_1_debugRiscv_dmToHart_valid = io_harts_1_dmToHart_regNext_valid;
  assign system_cores_1_debugRiscv_dmToHart_payload_op = io_harts_1_dmToHart_regNext_payload_op;
  assign system_cores_1_debugRiscv_dmToHart_payload_address = io_harts_1_dmToHart_regNext_payload_address;
  assign system_cores_1_debugRiscv_dmToHart_payload_data = io_harts_1_dmToHart_regNext_payload_data;
  assign system_cores_1_debugRiscv_dmToHart_payload_size = io_harts_1_dmToHart_regNext_payload_size;
  assign system_riscvJtag_debug_systemReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_fabric_iBus_bmb_cmd_valid = system_fabric_iBus_bmb_arbiter_io_output_cmd_valid;
  assign system_fabric_iBus_bmb_rsp_ready = system_fabric_iBus_bmb_arbiter_io_output_rsp_ready;
  assign system_fabric_iBus_bmb_cmd_payload_last = system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_last;
  assign system_fabric_iBus_bmb_cmd_payload_fragment_source = system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_source;
  assign system_fabric_iBus_bmb_cmd_payload_fragment_opcode = system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_opcode;
  assign system_fabric_iBus_bmb_cmd_payload_fragment_address = system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_address;
  assign system_fabric_iBus_bmb_cmd_payload_fragment_length = system_fabric_iBus_bmb_arbiter_io_output_cmd_payload_fragment_length;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready = system_fabric_iBus_bmb_arbiter_io_inputs_0_cmd_ready;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid = system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_valid;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last = system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_last;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode = system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data = system_fabric_iBus_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_ready = system_fabric_iBus_bmb_arbiter_io_inputs_1_cmd_ready;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_valid = system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_valid;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_last = system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_last;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_opcode = system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode;
  assign system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_data = system_fabric_iBus_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data;
  assign system_fabric_invalidationMonitor_logic_input_cmd_ready = system_fabric_invalidationMonitor_logic_monitor_io_input_cmd_ready;
  assign system_fabric_invalidationMonitor_logic_input_rsp_valid = system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_valid;
  assign system_fabric_invalidationMonitor_logic_input_rsp_payload_last = system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_last;
  assign system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_source = system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_source;
  assign system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_opcode = system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_opcode;
  assign system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_data = system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_data;
  assign system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_context = system_fabric_invalidationMonitor_logic_monitor_io_input_rsp_payload_fragment_context;
  assign system_fabric_invalidationMonitor_logic_input_inv_valid = system_fabric_invalidationMonitor_logic_monitor_io_input_inv_valid;
  assign system_fabric_invalidationMonitor_logic_input_ack_ready = system_fabric_invalidationMonitor_logic_monitor_io_input_ack_ready;
  assign system_fabric_invalidationMonitor_logic_input_inv_payload_source = system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_source;
  assign system_fabric_invalidationMonitor_logic_input_inv_payload_address = system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_address;
  assign system_fabric_invalidationMonitor_logic_input_inv_payload_length = system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_length;
  assign system_fabric_invalidationMonitor_logic_input_inv_payload_all = system_fabric_invalidationMonitor_logic_monitor_io_input_inv_payload_all;
  assign system_fabric_invalidationMonitor_logic_input_sync_valid = system_fabric_invalidationMonitor_logic_monitor_io_input_sync_valid;
  assign system_fabric_invalidationMonitor_logic_input_sync_payload_source = system_fabric_invalidationMonitor_logic_monitor_io_input_sync_payload_source;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_valid = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_ready;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_last = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_source = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_opcode = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_address = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_length = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_data = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_mask = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_context = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_ready = system_fabric_invalidationMonitor_logic_input_cmd_ready;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_fabric_invalidationMonitor_logic_input_rsp_valid;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_fabric_invalidationMonitor_logic_input_rsp_payload_last;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_source;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_opcode;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_data;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_fabric_invalidationMonitor_logic_input_rsp_payload_fragment_context;
  assign _zz_system_fabric_invalidationMonitor_logic_input_inv_ready = _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid = (_zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid || (! _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1));
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all = (_zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1 ? _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all : _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all_1);
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address = (_zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1 ? _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address : _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address_1);
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length = (_zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1 ? _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length : _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length_1);
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source = (_zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1 ? _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source : _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source_1);
  always @(*) begin
    system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_m2sPipe_ready;
    if(when_Stream_l375_16) begin
      system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready = 1'b1;
    end
  end

  assign when_Stream_l375_16 = (! system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_m2sPipe_valid);
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_m2sPipe_valid = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_rValid;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_m2sPipe_ready = system_fabric_invalidationMonitor_logic_input_ack_ready;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_valid = system_fabric_invalidationMonitor_logic_input_sync_valid;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_payload_source = system_fabric_invalidationMonitor_logic_input_sync_payload_source;
  assign system_fabric_invalidationMonitor_logic_input_cmd_valid = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_valid;
  assign system_fabric_invalidationMonitor_logic_input_rsp_ready = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_last = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_last;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_source = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_source;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_opcode = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_opcode;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_address = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_address;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_length = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_length;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_data = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_data;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_mask = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_mask;
  assign system_fabric_invalidationMonitor_logic_input_cmd_payload_fragment_context = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_context;
  assign _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid = system_fabric_invalidationMonitor_logic_input_inv_valid;
  assign system_fabric_invalidationMonitor_logic_input_inv_ready = _zz_system_fabric_invalidationMonitor_logic_input_inv_ready;
  assign system_fabric_invalidationMonitor_logic_input_ack_valid = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_m2sPipe_valid;
  assign _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source = system_fabric_invalidationMonitor_logic_input_inv_payload_source;
  assign _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address = system_fabric_invalidationMonitor_logic_input_inv_payload_address;
  assign _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length = system_fabric_invalidationMonitor_logic_input_inv_payload_length;
  assign _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all = system_fabric_invalidationMonitor_logic_input_inv_payload_all;
  assign system_fabric_invalidationMonitor_logic_input_sync_ready = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_ready;
  assign io_output_cmd_s2mPipe_valid = (system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_valid || (! io_output_cmd_rValidN));
  assign io_output_cmd_s2mPipe_payload_last = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_last : io_output_cmd_rData_last);
  assign io_output_cmd_s2mPipe_payload_fragment_source = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_source : io_output_cmd_rData_fragment_source);
  assign io_output_cmd_s2mPipe_payload_fragment_opcode = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_opcode : io_output_cmd_rData_fragment_opcode);
  assign io_output_cmd_s2mPipe_payload_fragment_address = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_address : io_output_cmd_rData_fragment_address);
  assign io_output_cmd_s2mPipe_payload_fragment_length = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_length : io_output_cmd_rData_fragment_length);
  assign io_output_cmd_s2mPipe_payload_fragment_data = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_data : io_output_cmd_rData_fragment_data);
  assign io_output_cmd_s2mPipe_payload_fragment_mask = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_mask : io_output_cmd_rData_fragment_mask);
  assign io_output_cmd_s2mPipe_payload_fragment_context = (io_output_cmd_rValidN ? system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_context : io_output_cmd_rData_fragment_context);
  always @(*) begin
    io_output_cmd_s2mPipe_ready = io_output_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_17) begin
      io_output_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_17 = (! io_output_cmd_s2mPipe_m2sPipe_valid);
  assign io_output_cmd_s2mPipe_m2sPipe_valid = io_output_cmd_s2mPipe_rValid;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_last = io_output_cmd_s2mPipe_rData_last;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_fragment_source = io_output_cmd_s2mPipe_rData_fragment_source;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_fragment_opcode = io_output_cmd_s2mPipe_rData_fragment_opcode;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_fragment_address = io_output_cmd_s2mPipe_rData_fragment_address;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_fragment_length = io_output_cmd_s2mPipe_rData_fragment_length;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_fragment_data = io_output_cmd_s2mPipe_rData_fragment_data;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_fragment_mask = io_output_cmd_s2mPipe_rData_fragment_mask;
  assign io_output_cmd_s2mPipe_m2sPipe_payload_fragment_context = io_output_cmd_s2mPipe_rData_fragment_context;
  assign io_output_cmd_s2mPipe_m2sPipe_ready = system_fabric_invalidationMonitor_output_connector_decoder_cmd_ready;
  always @(*) begin
    _zz_system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready = system_fabric_invalidationMonitor_logic_monitor_io_output_rsp_ready;
    if(when_Stream_l375_18) begin
      _zz_system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready = 1'b1;
    end
  end

  assign when_Stream_l375_18 = (! _zz_when_Stream_l375);
  assign _zz_when_Stream_l375 = _zz_when_Stream_l375_1;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_valid = io_output_cmd_s2mPipe_m2sPipe_valid;
  assign system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready = _zz_system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_last = io_output_cmd_s2mPipe_m2sPipe_payload_last;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_source = io_output_cmd_s2mPipe_m2sPipe_payload_fragment_source;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_opcode = io_output_cmd_s2mPipe_m2sPipe_payload_fragment_opcode;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_address = io_output_cmd_s2mPipe_m2sPipe_payload_fragment_address;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_length = io_output_cmd_s2mPipe_m2sPipe_payload_fragment_length;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_data = io_output_cmd_s2mPipe_m2sPipe_payload_fragment_data;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_mask = io_output_cmd_s2mPipe_m2sPipe_payload_fragment_mask;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_context = io_output_cmd_s2mPipe_m2sPipe_payload_fragment_context;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid || (! system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN));
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_exclusive = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_exclusive : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_exclusive);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context = (system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context : system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context);
  always @(*) begin
    system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_19) begin
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_19 = (! system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid);
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_exclusive = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_exclusive;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready = system_fabric_exclusiveMonitor_logic_io_input_cmd_ready;
  always @(*) begin
    _zz_io_input_rsp_ready = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
    if(when_Stream_l375_20) begin
      _zz_io_input_rsp_ready = 1'b1;
    end
  end

  assign when_Stream_l375_20 = (! _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid);
  assign _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_exclusive = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_exclusive;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid = system_fabric_exclusiveMonitor_logic_io_input_inv_valid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all = system_fabric_exclusiveMonitor_logic_io_input_inv_payload_all;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address = system_fabric_exclusiveMonitor_logic_io_input_inv_payload_address;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length = system_fabric_exclusiveMonitor_logic_io_input_inv_payload_length;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source = system_fabric_exclusiveMonitor_logic_io_input_inv_payload_source;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_combStage_valid = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_valid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_combStage_ready;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_combStage_ready = system_fabric_exclusiveMonitor_logic_io_input_ack_ready;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_valid = system_fabric_exclusiveMonitor_logic_io_input_sync_valid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_payload_source = system_fabric_exclusiveMonitor_logic_io_input_sync_payload_source;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_valid = system_fabric_exclusiveMonitor_logic_io_output_cmd_valid;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_rsp_ready = system_fabric_exclusiveMonitor_logic_io_output_rsp_ready;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_last = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_last;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_source = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_source;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_opcode = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_opcode;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_address = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_address;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_length = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_length;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_data = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_data;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_mask = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_mask;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_context = system_fabric_exclusiveMonitor_logic_io_output_cmd_payload_fragment_context;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_inv_ready = system_fabric_exclusiveMonitor_logic_io_output_inv_ready;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_ack_valid = system_fabric_exclusiveMonitor_logic_io_output_ack_valid;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_sync_ready = system_fabric_exclusiveMonitor_logic_io_output_sync_ready;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_valid;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_cmd_ready = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_rsp_valid = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_fabric_exclusiveMonitor_output_connector_decoder_rsp_ready;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_last;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_last = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_source;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_opcode;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_address;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_length;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_data;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_mask;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_fabric_exclusiveMonitor_output_connector_decoder_cmd_payload_fragment_context;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_source = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_opcode = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_data = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_rsp_payload_fragment_context = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_inv_valid = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_ready = system_fabric_exclusiveMonitor_output_connector_decoder_inv_ready;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_valid = system_fabric_exclusiveMonitor_output_connector_decoder_ack_valid;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_ack_ready = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_source = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_address = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_length = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_inv_payload_all = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_sync_valid = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_valid;
  assign system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_ready = system_fabric_exclusiveMonitor_output_connector_decoder_sync_ready;
  assign system_fabric_exclusiveMonitor_output_connector_decoder_sync_payload_source = system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_payload_source;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_valid = system_fabric_dBusCoherent_bmb_cmd_valid;
  assign system_fabric_dBusCoherent_bmb_cmd_ready = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_ready;
  assign system_fabric_dBusCoherent_bmb_rsp_valid = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_valid;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_ready = system_fabric_dBusCoherent_bmb_rsp_ready;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_last = system_fabric_dBusCoherent_bmb_cmd_payload_last;
  assign system_fabric_dBusCoherent_bmb_rsp_payload_last = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_last;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_source = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_source;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_opcode = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_opcode;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_address = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_address;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_length = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_length;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_data = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_data;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_mask = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_mask;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_context = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_exclusive = system_fabric_dBusCoherent_bmb_cmd_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_rsp_payload_fragment_source = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_source;
  assign system_fabric_dBusCoherent_bmb_rsp_payload_fragment_opcode = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_opcode;
  assign system_fabric_dBusCoherent_bmb_rsp_payload_fragment_data = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_data;
  assign system_fabric_dBusCoherent_bmb_rsp_payload_fragment_context = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_rsp_payload_fragment_exclusive = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_inv_valid = system_fabric_dBusCoherent_bmb_connector_decoder_inv_valid;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_inv_ready = system_fabric_dBusCoherent_bmb_inv_ready;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_ack_valid = system_fabric_dBusCoherent_bmb_ack_valid;
  assign system_fabric_dBusCoherent_bmb_ack_ready = system_fabric_dBusCoherent_bmb_connector_decoder_ack_ready;
  assign system_fabric_dBusCoherent_bmb_inv_payload_source = system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_source;
  assign system_fabric_dBusCoherent_bmb_inv_payload_address = system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_address;
  assign system_fabric_dBusCoherent_bmb_inv_payload_length = system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_length;
  assign system_fabric_dBusCoherent_bmb_inv_payload_all = system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_all;
  assign system_fabric_dBusCoherent_bmb_sync_valid = system_fabric_dBusCoherent_bmb_connector_decoder_sync_valid;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_sync_ready = system_fabric_dBusCoherent_bmb_sync_ready;
  assign system_fabric_dBusCoherent_bmb_sync_payload_source = system_fabric_dBusCoherent_bmb_connector_decoder_sync_payload_source;
  assign system_fabric_dBus_bmb_cmd_valid = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_fabric_dBus_bmb_cmd_ready;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_fabric_dBus_bmb_rsp_valid;
  assign system_fabric_dBus_bmb_rsp_ready = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  assign system_fabric_dBus_bmb_cmd_payload_last = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_fabric_dBus_bmb_rsp_payload_last;
  assign system_fabric_dBus_bmb_cmd_payload_fragment_source = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
  assign system_fabric_dBus_bmb_cmd_payload_fragment_opcode = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  assign system_fabric_dBus_bmb_cmd_payload_fragment_address = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  assign system_fabric_dBus_bmb_cmd_payload_fragment_length = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  assign system_fabric_dBus_bmb_cmd_payload_fragment_data = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  assign system_fabric_dBus_bmb_cmd_payload_fragment_mask = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  assign system_fabric_dBus_bmb_cmd_payload_fragment_context = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = system_fabric_dBus_bmb_rsp_payload_fragment_source;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_fabric_dBus_bmb_rsp_payload_fragment_opcode;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_fabric_dBus_bmb_rsp_payload_fragment_data;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_fabric_dBus_bmb_rsp_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_cmd_valid = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_valid;
  assign system_fabric_dBusCoherent_bmb_rsp_ready = system_fabric_dBusCoherent_bmb_arbiter_io_output_rsp_ready;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_last = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_last;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_source = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_source;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_opcode = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_opcode;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_address = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_address;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_length = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_length;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_data = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_data;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_mask = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_mask;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_context = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_cmd_payload_fragment_exclusive = system_fabric_dBusCoherent_bmb_arbiter_io_output_cmd_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_inv_ready = system_fabric_dBusCoherent_bmb_arbiter_io_output_inv_ready;
  assign system_fabric_dBusCoherent_bmb_ack_valid = system_fabric_dBusCoherent_bmb_arbiter_io_output_ack_valid;
  assign system_fabric_dBusCoherent_bmb_sync_ready = system_fabric_dBusCoherent_bmb_arbiter_io_output_sync_ready;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_valid;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_cmd_ready = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_valid = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_fabric_dBusCoherent_bmb_connector_decoder_rsp_ready;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_last;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_last = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_source;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_opcode;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_address;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_length;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_data;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_mask;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_context;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_exclusive = system_fabric_dBusCoherent_bmb_connector_decoder_cmd_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_source = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_opcode = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_data = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_context = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_rsp_payload_fragment_exclusive = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_inv_valid = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_ready = system_fabric_dBusCoherent_bmb_connector_decoder_inv_ready;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_valid = system_fabric_dBusCoherent_bmb_connector_decoder_ack_valid;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_ack_ready = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_source = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_address = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_length = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_inv_payload_all = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_sync_valid = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_valid;
  assign system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_ready = system_fabric_dBusCoherent_bmb_connector_decoder_sync_ready;
  assign system_fabric_dBusCoherent_bmb_connector_decoder_sync_payload_source = system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_sync_payload_source;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_fabric_invalidationMonitor_output_connector_decoder_cmd_valid;
  assign system_fabric_invalidationMonitor_output_connector_decoder_cmd_ready = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_fabric_invalidationMonitor_output_connector_decoder_rsp_valid = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_last;
  assign system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_last = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_source;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_opcode;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_address;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_length;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_data;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_mask;
  assign system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_fabric_invalidationMonitor_output_connector_decoder_cmd_payload_fragment_context;
  assign system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_source = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  assign system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_opcode = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_data = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_context = system_fabric_dBus_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_cmd_ready;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_last;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_context = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_exclusive = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_rsp_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_valid = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_ack_ready = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_ack_ready;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_address = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_address;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_length = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_length;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_all = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_inv_payload_all;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_valid = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_0_sync_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_cmd_ready = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_cmd_ready;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_valid = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_last = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_last;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_opcode = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_opcode;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_data = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_data;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_context = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_context;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_exclusive = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_rsp_payload_fragment_exclusive;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_valid = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_valid;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_ack_ready = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_ack_ready;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_address = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_address;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_length = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_length;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_all = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_inv_payload_all;
  assign system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_valid = system_fabric_dBusCoherent_bmb_arbiter_io_inputs_1_sync_valid;
  always @(*) begin
    system_fabric_iBus_bmb_cmd_ready = system_fabric_iBus_bmb_cmd_m2sPipe_ready;
    if(when_Stream_l375_21) begin
      system_fabric_iBus_bmb_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l375_21 = (! system_fabric_iBus_bmb_cmd_m2sPipe_valid);
  assign system_fabric_iBus_bmb_cmd_m2sPipe_valid = system_fabric_iBus_bmb_cmd_rValid;
  assign system_fabric_iBus_bmb_cmd_m2sPipe_payload_last = system_fabric_iBus_bmb_cmd_rData_last;
  assign system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_source = system_fabric_iBus_bmb_cmd_rData_fragment_source;
  assign system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_opcode = system_fabric_iBus_bmb_cmd_rData_fragment_opcode;
  assign system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_address = system_fabric_iBus_bmb_cmd_rData_fragment_address;
  assign system_fabric_iBus_bmb_cmd_m2sPipe_payload_fragment_length = system_fabric_iBus_bmb_cmd_rData_fragment_length;
  assign system_fabric_iBus_bmb_cmd_m2sPipe_ready = system_fabric_iBus_bmb_decoder_io_input_cmd_ready;
  assign system_fabric_iBus_bmb_rsp_valid = system_fabric_iBus_bmb_decoder_io_input_rsp_valid;
  assign system_fabric_iBus_bmb_rsp_payload_last = system_fabric_iBus_bmb_decoder_io_input_rsp_payload_last;
  assign system_fabric_iBus_bmb_rsp_payload_fragment_source = system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_source;
  assign system_fabric_iBus_bmb_rsp_payload_fragment_opcode = system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_opcode;
  assign system_fabric_iBus_bmb_rsp_payload_fragment_data = system_fabric_iBus_bmb_decoder_io_input_rsp_payload_fragment_data;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_valid = system_fabric_dBus_bmb_cmd_valid;
  assign system_fabric_dBus_bmb_cmd_ready = system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready;
  assign system_fabric_dBus_bmb_rsp_valid = system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready = system_fabric_dBus_bmb_rsp_ready;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_last = system_fabric_dBus_bmb_cmd_payload_last;
  assign system_fabric_dBus_bmb_rsp_payload_last = system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_source = system_fabric_dBus_bmb_cmd_payload_fragment_source;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_opcode = system_fabric_dBus_bmb_cmd_payload_fragment_opcode;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_address = system_fabric_dBus_bmb_cmd_payload_fragment_address;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_length = system_fabric_dBus_bmb_cmd_payload_fragment_length;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_data = system_fabric_dBus_bmb_cmd_payload_fragment_data;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_mask = system_fabric_dBus_bmb_cmd_payload_fragment_mask;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_payload_fragment_context = system_fabric_dBus_bmb_cmd_payload_fragment_context;
  assign system_fabric_dBus_bmb_rsp_payload_fragment_source = system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_source;
  assign system_fabric_dBus_bmb_rsp_payload_fragment_opcode = system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode;
  assign system_fabric_dBus_bmb_rsp_payload_fragment_data = system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data;
  assign system_fabric_dBus_bmb_rsp_payload_fragment_context = system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_context;
  assign system_bridge_bmb_cmd_valid = system_bridge_bmb_arbiter_io_output_cmd_valid;
  assign system_bridge_bmb_rsp_ready = system_bridge_bmb_arbiter_io_output_rsp_ready;
  assign system_bridge_bmb_cmd_payload_last = system_bridge_bmb_arbiter_io_output_cmd_payload_last;
  assign system_bridge_bmb_cmd_payload_fragment_source = system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_source;
  assign system_bridge_bmb_cmd_payload_fragment_opcode = system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_opcode;
  assign system_bridge_bmb_cmd_payload_fragment_address = system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_address;
  assign system_bridge_bmb_cmd_payload_fragment_length = system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_length;
  assign system_bridge_bmb_cmd_payload_fragment_data = system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_data;
  assign system_bridge_bmb_cmd_payload_fragment_mask = system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_mask;
  assign system_bridge_bmb_cmd_payload_fragment_context = system_bridge_bmb_arbiter_io_output_cmd_payload_fragment_context;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_cmd_ready = system_bridge_bmb_arbiter_io_inputs_0_cmd_ready;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid = system_bridge_bmb_arbiter_io_inputs_0_rsp_valid;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last = system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_last;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_source = system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_source;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode = system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_opcode;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data = system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_data;
  assign system_bridge_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_context = system_bridge_bmb_arbiter_io_inputs_0_rsp_payload_fragment_context;
  always @(*) begin
    system_ddr_ddrLogic_cc_fifo_io_output_cmd_ready = io_output_cmd_m2sPipe_ready;
    if(when_Stream_l375_22) begin
      system_ddr_ddrLogic_cc_fifo_io_output_cmd_ready = 1'b1;
    end
  end

  assign when_Stream_l375_22 = (! io_output_cmd_m2sPipe_valid);
  assign io_output_cmd_m2sPipe_valid = io_output_cmd_rValid;
  assign io_output_cmd_m2sPipe_payload_last = io_output_cmd_rData_last_1;
  assign io_output_cmd_m2sPipe_payload_fragment_source = io_output_cmd_rData_fragment_source_1;
  assign io_output_cmd_m2sPipe_payload_fragment_opcode = io_output_cmd_rData_fragment_opcode_1;
  assign io_output_cmd_m2sPipe_payload_fragment_address = io_output_cmd_rData_fragment_address_1;
  assign io_output_cmd_m2sPipe_payload_fragment_length = io_output_cmd_rData_fragment_length_1;
  assign io_output_cmd_m2sPipe_payload_fragment_data = io_output_cmd_rData_fragment_data_1;
  assign io_output_cmd_m2sPipe_payload_fragment_mask = io_output_cmd_rData_fragment_mask_1;
  assign io_output_cmd_m2sPipe_payload_fragment_context = io_output_cmd_rData_fragment_context_1;
  assign io_output_cmd_m2sPipe_ready = system_ddr_ddrLogic_bmbToAxiBridge_io_input_cmd_ready;
  always @(*) begin
    _zz_io_input_rsp_ready_1 = system_ddr_ddrLogic_cc_fifo_io_output_rsp_ready;
    if(when_Stream_l375_23) begin
      _zz_io_input_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_23 = (! _zz_when_Stream_l375_2);
  assign _zz_when_Stream_l375_2 = _zz_when_Stream_l375_3;
  assign io_output_arw_s2mPipe_valid = (system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_valid || (! io_output_arw_rValidN));
  assign io_output_arw_s2mPipe_payload_addr = (io_output_arw_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_addr : io_output_arw_rData_addr);
  assign io_output_arw_s2mPipe_payload_len = (io_output_arw_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_len : io_output_arw_rData_len);
  assign io_output_arw_s2mPipe_payload_size = (io_output_arw_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_size : io_output_arw_rData_size);
  assign io_output_arw_s2mPipe_payload_cache = (io_output_arw_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_cache : io_output_arw_rData_cache);
  assign io_output_arw_s2mPipe_payload_prot = (io_output_arw_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_prot : io_output_arw_rData_prot);
  assign io_output_arw_s2mPipe_payload_write = (io_output_arw_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_write : io_output_arw_rData_write);
  always @(*) begin
    io_output_arw_s2mPipe_ready = io_output_arw_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_24) begin
      io_output_arw_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_24 = (! io_output_arw_s2mPipe_m2sPipe_valid);
  assign io_output_arw_s2mPipe_m2sPipe_valid = io_output_arw_s2mPipe_rValid;
  assign io_output_arw_s2mPipe_m2sPipe_payload_addr = io_output_arw_s2mPipe_rData_addr;
  assign io_output_arw_s2mPipe_m2sPipe_payload_len = io_output_arw_s2mPipe_rData_len;
  assign io_output_arw_s2mPipe_m2sPipe_payload_size = io_output_arw_s2mPipe_rData_size;
  assign io_output_arw_s2mPipe_m2sPipe_payload_cache = io_output_arw_s2mPipe_rData_cache;
  assign io_output_arw_s2mPipe_m2sPipe_payload_prot = io_output_arw_s2mPipe_rData_prot;
  assign io_output_arw_s2mPipe_m2sPipe_payload_write = io_output_arw_s2mPipe_rData_write;
  always @(*) begin
    io_output_arw_s2mPipe_m2sPipe_ready = io_output_arw_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l375_25) begin
      io_output_arw_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_25 = (! io_output_arw_s2mPipe_m2sPipe_m2sPipe_valid);
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_valid = io_output_arw_s2mPipe_m2sPipe_rValid;
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_addr = io_output_arw_s2mPipe_m2sPipe_rData_addr;
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_len = io_output_arw_s2mPipe_m2sPipe_rData_len;
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_size = io_output_arw_s2mPipe_m2sPipe_rData_size;
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_cache = io_output_arw_s2mPipe_m2sPipe_rData_cache;
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_prot = io_output_arw_s2mPipe_m2sPipe_rData_prot;
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_write = io_output_arw_s2mPipe_m2sPipe_rData_write;
  assign system_ddr_ddrLogic_cpuAccess_arw_valid = io_output_arw_s2mPipe_m2sPipe_m2sPipe_valid;
  assign io_output_arw_s2mPipe_m2sPipe_m2sPipe_ready = system_ddr_ddrLogic_cpuAccess_arw_ready;
  assign system_ddr_ddrLogic_cpuAccess_arw_payload_addr = io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_addr;
  assign system_ddr_ddrLogic_cpuAccess_arw_payload_len = io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_len;
  assign system_ddr_ddrLogic_cpuAccess_arw_payload_size = io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_size;
  assign system_ddr_ddrLogic_cpuAccess_arw_payload_cache = io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_cache;
  assign system_ddr_ddrLogic_cpuAccess_arw_payload_prot = io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_prot;
  assign system_ddr_ddrLogic_cpuAccess_arw_payload_write = io_output_arw_s2mPipe_m2sPipe_m2sPipe_payload_write;
  assign io_output_w_s2mPipe_valid = (system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_valid || (! io_output_w_rValidN));
  assign io_output_w_s2mPipe_payload_data = (io_output_w_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_data : io_output_w_rData_data);
  assign io_output_w_s2mPipe_payload_strb = (io_output_w_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_strb : io_output_w_rData_strb);
  assign io_output_w_s2mPipe_payload_last = (io_output_w_rValidN ? system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_last : io_output_w_rData_last);
  always @(*) begin
    io_output_w_s2mPipe_ready = io_output_w_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_26) begin
      io_output_w_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_26 = (! io_output_w_s2mPipe_m2sPipe_valid);
  assign io_output_w_s2mPipe_m2sPipe_valid = io_output_w_s2mPipe_rValid;
  assign io_output_w_s2mPipe_m2sPipe_payload_data = io_output_w_s2mPipe_rData_data;
  assign io_output_w_s2mPipe_m2sPipe_payload_strb = io_output_w_s2mPipe_rData_strb;
  assign io_output_w_s2mPipe_m2sPipe_payload_last = io_output_w_s2mPipe_rData_last;
  always @(*) begin
    io_output_w_s2mPipe_m2sPipe_ready = io_output_w_s2mPipe_m2sPipe_m2sPipe_ready;
    if(when_Stream_l375_27) begin
      io_output_w_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_27 = (! io_output_w_s2mPipe_m2sPipe_m2sPipe_valid);
  assign io_output_w_s2mPipe_m2sPipe_m2sPipe_valid = io_output_w_s2mPipe_m2sPipe_rValid;
  assign io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_data = io_output_w_s2mPipe_m2sPipe_rData_data;
  assign io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_strb = io_output_w_s2mPipe_m2sPipe_rData_strb;
  assign io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_last = io_output_w_s2mPipe_m2sPipe_rData_last;
  assign system_ddr_ddrLogic_cpuAccess_w_valid = io_output_w_s2mPipe_m2sPipe_m2sPipe_valid;
  assign io_output_w_s2mPipe_m2sPipe_m2sPipe_ready = system_ddr_ddrLogic_cpuAccess_w_ready;
  assign system_ddr_ddrLogic_cpuAccess_w_payload_data = io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_data;
  assign system_ddr_ddrLogic_cpuAccess_w_payload_strb = io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_strb;
  assign system_ddr_ddrLogic_cpuAccess_w_payload_last = io_output_w_s2mPipe_m2sPipe_m2sPipe_payload_last;
  assign system_ddr_ddrLogic_cpuAccess_b_ready = system_ddr_ddrLogic_cpuAccess_b_rValidN;
  assign system_ddr_ddrLogic_cpuAccess_b_s2mPipe_valid = (system_ddr_ddrLogic_cpuAccess_b_valid || (! system_ddr_ddrLogic_cpuAccess_b_rValidN));
  assign system_ddr_ddrLogic_cpuAccess_b_s2mPipe_payload_resp = (system_ddr_ddrLogic_cpuAccess_b_rValidN ? system_ddr_ddrLogic_cpuAccess_b_payload_resp : system_ddr_ddrLogic_cpuAccess_b_rData_resp);
  always @(*) begin
    system_ddr_ddrLogic_cpuAccess_b_s2mPipe_ready = system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_28) begin
      system_ddr_ddrLogic_cpuAccess_b_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_28 = (! system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_cpuAccess_b_s2mPipe_rValid;
  assign system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_payload_resp = system_ddr_ddrLogic_cpuAccess_b_s2mPipe_rData_resp;
  assign system_ddr_ddrLogic_cpuAccess_b_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_bmbToAxiBridge_io_output_b_ready;
  assign system_ddr_ddrLogic_cpuAccess_r_ready = system_ddr_ddrLogic_cpuAccess_r_rValidN;
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_valid = (system_ddr_ddrLogic_cpuAccess_r_valid || (! system_ddr_ddrLogic_cpuAccess_r_rValidN));
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_data = (system_ddr_ddrLogic_cpuAccess_r_rValidN ? system_ddr_ddrLogic_cpuAccess_r_payload_data : system_ddr_ddrLogic_cpuAccess_r_rData_data);
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_resp = (system_ddr_ddrLogic_cpuAccess_r_rValidN ? system_ddr_ddrLogic_cpuAccess_r_payload_resp : system_ddr_ddrLogic_cpuAccess_r_rData_resp);
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_last = (system_ddr_ddrLogic_cpuAccess_r_rValidN ? system_ddr_ddrLogic_cpuAccess_r_payload_last : system_ddr_ddrLogic_cpuAccess_r_rData_last);
  always @(*) begin
    system_ddr_ddrLogic_cpuAccess_r_s2mPipe_ready = system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_29) begin
      system_ddr_ddrLogic_cpuAccess_r_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_29 = (! system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rValid;
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_data = system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_data;
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_resp = system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_resp;
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_payload_last = system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_last;
  assign system_ddr_ddrLogic_cpuAccess_r_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_bmbToAxiBridge_io_output_r_ready;
  assign system_ddr_ddrLogic_cpuAccess_arw_ready = (system_ddr_ddrLogic_cpuAccess_arw_payload_write ? system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_aw_ready : system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_ar_ready);
  assign system_ddr_ddrLogic_cpuAccess_w_ready = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_w_ready;
  assign system_ddr_ddrLogic_cpuAccess_r_valid = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_valid;
  assign system_ddr_ddrLogic_cpuAccess_r_payload_data = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_data;
  assign system_ddr_ddrLogic_cpuAccess_r_payload_resp = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_resp;
  assign system_ddr_ddrLogic_cpuAccess_r_payload_last = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_r_payload_last;
  assign system_ddr_ddrLogic_cpuAccess_b_valid = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_valid;
  assign system_ddr_ddrLogic_cpuAccess_b_payload_resp = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_b_payload_resp;
  assign system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_0_ar_valid = (system_ddr_ddrLogic_cpuAccess_arw_valid && (! system_ddr_ddrLogic_cpuAccess_arw_payload_write));
  assign _zz_io_inputs_0_ar_payload_region[3 : 0] = 4'b0000;
  assign system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_0_aw_valid = (system_ddr_ddrLogic_cpuAccess_arw_valid && system_ddr_ddrLogic_cpuAccess_arw_payload_write);
  assign _zz_io_inputs_0_aw_payload_region[3 : 0] = 4'b0000;
  assign io_ddrMasters_1_reset_read_buffer = ddrCd_logic_outputReset_buffercc_io_dataOut;
  assign io_ddrMasters_1_aw_ready = io_ddrMasters_1_aw_rValidN;
  assign io_ddrMasters_1_aw_s2mPipe_valid = (io_ddrMasters_1_aw_valid || (! io_ddrMasters_1_aw_rValidN));
  assign io_ddrMasters_1_aw_s2mPipe_payload_addr = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_addr : io_ddrMasters_1_aw_rData_addr);
  assign io_ddrMasters_1_aw_s2mPipe_payload_id = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_id : io_ddrMasters_1_aw_rData_id);
  assign io_ddrMasters_1_aw_s2mPipe_payload_region = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_region : io_ddrMasters_1_aw_rData_region);
  assign io_ddrMasters_1_aw_s2mPipe_payload_len = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_len : io_ddrMasters_1_aw_rData_len);
  assign io_ddrMasters_1_aw_s2mPipe_payload_size = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_size : io_ddrMasters_1_aw_rData_size);
  assign io_ddrMasters_1_aw_s2mPipe_payload_burst = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_burst : io_ddrMasters_1_aw_rData_burst);
  assign io_ddrMasters_1_aw_s2mPipe_payload_lock = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_lock : io_ddrMasters_1_aw_rData_lock);
  assign io_ddrMasters_1_aw_s2mPipe_payload_cache = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_cache : io_ddrMasters_1_aw_rData_cache);
  assign io_ddrMasters_1_aw_s2mPipe_payload_qos = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_qos : io_ddrMasters_1_aw_rData_qos);
  assign io_ddrMasters_1_aw_s2mPipe_payload_prot = (io_ddrMasters_1_aw_rValidN ? io_ddrMasters_1_aw_payload_prot : io_ddrMasters_1_aw_rData_prot);
  always @(*) begin
    io_ddrMasters_1_aw_s2mPipe_ready = io_ddrMasters_1_aw_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_30) begin
      io_ddrMasters_1_aw_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_30 = (! io_ddrMasters_1_aw_s2mPipe_m2sPipe_valid);
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_valid = io_ddrMasters_1_aw_s2mPipe_rValid;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_addr = io_ddrMasters_1_aw_s2mPipe_rData_addr;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_id = io_ddrMasters_1_aw_s2mPipe_rData_id;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_region = io_ddrMasters_1_aw_s2mPipe_rData_region;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_len = io_ddrMasters_1_aw_s2mPipe_rData_len;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_size = io_ddrMasters_1_aw_s2mPipe_rData_size;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_burst = io_ddrMasters_1_aw_s2mPipe_rData_burst;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_lock = io_ddrMasters_1_aw_s2mPipe_rData_lock;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_cache = io_ddrMasters_1_aw_s2mPipe_rData_cache;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_qos = io_ddrMasters_1_aw_s2mPipe_rData_qos;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_payload_prot = io_ddrMasters_1_aw_s2mPipe_rData_prot;
  assign io_ddrMasters_1_aw_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_0_bridge_io_input_aw_ready;
  assign io_ddrMasters_1_ar_halfPipe_fire = (io_ddrMasters_1_ar_halfPipe_valid && io_ddrMasters_1_ar_halfPipe_ready);
  assign io_ddrMasters_1_ar_ready = (! io_ddrMasters_1_ar_rValid);
  assign io_ddrMasters_1_ar_halfPipe_valid = io_ddrMasters_1_ar_rValid;
  assign io_ddrMasters_1_ar_halfPipe_payload_addr = io_ddrMasters_1_ar_rData_addr;
  assign io_ddrMasters_1_ar_halfPipe_payload_id = io_ddrMasters_1_ar_rData_id;
  assign io_ddrMasters_1_ar_halfPipe_payload_region = io_ddrMasters_1_ar_rData_region;
  assign io_ddrMasters_1_ar_halfPipe_payload_len = io_ddrMasters_1_ar_rData_len;
  assign io_ddrMasters_1_ar_halfPipe_payload_size = io_ddrMasters_1_ar_rData_size;
  assign io_ddrMasters_1_ar_halfPipe_payload_burst = io_ddrMasters_1_ar_rData_burst;
  assign io_ddrMasters_1_ar_halfPipe_payload_lock = io_ddrMasters_1_ar_rData_lock;
  assign io_ddrMasters_1_ar_halfPipe_payload_cache = io_ddrMasters_1_ar_rData_cache;
  assign io_ddrMasters_1_ar_halfPipe_payload_qos = io_ddrMasters_1_ar_rData_qos;
  assign io_ddrMasters_1_ar_halfPipe_payload_prot = io_ddrMasters_1_ar_rData_prot;
  assign io_ddrMasters_1_ar_halfPipe_ready = system_ddr_ddrLogic_userAdapters_0_bridge_io_input_ar_ready;
  assign io_ddrMasters_1_w_ready = io_ddrMasters_1_w_rValidN;
  assign io_ddrMasters_1_w_s2mPipe_valid = (io_ddrMasters_1_w_valid || (! io_ddrMasters_1_w_rValidN));
  assign io_ddrMasters_1_w_s2mPipe_payload_data = (io_ddrMasters_1_w_rValidN ? io_ddrMasters_1_w_payload_data : io_ddrMasters_1_w_rData_data);
  assign io_ddrMasters_1_w_s2mPipe_payload_strb = (io_ddrMasters_1_w_rValidN ? io_ddrMasters_1_w_payload_strb : io_ddrMasters_1_w_rData_strb);
  assign io_ddrMasters_1_w_s2mPipe_payload_last = (io_ddrMasters_1_w_rValidN ? io_ddrMasters_1_w_payload_last : io_ddrMasters_1_w_rData_last);
  always @(*) begin
    io_ddrMasters_1_w_s2mPipe_ready = io_ddrMasters_1_w_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_31) begin
      io_ddrMasters_1_w_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_31 = (! io_ddrMasters_1_w_s2mPipe_m2sPipe_valid);
  assign io_ddrMasters_1_w_s2mPipe_m2sPipe_valid = io_ddrMasters_1_w_s2mPipe_rValid;
  assign io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_data = io_ddrMasters_1_w_s2mPipe_rData_data;
  assign io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_strb = io_ddrMasters_1_w_s2mPipe_rData_strb;
  assign io_ddrMasters_1_w_s2mPipe_m2sPipe_payload_last = io_ddrMasters_1_w_s2mPipe_rData_last;
  assign io_ddrMasters_1_w_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_0_bridge_io_input_w_ready;
  always @(*) begin
    system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_ready = io_input_r_m2sPipe_ready;
    if(when_Stream_l375_32) begin
      system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_ready = 1'b1;
    end
  end

  assign when_Stream_l375_32 = (! io_input_r_m2sPipe_valid);
  assign io_input_r_m2sPipe_valid = io_input_r_rValid;
  assign io_input_r_m2sPipe_payload_data = io_input_r_rData_data;
  assign io_input_r_m2sPipe_payload_id = io_input_r_rData_id;
  assign io_input_r_m2sPipe_payload_resp = io_input_r_rData_resp;
  assign io_input_r_m2sPipe_payload_last = io_input_r_rData_last;
  assign io_ddrMasters_1_r_valid = io_input_r_m2sPipe_valid;
  assign io_input_r_m2sPipe_ready = io_ddrMasters_1_r_ready;
  assign io_ddrMasters_1_r_payload_data = io_input_r_m2sPipe_payload_data;
  assign io_ddrMasters_1_r_payload_id = io_input_r_m2sPipe_payload_id;
  assign io_ddrMasters_1_r_payload_resp = io_input_r_m2sPipe_payload_resp;
  assign io_ddrMasters_1_r_payload_last = io_input_r_m2sPipe_payload_last;
  assign io_input_b_s2mPipe_valid = (system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_valid || (! io_input_b_rValidN));
  assign io_input_b_s2mPipe_payload_id = (io_input_b_rValidN ? system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_id : io_input_b_rData_id);
  assign io_input_b_s2mPipe_payload_resp = (io_input_b_rValidN ? system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_resp : io_input_b_rData_resp);
  always @(*) begin
    io_input_b_s2mPipe_ready = io_input_b_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_33) begin
      io_input_b_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_33 = (! io_input_b_s2mPipe_m2sPipe_valid);
  assign io_input_b_s2mPipe_m2sPipe_valid = io_input_b_s2mPipe_rValid;
  assign io_input_b_s2mPipe_m2sPipe_payload_id = io_input_b_s2mPipe_rData_id;
  assign io_input_b_s2mPipe_m2sPipe_payload_resp = io_input_b_s2mPipe_rData_resp;
  assign io_ddrMasters_1_b_valid = io_input_b_s2mPipe_m2sPipe_valid;
  assign io_input_b_s2mPipe_m2sPipe_ready = io_ddrMasters_1_b_ready;
  assign io_ddrMasters_1_b_payload_id = io_input_b_s2mPipe_m2sPipe_payload_id;
  assign io_ddrMasters_1_b_payload_resp = io_input_b_s2mPipe_m2sPipe_payload_resp;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_valid = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_valid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_addr = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_id = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_id;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_region = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_region;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_len = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_len;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_size = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_size;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_burst = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_lock = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_cache = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_qos = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_prot = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_ar_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_valid = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_valid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_addr = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_id = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_id;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_region = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_region;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_len = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_len;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_size = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_size;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_burst = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_lock = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_cache = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_qos = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_prot = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_aw_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_valid = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_valid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_data = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_data;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_strb = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_strb;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_last = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_w_payload_last;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_r_ready = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_r_ready;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_b_ready = system_ddr_ddrLogic_userAdapters_0_upsizer_logic_io_output_b_ready;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_fire = (system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_valid && system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_ready);
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_ready = (! system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rValid);
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_valid = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rValid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_addr = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_addr;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_id = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_id;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_region = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_region;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_len = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_len;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_size = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_size;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_burst = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_burst;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_lock = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_lock;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_cache = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_cache;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_qos = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_qos;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_prot = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_prot;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_valid = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_ready = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_ready;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_addr = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_id = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_region = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_region;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_len = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_len;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_size = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_size;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_burst = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_lock = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_cache = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_qos = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_prot = system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_fire = (system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_valid && system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_ready);
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_ready = (! system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rValid);
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_valid = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rValid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_addr = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_addr;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_id = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_id;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_region = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_region;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_len = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_len;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_size = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_size;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_burst = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_burst;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_lock = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_lock;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_cache = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_cache;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_qos = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_qos;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_prot = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_prot;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_valid = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_ready = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_ready;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_addr = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_id = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_region = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_region;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_len = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_len;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_size = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_size;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_burst = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_lock = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_cache = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_qos = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_prot = system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_ready = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_valid = (system_ddr_ddrLogic_userAdapters_0_userAxi4_w_valid || (! system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN));
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_data = (system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN ? system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_data : system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_data);
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_strb = (system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN ? system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_strb : system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_strb);
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_last = (system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN ? system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_last : system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_last);
  always @(*) begin
    system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_ready = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_34) begin
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_34 = (! system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rValid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_data = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_data;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_strb = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_strb;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_last = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_last;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_valid = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_ready;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_data = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_data;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_strb = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_strb;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_payload_last = system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_m2sPipe_payload_last;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_ready = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_valid = (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_valid || (! system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN));
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_data = (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_data : system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_data);
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_id = (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_id : system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_id);
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_resp = (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_resp : system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_resp);
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_last = (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_last : system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_last);
  always @(*) begin
    system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_ready = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_35) begin
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_35 = (! system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rValid;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_data = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_data;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_id = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_id;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_resp = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_resp;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_last = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_last;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_r_valid = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_0_userAxi4_r_ready;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_data = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_data;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_id = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_resp = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_resp;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_r_payload_last = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_m2sPipe_payload_last;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_fire = (system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_valid && system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_ready);
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_ready = (! system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rValid);
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_valid = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rValid;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_payload_id = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rData_id;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_payload_resp = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rData_resp;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_b_valid = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_ready = system_ddr_ddrLogic_userAdapters_0_userAxi4_b_ready;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_b_payload_id = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_0_userAxi4_b_payload_resp = system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_payload_resp;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_ready = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_ar_ready;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_valid = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_valid;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_data = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_data;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_last = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_last;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_id = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_id[3:0];
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_resp = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_r_payload_resp;
  assign system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_1_ar_payload_id = {2'd0, system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_ar_payload_id};
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_ready = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_aw_ready;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_w_ready = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_w_ready;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_valid = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_valid;
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_payload_id = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_payload_id[3:0];
  assign system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_payload_resp = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_b_payload_resp;
  assign system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_1_aw_payload_id = {2'd0, system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_aw_payload_id};
  assign io_ddrMasters_0_reset_read_buffer = ddrCd_logic_outputReset_buffercc_1_io_dataOut;
  assign io_ddrMasters_0_aw_ready = io_ddrMasters_0_aw_rValidN;
  assign io_ddrMasters_0_aw_s2mPipe_valid = (io_ddrMasters_0_aw_valid || (! io_ddrMasters_0_aw_rValidN));
  assign io_ddrMasters_0_aw_s2mPipe_payload_addr = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_addr : io_ddrMasters_0_aw_rData_addr);
  assign io_ddrMasters_0_aw_s2mPipe_payload_id = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_id : io_ddrMasters_0_aw_rData_id);
  assign io_ddrMasters_0_aw_s2mPipe_payload_region = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_region : io_ddrMasters_0_aw_rData_region);
  assign io_ddrMasters_0_aw_s2mPipe_payload_len = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_len : io_ddrMasters_0_aw_rData_len);
  assign io_ddrMasters_0_aw_s2mPipe_payload_size = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_size : io_ddrMasters_0_aw_rData_size);
  assign io_ddrMasters_0_aw_s2mPipe_payload_burst = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_burst : io_ddrMasters_0_aw_rData_burst);
  assign io_ddrMasters_0_aw_s2mPipe_payload_lock = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_lock : io_ddrMasters_0_aw_rData_lock);
  assign io_ddrMasters_0_aw_s2mPipe_payload_cache = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_cache : io_ddrMasters_0_aw_rData_cache);
  assign io_ddrMasters_0_aw_s2mPipe_payload_qos = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_qos : io_ddrMasters_0_aw_rData_qos);
  assign io_ddrMasters_0_aw_s2mPipe_payload_prot = (io_ddrMasters_0_aw_rValidN ? io_ddrMasters_0_aw_payload_prot : io_ddrMasters_0_aw_rData_prot);
  always @(*) begin
    io_ddrMasters_0_aw_s2mPipe_ready = io_ddrMasters_0_aw_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_36) begin
      io_ddrMasters_0_aw_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_36 = (! io_ddrMasters_0_aw_s2mPipe_m2sPipe_valid);
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_valid = io_ddrMasters_0_aw_s2mPipe_rValid;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_addr = io_ddrMasters_0_aw_s2mPipe_rData_addr;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_id = io_ddrMasters_0_aw_s2mPipe_rData_id;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_region = io_ddrMasters_0_aw_s2mPipe_rData_region;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_len = io_ddrMasters_0_aw_s2mPipe_rData_len;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_size = io_ddrMasters_0_aw_s2mPipe_rData_size;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_burst = io_ddrMasters_0_aw_s2mPipe_rData_burst;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_lock = io_ddrMasters_0_aw_s2mPipe_rData_lock;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_cache = io_ddrMasters_0_aw_s2mPipe_rData_cache;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_qos = io_ddrMasters_0_aw_s2mPipe_rData_qos;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_payload_prot = io_ddrMasters_0_aw_s2mPipe_rData_prot;
  assign io_ddrMasters_0_aw_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_1_bridge_io_input_aw_ready;
  assign io_ddrMasters_0_ar_halfPipe_fire = (io_ddrMasters_0_ar_halfPipe_valid && io_ddrMasters_0_ar_halfPipe_ready);
  assign io_ddrMasters_0_ar_ready = (! io_ddrMasters_0_ar_rValid);
  assign io_ddrMasters_0_ar_halfPipe_valid = io_ddrMasters_0_ar_rValid;
  assign io_ddrMasters_0_ar_halfPipe_payload_addr = io_ddrMasters_0_ar_rData_addr;
  assign io_ddrMasters_0_ar_halfPipe_payload_id = io_ddrMasters_0_ar_rData_id;
  assign io_ddrMasters_0_ar_halfPipe_payload_region = io_ddrMasters_0_ar_rData_region;
  assign io_ddrMasters_0_ar_halfPipe_payload_len = io_ddrMasters_0_ar_rData_len;
  assign io_ddrMasters_0_ar_halfPipe_payload_size = io_ddrMasters_0_ar_rData_size;
  assign io_ddrMasters_0_ar_halfPipe_payload_burst = io_ddrMasters_0_ar_rData_burst;
  assign io_ddrMasters_0_ar_halfPipe_payload_lock = io_ddrMasters_0_ar_rData_lock;
  assign io_ddrMasters_0_ar_halfPipe_payload_cache = io_ddrMasters_0_ar_rData_cache;
  assign io_ddrMasters_0_ar_halfPipe_payload_qos = io_ddrMasters_0_ar_rData_qos;
  assign io_ddrMasters_0_ar_halfPipe_payload_prot = io_ddrMasters_0_ar_rData_prot;
  assign io_ddrMasters_0_ar_halfPipe_ready = system_ddr_ddrLogic_userAdapters_1_bridge_io_input_ar_ready;
  assign io_ddrMasters_0_w_ready = io_ddrMasters_0_w_rValidN;
  assign io_ddrMasters_0_w_s2mPipe_valid = (io_ddrMasters_0_w_valid || (! io_ddrMasters_0_w_rValidN));
  assign io_ddrMasters_0_w_s2mPipe_payload_data = (io_ddrMasters_0_w_rValidN ? io_ddrMasters_0_w_payload_data : io_ddrMasters_0_w_rData_data);
  assign io_ddrMasters_0_w_s2mPipe_payload_strb = (io_ddrMasters_0_w_rValidN ? io_ddrMasters_0_w_payload_strb : io_ddrMasters_0_w_rData_strb);
  assign io_ddrMasters_0_w_s2mPipe_payload_last = (io_ddrMasters_0_w_rValidN ? io_ddrMasters_0_w_payload_last : io_ddrMasters_0_w_rData_last);
  always @(*) begin
    io_ddrMasters_0_w_s2mPipe_ready = io_ddrMasters_0_w_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_37) begin
      io_ddrMasters_0_w_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_37 = (! io_ddrMasters_0_w_s2mPipe_m2sPipe_valid);
  assign io_ddrMasters_0_w_s2mPipe_m2sPipe_valid = io_ddrMasters_0_w_s2mPipe_rValid;
  assign io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_data = io_ddrMasters_0_w_s2mPipe_rData_data;
  assign io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_strb = io_ddrMasters_0_w_s2mPipe_rData_strb;
  assign io_ddrMasters_0_w_s2mPipe_m2sPipe_payload_last = io_ddrMasters_0_w_s2mPipe_rData_last;
  assign io_ddrMasters_0_w_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_1_bridge_io_input_w_ready;
  always @(*) begin
    system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_ready = io_input_r_m2sPipe_ready_1;
    if(when_Stream_l375_38) begin
      system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_ready = 1'b1;
    end
  end

  assign when_Stream_l375_38 = (! io_input_r_m2sPipe_valid_1);
  assign io_input_r_m2sPipe_valid_1 = io_input_r_rValid_1;
  assign io_input_r_m2sPipe_payload_data_1 = io_input_r_rData_data_1;
  assign io_input_r_m2sPipe_payload_id_1 = io_input_r_rData_id_1;
  assign io_input_r_m2sPipe_payload_resp_1 = io_input_r_rData_resp_1;
  assign io_input_r_m2sPipe_payload_last_1 = io_input_r_rData_last_1;
  assign io_ddrMasters_0_r_valid = io_input_r_m2sPipe_valid_1;
  assign io_input_r_m2sPipe_ready_1 = io_ddrMasters_0_r_ready;
  assign io_ddrMasters_0_r_payload_data = io_input_r_m2sPipe_payload_data_1;
  assign io_ddrMasters_0_r_payload_id = io_input_r_m2sPipe_payload_id_1;
  assign io_ddrMasters_0_r_payload_resp = io_input_r_m2sPipe_payload_resp_1;
  assign io_ddrMasters_0_r_payload_last = io_input_r_m2sPipe_payload_last_1;
  assign io_input_b_s2mPipe_valid_1 = (system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_valid || (! io_input_b_rValidN_1));
  assign io_input_b_s2mPipe_payload_id_1 = (io_input_b_rValidN_1 ? system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_id : io_input_b_rData_id_1);
  assign io_input_b_s2mPipe_payload_resp_1 = (io_input_b_rValidN_1 ? system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_resp : io_input_b_rData_resp_1);
  always @(*) begin
    io_input_b_s2mPipe_ready_1 = io_input_b_s2mPipe_m2sPipe_ready_1;
    if(when_Stream_l375_39) begin
      io_input_b_s2mPipe_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_39 = (! io_input_b_s2mPipe_m2sPipe_valid_1);
  assign io_input_b_s2mPipe_m2sPipe_valid_1 = io_input_b_s2mPipe_rValid_1;
  assign io_input_b_s2mPipe_m2sPipe_payload_id_1 = io_input_b_s2mPipe_rData_id_1;
  assign io_input_b_s2mPipe_m2sPipe_payload_resp_1 = io_input_b_s2mPipe_rData_resp_1;
  assign io_ddrMasters_0_b_valid = io_input_b_s2mPipe_m2sPipe_valid_1;
  assign io_input_b_s2mPipe_m2sPipe_ready_1 = io_ddrMasters_0_b_ready;
  assign io_ddrMasters_0_b_payload_id = io_input_b_s2mPipe_m2sPipe_payload_id_1;
  assign io_ddrMasters_0_b_payload_resp = io_input_b_s2mPipe_m2sPipe_payload_resp_1;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_valid = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_valid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_addr = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_id = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_id;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_region = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_region;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_len = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_len;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_size = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_size;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_burst = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_lock = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_cache = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_qos = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_prot = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_ar_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_valid = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_valid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_addr = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_id = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_id;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_region = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_region;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_len = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_len;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_size = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_size;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_burst = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_lock = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_cache = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_qos = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_prot = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_aw_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_valid = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_valid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_data = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_data;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_strb = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_strb;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_last = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_w_payload_last;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_r_ready = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_r_ready;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_b_ready = system_ddr_ddrLogic_userAdapters_1_upsizer_logic_io_output_b_ready;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_fire = (system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_valid && system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_ready);
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_ready = (! system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rValid);
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_valid = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rValid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_addr = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_addr;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_id = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_id;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_region = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_region;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_len = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_len;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_size = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_size;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_burst = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_burst;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_lock = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_lock;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_cache = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_cache;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_qos = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_qos;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_prot = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_prot;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_valid = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_ready = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_ready;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_addr = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_id = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_region = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_region;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_len = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_len;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_size = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_size;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_burst = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_lock = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_cache = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_qos = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_prot = system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_fire = (system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_valid && system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_ready);
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_ready = (! system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rValid);
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_valid = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rValid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_addr = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_addr;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_id = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_id;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_region = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_region;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_len = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_len;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_size = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_size;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_burst = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_burst;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_lock = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_lock;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_cache = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_cache;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_qos = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_qos;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_prot = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_prot;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_valid = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_ready = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_ready;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_addr = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_addr;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_id = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_region = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_region;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_len = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_len;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_size = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_size;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_burst = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_burst;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_lock = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_lock;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_cache = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_cache;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_qos = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_qos;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_prot = system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_payload_prot;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_ready = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_valid = (system_ddr_ddrLogic_userAdapters_1_userAxi4_w_valid || (! system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN));
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_data = (system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN ? system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_data : system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_data);
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_strb = (system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN ? system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_strb : system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_strb);
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_last = (system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN ? system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_last : system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_last);
  always @(*) begin
    system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_ready = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_40) begin
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_40 = (! system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rValid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_data = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_data;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_strb = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_strb;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_last = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_last;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_valid = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_ready;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_data = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_data;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_strb = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_strb;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_payload_last = system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_m2sPipe_payload_last;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_ready = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_valid = (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_valid || (! system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN));
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_data = (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_data : system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_data);
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_id = (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_id : system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_id);
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_resp = (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_resp : system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_resp);
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_last = (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN ? system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_last : system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_last);
  always @(*) begin
    system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_ready = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_41) begin
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_41 = (! system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rValid;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_data = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_data;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_id = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_id;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_resp = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_resp;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_last = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_last;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_r_valid = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_userAdapters_1_userAxi4_r_ready;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_data = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_data;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_id = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_resp = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_resp;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_r_payload_last = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_m2sPipe_payload_last;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_fire = (system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_valid && system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_ready);
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_ready = (! system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rValid);
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_valid = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rValid;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_payload_id = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rData_id;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_payload_resp = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rData_resp;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_b_valid = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_valid;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_ready = system_ddr_ddrLogic_userAdapters_1_userAxi4_b_ready;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_b_payload_id = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_payload_id;
  assign system_ddr_ddrLogic_userAdapters_1_userAxi4_b_payload_resp = system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_payload_resp;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_ready = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_ar_ready;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_valid = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_valid;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_data = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_data;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_last = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_last;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_id = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_id[3:0];
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_resp = system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_r_payload_resp;
  assign system_ddr_ddrLogic_arbiterAxi4Read_io_inputs_2_ar_payload_id = {2'd0, system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_ar_payload_id};
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_ready = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_aw_ready;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_w_ready = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_w_ready;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_valid = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_valid;
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_payload_id = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_payload_id[3:0];
  assign system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_payload_resp = system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_b_payload_resp;
  assign system_ddr_ddrLogic_arbiterAxi4Write_io_inputs_2_aw_payload_id = {2'd0, system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_aw_payload_id};
  assign io_output_aw_s2mPipe_valid = (system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_valid || (! io_output_aw_rValidN));
  assign io_output_aw_s2mPipe_payload_addr = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_addr : io_output_aw_rData_addr);
  assign io_output_aw_s2mPipe_payload_id = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_id : io_output_aw_rData_id);
  assign io_output_aw_s2mPipe_payload_region = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_region : io_output_aw_rData_region);
  assign io_output_aw_s2mPipe_payload_len = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_len : io_output_aw_rData_len);
  assign io_output_aw_s2mPipe_payload_size = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_size : io_output_aw_rData_size);
  assign io_output_aw_s2mPipe_payload_burst = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_burst : io_output_aw_rData_burst);
  assign io_output_aw_s2mPipe_payload_lock = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_lock : io_output_aw_rData_lock);
  assign io_output_aw_s2mPipe_payload_cache = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_cache : io_output_aw_rData_cache);
  assign io_output_aw_s2mPipe_payload_qos = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_qos : io_output_aw_rData_qos);
  assign io_output_aw_s2mPipe_payload_prot = (io_output_aw_rValidN ? system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_prot : io_output_aw_rData_prot);
  always @(*) begin
    io_output_aw_s2mPipe_ready = io_output_aw_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_42) begin
      io_output_aw_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_42 = (! io_output_aw_s2mPipe_m2sPipe_valid);
  assign io_output_aw_s2mPipe_m2sPipe_valid = io_output_aw_s2mPipe_rValid;
  assign io_output_aw_s2mPipe_m2sPipe_payload_addr = io_output_aw_s2mPipe_rData_addr;
  assign io_output_aw_s2mPipe_m2sPipe_payload_id = io_output_aw_s2mPipe_rData_id;
  assign io_output_aw_s2mPipe_m2sPipe_payload_region = io_output_aw_s2mPipe_rData_region;
  assign io_output_aw_s2mPipe_m2sPipe_payload_len = io_output_aw_s2mPipe_rData_len;
  assign io_output_aw_s2mPipe_m2sPipe_payload_size = io_output_aw_s2mPipe_rData_size;
  assign io_output_aw_s2mPipe_m2sPipe_payload_burst = io_output_aw_s2mPipe_rData_burst;
  assign io_output_aw_s2mPipe_m2sPipe_payload_lock = io_output_aw_s2mPipe_rData_lock;
  assign io_output_aw_s2mPipe_m2sPipe_payload_cache = io_output_aw_s2mPipe_rData_cache;
  assign io_output_aw_s2mPipe_m2sPipe_payload_qos = io_output_aw_s2mPipe_rData_qos;
  assign io_output_aw_s2mPipe_m2sPipe_payload_prot = io_output_aw_s2mPipe_rData_prot;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_valid = io_output_aw_s2mPipe_m2sPipe_valid;
  assign io_output_aw_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_ddrAAxi4_aw_ready;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_addr = io_output_aw_s2mPipe_m2sPipe_payload_addr;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_id = io_output_aw_s2mPipe_m2sPipe_payload_id;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_region = io_output_aw_s2mPipe_m2sPipe_payload_region;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_len = io_output_aw_s2mPipe_m2sPipe_payload_len;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_size = io_output_aw_s2mPipe_m2sPipe_payload_size;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_burst = io_output_aw_s2mPipe_m2sPipe_payload_burst;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_lock = io_output_aw_s2mPipe_m2sPipe_payload_lock;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_cache = io_output_aw_s2mPipe_m2sPipe_payload_cache;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_qos = io_output_aw_s2mPipe_m2sPipe_payload_qos;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_payload_prot = io_output_aw_s2mPipe_m2sPipe_payload_prot;
  assign io_output_ar_s2mPipe_valid = (system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_valid || (! io_output_ar_rValidN));
  assign io_output_ar_s2mPipe_payload_addr = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_addr : io_output_ar_rData_addr);
  assign io_output_ar_s2mPipe_payload_id = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_id : io_output_ar_rData_id);
  assign io_output_ar_s2mPipe_payload_region = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_region : io_output_ar_rData_region);
  assign io_output_ar_s2mPipe_payload_len = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_len : io_output_ar_rData_len);
  assign io_output_ar_s2mPipe_payload_size = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_size : io_output_ar_rData_size);
  assign io_output_ar_s2mPipe_payload_burst = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_burst : io_output_ar_rData_burst);
  assign io_output_ar_s2mPipe_payload_lock = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_lock : io_output_ar_rData_lock);
  assign io_output_ar_s2mPipe_payload_cache = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_cache : io_output_ar_rData_cache);
  assign io_output_ar_s2mPipe_payload_qos = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_qos : io_output_ar_rData_qos);
  assign io_output_ar_s2mPipe_payload_prot = (io_output_ar_rValidN ? system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_prot : io_output_ar_rData_prot);
  always @(*) begin
    io_output_ar_s2mPipe_ready = io_output_ar_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_43) begin
      io_output_ar_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_43 = (! io_output_ar_s2mPipe_m2sPipe_valid);
  assign io_output_ar_s2mPipe_m2sPipe_valid = io_output_ar_s2mPipe_rValid;
  assign io_output_ar_s2mPipe_m2sPipe_payload_addr = io_output_ar_s2mPipe_rData_addr;
  assign io_output_ar_s2mPipe_m2sPipe_payload_id = io_output_ar_s2mPipe_rData_id;
  assign io_output_ar_s2mPipe_m2sPipe_payload_region = io_output_ar_s2mPipe_rData_region;
  assign io_output_ar_s2mPipe_m2sPipe_payload_len = io_output_ar_s2mPipe_rData_len;
  assign io_output_ar_s2mPipe_m2sPipe_payload_size = io_output_ar_s2mPipe_rData_size;
  assign io_output_ar_s2mPipe_m2sPipe_payload_burst = io_output_ar_s2mPipe_rData_burst;
  assign io_output_ar_s2mPipe_m2sPipe_payload_lock = io_output_ar_s2mPipe_rData_lock;
  assign io_output_ar_s2mPipe_m2sPipe_payload_cache = io_output_ar_s2mPipe_rData_cache;
  assign io_output_ar_s2mPipe_m2sPipe_payload_qos = io_output_ar_s2mPipe_rData_qos;
  assign io_output_ar_s2mPipe_m2sPipe_payload_prot = io_output_ar_s2mPipe_rData_prot;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_valid = io_output_ar_s2mPipe_m2sPipe_valid;
  assign io_output_ar_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_ddrAAxi4_ar_ready;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_addr = io_output_ar_s2mPipe_m2sPipe_payload_addr;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_id = io_output_ar_s2mPipe_m2sPipe_payload_id;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_region = io_output_ar_s2mPipe_m2sPipe_payload_region;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_len = io_output_ar_s2mPipe_m2sPipe_payload_len;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_size = io_output_ar_s2mPipe_m2sPipe_payload_size;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_burst = io_output_ar_s2mPipe_m2sPipe_payload_burst;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_lock = io_output_ar_s2mPipe_m2sPipe_payload_lock;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_cache = io_output_ar_s2mPipe_m2sPipe_payload_cache;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_qos = io_output_ar_s2mPipe_m2sPipe_payload_qos;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_payload_prot = io_output_ar_s2mPipe_m2sPipe_payload_prot;
  always @(*) begin
    system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_ready = io_output_w_m2sPipe_ready;
    if(when_Stream_l375_44) begin
      system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_ready = 1'b1;
    end
  end

  assign when_Stream_l375_44 = (! io_output_w_m2sPipe_valid);
  assign io_output_w_m2sPipe_valid = io_output_w_rValid;
  assign io_output_w_m2sPipe_payload_data = io_output_w_rData_data_1;
  assign io_output_w_m2sPipe_payload_strb = io_output_w_rData_strb_1;
  assign io_output_w_m2sPipe_payload_last = io_output_w_rData_last_1;
  always @(*) begin
    system_ddr_ddrLogic_ddrAAxi4_w_valid = io_output_w_m2sPipe_valid;
    if(when_TrionDdrGenerator_l363) begin
      system_ddr_ddrLogic_ddrAAxi4_w_valid = 1'b1;
    end
  end

  assign io_output_w_m2sPipe_ready = system_ddr_ddrLogic_ddrAAxi4_w_ready;
  assign system_ddr_ddrLogic_ddrAAxi4_w_payload_data = io_output_w_m2sPipe_payload_data;
  assign system_ddr_ddrLogic_ddrAAxi4_w_payload_strb = io_output_w_m2sPipe_payload_strb;
  always @(*) begin
    system_ddr_ddrLogic_ddrAAxi4_w_payload_last = io_output_w_m2sPipe_payload_last;
    if(when_TrionDdrGenerator_l363) begin
      system_ddr_ddrLogic_ddrAAxi4_w_payload_last = (system_ddr_ddrLogic_ddrAToAxi4_widStream_payload_len == system_ddr_ddrLogic_ddrAToAxi4_ddrA_wCounter);
    end
  end

  assign system_ddr_ddrLogic_ddrAAxi4_r_ready = system_ddr_ddrLogic_arbiterAxi4Read_io_output_r_ready;
  assign system_ddr_ddrLogic_ddrAAxi4_b_ready = system_ddr_ddrLogic_ddrAAxi4_b_rValidN;
  assign system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_valid = (system_ddr_ddrLogic_ddrAAxi4_b_valid || (! system_ddr_ddrLogic_ddrAAxi4_b_rValidN));
  assign system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_payload_id = (system_ddr_ddrLogic_ddrAAxi4_b_rValidN ? system_ddr_ddrLogic_ddrAAxi4_b_payload_id : system_ddr_ddrLogic_ddrAAxi4_b_rData_id);
  assign system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_payload_resp = (system_ddr_ddrLogic_ddrAAxi4_b_rValidN ? system_ddr_ddrLogic_ddrAAxi4_b_payload_resp : system_ddr_ddrLogic_ddrAAxi4_b_rData_resp);
  always @(*) begin
    system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_ready = system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_45) begin
      system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_45 = (! system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rValid;
  assign system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_payload_id = system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rData_id;
  assign system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_payload_resp = system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rData_resp;
  assign system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_arbiterAxi4Write_io_output_b_ready;
  always @(*) begin
    system_ddr_ddrLogic_ddrAReset_resetUnbuffered = 1'b0;
    if(when_TrionDdrGenerator_l257) begin
      system_ddr_ddrLogic_ddrAReset_resetUnbuffered = 1'b1;
    end
  end

  assign _zz_when_TrionDdrGenerator_l257[4 : 0] = 5'h1f;
  assign when_TrionDdrGenerator_l257 = (system_ddr_ddrLogic_ddrAReset_counter != _zz_when_TrionDdrGenerator_l257);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_addr = system_ddr_ddrLogic_ddrAAxi4_aw_payload_addr;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_id = system_ddr_ddrLogic_ddrAAxi4_aw_payload_id;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_region = system_ddr_ddrLogic_ddrAAxi4_aw_payload_region;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_len = system_ddr_ddrLogic_ddrAAxi4_aw_payload_len;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_size = system_ddr_ddrLogic_ddrAAxi4_aw_payload_size;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_burst = system_ddr_ddrLogic_ddrAAxi4_aw_payload_burst;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_lock = system_ddr_ddrLogic_ddrAAxi4_aw_payload_lock;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_cache = system_ddr_ddrLogic_ddrAAxi4_aw_payload_cache;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_qos = system_ddr_ddrLogic_ddrAAxi4_aw_payload_qos;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_prot = system_ddr_ddrLogic_ddrAAxi4_aw_payload_prot;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_addr = system_ddr_ddrLogic_ddrAAxi4_aw_payload_addr;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_id = system_ddr_ddrLogic_ddrAAxi4_aw_payload_id;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_region = system_ddr_ddrLogic_ddrAAxi4_aw_payload_region;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_len = system_ddr_ddrLogic_ddrAAxi4_aw_payload_len;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_size = system_ddr_ddrLogic_ddrAAxi4_aw_payload_size;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_burst = system_ddr_ddrLogic_ddrAAxi4_aw_payload_burst;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_lock = system_ddr_ddrLogic_ddrAAxi4_aw_payload_lock;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_cache = system_ddr_ddrLogic_ddrAAxi4_aw_payload_cache;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_qos = system_ddr_ddrLogic_ddrAAxi4_aw_payload_qos;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_prot = system_ddr_ddrLogic_ddrAAxi4_aw_payload_prot;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_fire = (system_ddr_ddrLogic_ddrAAxi4_aw_valid && system_ddr_ddrLogic_ddrAAxi4_aw_ready);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_valid = system_ddr_ddrLogic_ddrAAxi4_aw_fire;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_valid = system_ddr_ddrLogic_ddrAAxi4_aw_fire;
  assign system_ddr_ddrLogic_ddrAAxi4_aw_ready = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_ready && system_ddr_ddrLogic_ddrAToAxi4_patchAw_ready);
  assign system_ddr_ddrLogic_ddrAToAxi4_a2wPayload_len = system_ddr_ddrLogic_ddrAToAxi4_patchAw_payload_len;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_valid = system_ddr_ddrLogic_ddrAToAxi4_patchAw_valid;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_ready = system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_ready;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_payload_len = system_ddr_ddrLogic_ddrAToAxi4_a2wPayload_len;
  assign system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_ready = system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_push_ready;
  assign io_pop_s2mPipe_valid_2 = (system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_valid || (! io_pop_rValidN_2));
  assign io_pop_s2mPipe_payload_len = (io_pop_rValidN_2 ? system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_payload_len : io_pop_rData_len);
  always @(*) begin
    io_pop_s2mPipe_ready_2 = system_ddr_ddrLogic_ddrAToAxi4_widStream_ready;
    if(when_Stream_l375_46) begin
      io_pop_s2mPipe_ready_2 = 1'b1;
    end
  end

  assign when_Stream_l375_46 = (! system_ddr_ddrLogic_ddrAToAxi4_widStream_valid);
  assign system_ddr_ddrLogic_ddrAToAxi4_widStream_valid = io_pop_s2mPipe_rValid_2;
  assign system_ddr_ddrLogic_ddrAToAxi4_widStream_payload_len = io_pop_s2mPipe_rData_len;
  assign system_ddr_ddrLogic_ddrAAxi4_w_fire = (system_ddr_ddrLogic_ddrAAxi4_w_valid && system_ddr_ddrLogic_ddrAAxi4_w_ready);
  assign system_ddr_ddrLogic_ddrAToAxi4_widStream_ready = (system_ddr_ddrLogic_ddrAAxi4_w_fire && system_ddr_ddrLogic_ddrAAxi4_w_payload_last);
  assign when_TrionDdrGenerator_l363 = (ddrCd_logic_outputReset_regNext && system_ddr_ddrLogic_ddrAToAxi4_widStream_valid);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_ready = system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_valid = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_valid || (! system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN));
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_addr = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_addr : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_addr);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_id = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_id : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_id);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_region = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_region : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_region);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_len = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_len : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_len);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_size = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_size : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_size);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_burst = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_burst : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_burst);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_lock = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_lock : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_lock);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_cache = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_cache : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_cache);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_qos = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_qos : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_qos);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_prot = (system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN ? system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_prot : system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_prot);
  always @(*) begin
    system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_ready = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_47) begin
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_47 = (! system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rValid;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_addr = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_addr;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_id = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_id;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_region = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_region;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_len = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_len;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_size = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_size;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_burst = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_burst;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_lock = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_lock;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_cache = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_cache;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_qos = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_qos;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_prot = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_prot;
  assign io_ddrA_aw_valid = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_valid;
  assign system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_ready = io_ddrA_aw_ready;
  assign io_ddrA_aw_payload_addr = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_addr;
  assign io_ddrA_aw_payload_id = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_id;
  assign io_ddrA_aw_payload_region = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_region;
  assign io_ddrA_aw_payload_len = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_len;
  assign io_ddrA_aw_payload_size = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_size;
  assign io_ddrA_aw_payload_burst = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_burst;
  assign io_ddrA_aw_payload_lock = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_lock;
  assign io_ddrA_aw_payload_cache = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_cache;
  assign io_ddrA_aw_payload_qos = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_qos;
  assign io_ddrA_aw_payload_prot = system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_m2sPipe_payload_prot;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_ready = system_ddr_ddrLogic_ddrAAxi4_ar_rValidN;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_valid = (system_ddr_ddrLogic_ddrAAxi4_ar_valid || (! system_ddr_ddrLogic_ddrAAxi4_ar_rValidN));
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_addr = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_addr : system_ddr_ddrLogic_ddrAAxi4_ar_rData_addr);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_id = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_id : system_ddr_ddrLogic_ddrAAxi4_ar_rData_id);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_region = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_region : system_ddr_ddrLogic_ddrAAxi4_ar_rData_region);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_len = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_len : system_ddr_ddrLogic_ddrAAxi4_ar_rData_len);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_size = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_size : system_ddr_ddrLogic_ddrAAxi4_ar_rData_size);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_burst = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_burst : system_ddr_ddrLogic_ddrAAxi4_ar_rData_burst);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_lock = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_lock : system_ddr_ddrLogic_ddrAAxi4_ar_rData_lock);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_cache = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_cache : system_ddr_ddrLogic_ddrAAxi4_ar_rData_cache);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_qos = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_qos : system_ddr_ddrLogic_ddrAAxi4_ar_rData_qos);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_prot = (system_ddr_ddrLogic_ddrAAxi4_ar_rValidN ? system_ddr_ddrLogic_ddrAAxi4_ar_payload_prot : system_ddr_ddrLogic_ddrAAxi4_ar_rData_prot);
  always @(*) begin
    system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_ready = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_48) begin
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_48 = (! system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_valid);
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_valid = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rValid;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_addr = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_addr;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_id = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_id;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_region = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_region;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_len = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_len;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_size = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_size;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_burst = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_burst;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_lock = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_lock;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_cache = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_cache;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_qos = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_qos;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_prot = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_prot;
  assign io_ddrA_ar_valid = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_valid;
  assign system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_ready = io_ddrA_ar_ready;
  assign io_ddrA_ar_payload_addr = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_addr;
  assign io_ddrA_ar_payload_id = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_id;
  assign io_ddrA_ar_payload_region = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_region;
  assign io_ddrA_ar_payload_len = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_len;
  assign io_ddrA_ar_payload_size = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_size;
  assign io_ddrA_ar_payload_burst = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_burst;
  assign io_ddrA_ar_payload_lock = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_lock;
  assign io_ddrA_ar_payload_cache = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_cache;
  assign io_ddrA_ar_payload_qos = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_qos;
  assign io_ddrA_ar_payload_prot = system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_m2sPipe_payload_prot;
  assign _zz_io_ddrA_w_valid = (! (! system_ddr_ddrLogic_ddrAToAxi4_widStream_valid));
  assign system_ddr_ddrLogic_ddrAAxi4_w_ready = (io_ddrA_w_ready && _zz_io_ddrA_w_valid);
  assign io_ddrA_w_valid = (system_ddr_ddrLogic_ddrAAxi4_w_valid && _zz_io_ddrA_w_valid);
  assign io_ddrA_w_payload_data = system_ddr_ddrLogic_ddrAAxi4_w_payload_data;
  assign io_ddrA_w_payload_strb = system_ddr_ddrLogic_ddrAAxi4_w_payload_strb;
  assign io_ddrA_w_payload_last = system_ddr_ddrLogic_ddrAAxi4_w_payload_last;
  always @(*) begin
    io_ddrA_r_ready = io_ddrA_r_m2sPipe_ready;
    if(when_Stream_l375_49) begin
      io_ddrA_r_ready = 1'b1;
    end
    if(ddrCd_logic_outputReset_regNext_1) begin
      io_ddrA_r_ready = 1'b1;
    end
  end

  assign when_Stream_l375_49 = (! io_ddrA_r_m2sPipe_valid);
  assign io_ddrA_r_m2sPipe_valid = io_ddrA_r_rValid;
  assign io_ddrA_r_m2sPipe_payload_data = io_ddrA_r_rData_data;
  assign io_ddrA_r_m2sPipe_payload_id = io_ddrA_r_rData_id;
  assign io_ddrA_r_m2sPipe_payload_resp = io_ddrA_r_rData_resp;
  assign io_ddrA_r_m2sPipe_payload_last = io_ddrA_r_rData_last;
  assign system_ddr_ddrLogic_ddrAAxi4_r_valid = io_ddrA_r_m2sPipe_valid;
  assign io_ddrA_r_m2sPipe_ready = system_ddr_ddrLogic_ddrAAxi4_r_ready;
  assign system_ddr_ddrLogic_ddrAAxi4_r_payload_data = io_ddrA_r_m2sPipe_payload_data;
  assign system_ddr_ddrLogic_ddrAAxi4_r_payload_id = io_ddrA_r_m2sPipe_payload_id;
  assign system_ddr_ddrLogic_ddrAAxi4_r_payload_resp = io_ddrA_r_m2sPipe_payload_resp;
  assign system_ddr_ddrLogic_ddrAAxi4_r_payload_last = io_ddrA_r_m2sPipe_payload_last;
  always @(*) begin
    io_ddrA_b_ready = io_ddrA_b_rValidN;
    if(ddrCd_logic_outputReset_regNext_1) begin
      io_ddrA_b_ready = 1'b1;
    end
  end

  assign io_ddrA_b_s2mPipe_valid = (io_ddrA_b_valid || (! io_ddrA_b_rValidN));
  assign io_ddrA_b_s2mPipe_payload_id = (io_ddrA_b_rValidN ? io_ddrA_b_payload_id : io_ddrA_b_rData_id);
  assign io_ddrA_b_s2mPipe_payload_resp = (io_ddrA_b_rValidN ? io_ddrA_b_payload_resp : io_ddrA_b_rData_resp);
  always @(*) begin
    io_ddrA_b_s2mPipe_ready = io_ddrA_b_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_50) begin
      io_ddrA_b_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_50 = (! io_ddrA_b_s2mPipe_m2sPipe_valid);
  assign io_ddrA_b_s2mPipe_m2sPipe_valid = io_ddrA_b_s2mPipe_rValid;
  assign io_ddrA_b_s2mPipe_m2sPipe_payload_id = io_ddrA_b_s2mPipe_rData_id;
  assign io_ddrA_b_s2mPipe_m2sPipe_payload_resp = io_ddrA_b_s2mPipe_rData_resp;
  assign system_ddr_ddrLogic_ddrAAxi4_b_valid = io_ddrA_b_s2mPipe_m2sPipe_valid;
  assign io_ddrA_b_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_ddrAAxi4_b_ready;
  assign system_ddr_ddrLogic_ddrAAxi4_b_payload_id = io_ddrA_b_s2mPipe_m2sPipe_payload_id;
  assign system_ddr_ddrLogic_ddrAAxi4_b_payload_resp = io_ddrA_b_s2mPipe_m2sPipe_payload_resp;
  assign system_axiA_logic_bmbToAxiBridge_io_output_arw_ready = (system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_write ? system_axiA_logic_axiAAdapted_aw_ready : system_axiA_logic_axiAAdapted_ar_ready);
  assign system_axiA_logic_axiAAdapted_ar_valid = (system_axiA_logic_bmbToAxiBridge_io_output_arw_valid && (! system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_write));
  assign system_axiA_logic_axiAAdapted_ar_payload_addr = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_addr;
  assign system_axiA_logic_axiAAdapted_ar_payload_id = 8'h0;
  assign _zz_system_axiA_logic_axiAAdapted_ar_payload_region[3 : 0] = 4'b0000;
  assign system_axiA_logic_axiAAdapted_ar_payload_region = _zz_system_axiA_logic_axiAAdapted_ar_payload_region;
  assign system_axiA_logic_axiAAdapted_ar_payload_len = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_len;
  assign system_axiA_logic_axiAAdapted_ar_payload_size = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_size;
  assign system_axiA_logic_axiAAdapted_ar_payload_burst = 2'b01;
  assign system_axiA_logic_axiAAdapted_ar_payload_lock = 1'b0;
  assign system_axiA_logic_axiAAdapted_ar_payload_cache = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_cache;
  assign system_axiA_logic_axiAAdapted_ar_payload_qos = 4'b0000;
  assign system_axiA_logic_axiAAdapted_ar_payload_prot = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_prot;
  assign system_axiA_logic_axiAAdapted_aw_valid = (system_axiA_logic_bmbToAxiBridge_io_output_arw_valid && system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_write);
  assign system_axiA_logic_axiAAdapted_aw_payload_addr = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_addr;
  assign system_axiA_logic_axiAAdapted_aw_payload_id = 8'h0;
  assign _zz_system_axiA_logic_axiAAdapted_aw_payload_region[3 : 0] = 4'b0000;
  assign system_axiA_logic_axiAAdapted_aw_payload_region = _zz_system_axiA_logic_axiAAdapted_aw_payload_region;
  assign system_axiA_logic_axiAAdapted_aw_payload_len = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_len;
  assign system_axiA_logic_axiAAdapted_aw_payload_size = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_size;
  assign system_axiA_logic_axiAAdapted_aw_payload_burst = 2'b01;
  assign system_axiA_logic_axiAAdapted_aw_payload_lock = 1'b0;
  assign system_axiA_logic_axiAAdapted_aw_payload_cache = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_cache;
  assign system_axiA_logic_axiAAdapted_aw_payload_qos = 4'b0000;
  assign system_axiA_logic_axiAAdapted_aw_payload_prot = system_axiA_logic_bmbToAxiBridge_io_output_arw_payload_prot;
  assign system_axiA_logic_axiAAdapted_w_valid = system_axiA_logic_bmbToAxiBridge_io_output_w_valid;
  assign system_axiA_logic_axiAAdapted_w_payload_data = system_axiA_logic_bmbToAxiBridge_io_output_w_payload_data;
  assign system_axiA_logic_axiAAdapted_w_payload_strb = system_axiA_logic_bmbToAxiBridge_io_output_w_payload_strb;
  assign system_axiA_logic_axiAAdapted_w_payload_last = system_axiA_logic_bmbToAxiBridge_io_output_w_payload_last;
  assign system_axiA_logic_axiAAdapted_r_ready = system_axiA_logic_bmbToAxiBridge_io_output_r_ready;
  assign system_axiA_logic_axiAAdapted_b_ready = system_axiA_logic_bmbToAxiBridge_io_output_b_ready;
  assign axiA_arvalid = system_axiA_logic_axiAAdapted_ar_valid;
  assign system_axiA_logic_axiAAdapted_ar_ready = axiA_arready;
  assign axiA_araddr = system_axiA_logic_axiAAdapted_ar_payload_addr;
  assign axiA_arid = system_axiA_logic_axiAAdapted_ar_payload_id;
  assign axiA_arregion = system_axiA_logic_axiAAdapted_ar_payload_region;
  assign axiA_arlen = system_axiA_logic_axiAAdapted_ar_payload_len;
  assign axiA_arsize = system_axiA_logic_axiAAdapted_ar_payload_size;
  assign axiA_arburst = system_axiA_logic_axiAAdapted_ar_payload_burst;
  assign axiA_arlock = system_axiA_logic_axiAAdapted_ar_payload_lock;
  assign axiA_arcache = system_axiA_logic_axiAAdapted_ar_payload_cache;
  assign axiA_arqos = system_axiA_logic_axiAAdapted_ar_payload_qos;
  assign axiA_arprot = system_axiA_logic_axiAAdapted_ar_payload_prot;
  assign axiA_awvalid = system_axiA_logic_axiAAdapted_aw_valid;
  assign system_axiA_logic_axiAAdapted_aw_ready = axiA_awready;
  assign axiA_awaddr = system_axiA_logic_axiAAdapted_aw_payload_addr;
  assign axiA_awid = system_axiA_logic_axiAAdapted_aw_payload_id;
  assign axiA_awregion = system_axiA_logic_axiAAdapted_aw_payload_region;
  assign axiA_awlen = system_axiA_logic_axiAAdapted_aw_payload_len;
  assign axiA_awsize = system_axiA_logic_axiAAdapted_aw_payload_size;
  assign axiA_awburst = system_axiA_logic_axiAAdapted_aw_payload_burst;
  assign axiA_awlock = system_axiA_logic_axiAAdapted_aw_payload_lock;
  assign axiA_awcache = system_axiA_logic_axiAAdapted_aw_payload_cache;
  assign axiA_awqos = system_axiA_logic_axiAAdapted_aw_payload_qos;
  assign axiA_awprot = system_axiA_logic_axiAAdapted_aw_payload_prot;
  assign axiA_wvalid = system_axiA_logic_axiAAdapted_w_valid;
  assign system_axiA_logic_axiAAdapted_w_ready = axiA_wready;
  assign axiA_wdata = system_axiA_logic_axiAAdapted_w_payload_data;
  assign axiA_wstrb = system_axiA_logic_axiAAdapted_w_payload_strb;
  assign axiA_wlast = system_axiA_logic_axiAAdapted_w_payload_last;
  always @(*) begin
    axiA_rready = axiA_r_m2sPipe_ready;
    if(when_Stream_l375_51) begin
      axiA_rready = 1'b1;
    end
  end

  assign when_Stream_l375_51 = (! axiA_r_m2sPipe_valid);
  assign axiA_r_m2sPipe_valid = axiA_r_rValid;
  assign axiA_r_m2sPipe_payload_data = axiA_r_rData_data;
  assign axiA_r_m2sPipe_payload_id = axiA_r_rData_id;
  assign axiA_r_m2sPipe_payload_resp = axiA_r_rData_resp;
  assign axiA_r_m2sPipe_payload_last = axiA_r_rData_last;
  assign system_axiA_logic_axiAAdapted_r_valid = axiA_r_m2sPipe_valid;
  assign axiA_r_m2sPipe_ready = system_axiA_logic_axiAAdapted_r_ready;
  assign system_axiA_logic_axiAAdapted_r_payload_data = axiA_r_m2sPipe_payload_data;
  assign system_axiA_logic_axiAAdapted_r_payload_id = axiA_r_m2sPipe_payload_id;
  assign system_axiA_logic_axiAAdapted_r_payload_resp = axiA_r_m2sPipe_payload_resp;
  assign system_axiA_logic_axiAAdapted_r_payload_last = axiA_r_m2sPipe_payload_last;
  assign system_axiA_logic_axiAAdapted_b_valid = axiA_bvalid;
  assign axiA_bready = system_axiA_logic_axiAAdapted_b_ready;
  assign system_axiA_logic_axiAAdapted_b_payload_id = axiA_bid;
  assign system_axiA_logic_axiAAdapted_b_payload_resp = axiA_bresp;
  assign system_bridge_bmb_cmd_ready = system_bridge_bmb_cmd_rValidN;
  assign system_bridge_bmb_cmd_s2mPipe_valid = (system_bridge_bmb_cmd_valid || (! system_bridge_bmb_cmd_rValidN));
  assign system_bridge_bmb_cmd_s2mPipe_payload_last = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_last : system_bridge_bmb_cmd_rData_last);
  assign system_bridge_bmb_cmd_s2mPipe_payload_fragment_source = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_fragment_source : system_bridge_bmb_cmd_rData_fragment_source);
  assign system_bridge_bmb_cmd_s2mPipe_payload_fragment_opcode = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_fragment_opcode : system_bridge_bmb_cmd_rData_fragment_opcode);
  assign system_bridge_bmb_cmd_s2mPipe_payload_fragment_address = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_fragment_address : system_bridge_bmb_cmd_rData_fragment_address);
  assign system_bridge_bmb_cmd_s2mPipe_payload_fragment_length = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_fragment_length : system_bridge_bmb_cmd_rData_fragment_length);
  assign system_bridge_bmb_cmd_s2mPipe_payload_fragment_data = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_fragment_data : system_bridge_bmb_cmd_rData_fragment_data);
  assign system_bridge_bmb_cmd_s2mPipe_payload_fragment_mask = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_fragment_mask : system_bridge_bmb_cmd_rData_fragment_mask);
  assign system_bridge_bmb_cmd_s2mPipe_payload_fragment_context = (system_bridge_bmb_cmd_rValidN ? system_bridge_bmb_cmd_payload_fragment_context : system_bridge_bmb_cmd_rData_fragment_context);
  always @(*) begin
    system_bridge_bmb_cmd_s2mPipe_ready = system_bridge_bmb_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_52) begin
      system_bridge_bmb_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_52 = (! system_bridge_bmb_cmd_s2mPipe_m2sPipe_valid);
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_valid = system_bridge_bmb_cmd_s2mPipe_rValid;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_last = system_bridge_bmb_cmd_s2mPipe_rData_last;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_source = system_bridge_bmb_cmd_s2mPipe_rData_fragment_source;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_opcode = system_bridge_bmb_cmd_s2mPipe_rData_fragment_opcode;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_address = system_bridge_bmb_cmd_s2mPipe_rData_fragment_address;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_length = system_bridge_bmb_cmd_s2mPipe_rData_fragment_length;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_data = system_bridge_bmb_cmd_s2mPipe_rData_fragment_data;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_mask = system_bridge_bmb_cmd_s2mPipe_rData_fragment_mask;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_payload_fragment_context = system_bridge_bmb_cmd_s2mPipe_rData_fragment_context;
  assign system_bridge_bmb_cmd_s2mPipe_m2sPipe_ready = system_bridge_bmb_decoder_io_input_cmd_ready;
  assign system_bridge_bmb_rsp_valid = system_bridge_bmb_decoder_io_input_rsp_valid;
  assign system_bridge_bmb_rsp_payload_last = system_bridge_bmb_decoder_io_input_rsp_payload_last;
  assign system_bridge_bmb_rsp_payload_fragment_source = system_bridge_bmb_decoder_io_input_rsp_payload_fragment_source;
  assign system_bridge_bmb_rsp_payload_fragment_opcode = system_bridge_bmb_decoder_io_input_rsp_payload_fragment_opcode;
  assign system_bridge_bmb_rsp_payload_fragment_data = system_bridge_bmb_decoder_io_input_rsp_payload_fragment_data;
  assign system_bridge_bmb_rsp_payload_fragment_context = system_bridge_bmb_decoder_io_input_rsp_payload_fragment_context;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid || (! system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN));
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context = (system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context : system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context);
  always @(*) begin
    system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_53) begin
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_53 = (! system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid);
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready = system_ddr_ddrLogic_cc_fifo_io_input_cmd_ready;
  always @(*) begin
    _zz_io_input_rsp_ready_2 = system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
    if(when_Stream_l375_54) begin
      _zz_io_input_rsp_ready_2 = 1'b1;
    end
  end

  assign when_Stream_l375_54 = (! _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid);
  assign _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bridge_bmb_upSizer_io_output_cmd_valid;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bridge_bmb_upSizer_io_output_rsp_ready;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bridge_bmb_upSizer_io_output_cmd_payload_last;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source = system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_source;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_opcode;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_address;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_length;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_data;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_mask;
  assign system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bridge_bmb_upSizer_io_output_cmd_payload_fragment_context;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid || (! system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN));
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context = (system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN ? system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context : system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context);
  always @(*) begin
    system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_55) begin
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_55 = (! system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_valid = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_last = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_source = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_opcode = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_address = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_length = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_data = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_mask = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_payload_fragment_context = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_m2sPipe_ready = system_axiA_logic_bmbToAxiBridge_io_input_cmd_ready;
  assign _zz_io_input_rsp_ready_3 = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1;
  always @(*) begin
    _zz_2 = system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
    if(when_Stream_l375_56) begin
      _zz_2 = 1'b1;
    end
  end

  assign when_Stream_l375_56 = (! _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1);
  assign _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_2;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_3;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source_2;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode_2;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data_2;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context_2;
  assign _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_axiA_logic_bmbToAxiBridge_io_input_rsp_valid;
  assign _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_last;
  assign _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source = system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_source;
  assign _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_opcode;
  assign _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_data;
  assign _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_axiA_logic_bmbToAxiBridge_io_input_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_4 = (! system_axiA_interrupt_plic_gateway_waitCompletion);
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bridge_bmb_crossClock_io_output_cmd_valid;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bridge_bmb_crossClock_io_output_rsp_ready;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bridge_bmb_crossClock_io_output_cmd_payload_last;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source = system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_source;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_opcode;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_address;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_length;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_data;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_mask;
  assign system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bridge_bmb_crossClock_io_output_cmd_payload_fragment_context;
  assign system_bmbPeripheral_bmb_cmd_valid = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_bmbPeripheral_bmb_cmd_ready;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_bmbPeripheral_bmb_rsp_valid;
  assign system_bmbPeripheral_bmb_rsp_ready = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  assign system_bmbPeripheral_bmb_cmd_payload_last = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_bmbPeripheral_bmb_rsp_payload_last;
  assign system_bmbPeripheral_bmb_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_cmd_payload_fragment_address = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_cmd_payload_fragment_length = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_cmd_payload_fragment_data = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_cmd_payload_fragment_mask = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  assign system_bmbPeripheral_bmb_cmd_payload_fragment_context = system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_bmbPeripheral_bmb_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_bmbPeripheral_bmb_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_bmbPeripheral_bmb_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bridge_bmb_crossClock_1_io_output_cmd_valid;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bridge_bmb_crossClock_1_io_output_rsp_ready;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bridge_bmb_crossClock_1_io_output_cmd_payload_last;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_address[23:0];
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_mask;
  assign system_bmbPeripheral_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bridge_bmb_crossClock_1_io_output_cmd_payload_fragment_context;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_valid = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_ready;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_last = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_opcode = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_address = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_length = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_data = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_mask = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_payload_fragment_context = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_combStage_ready = system_ramA_logic_io_bus_cmd_ready;
  always @(*) begin
    _zz_io_bus_rsp_ready = system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
    if(when_Stream_l375_57) begin
      _zz_io_bus_rsp_ready = 1'b1;
    end
  end

  assign when_Stream_l375_57 = (! _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid);
  assign _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bridge_bmb_unburstify_1_io_output_cmd_valid;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bridge_bmb_unburstify_1_io_output_rsp_ready;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bridge_bmb_unburstify_1_io_output_cmd_payload_last;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_opcode;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_address[10:0];
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_length;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_data;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask = system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_mask;
  assign system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bridge_bmb_unburstify_1_io_output_cmd_payload_fragment_context;
  assign system_bmbPeripheral_bmb_cmd_combStage_valid = system_bmbPeripheral_bmb_cmd_valid;
  assign system_bmbPeripheral_bmb_cmd_ready = system_bmbPeripheral_bmb_cmd_combStage_ready;
  assign system_bmbPeripheral_bmb_cmd_combStage_payload_last = system_bmbPeripheral_bmb_cmd_payload_last;
  assign system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_opcode = system_bmbPeripheral_bmb_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_address = system_bmbPeripheral_bmb_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_length = system_bmbPeripheral_bmb_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_data = system_bmbPeripheral_bmb_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_mask = system_bmbPeripheral_bmb_cmd_payload_fragment_mask;
  assign system_bmbPeripheral_bmb_cmd_combStage_payload_fragment_context = system_bmbPeripheral_bmb_cmd_payload_fragment_context;
  assign system_bmbPeripheral_bmb_cmd_combStage_ready = system_bmbPeripheral_bmb_decoder_io_input_cmd_ready;
  assign _zz_io_input_rsp_ready_4 = (! _zz_system_bmbPeripheral_bmb_rsp_valid_1);
  assign _zz_system_bmbPeripheral_bmb_rsp_valid = _zz_system_bmbPeripheral_bmb_rsp_valid_1;
  assign system_bmbPeripheral_bmb_rsp_valid = _zz_system_bmbPeripheral_bmb_rsp_valid;
  assign system_bmbPeripheral_bmb_rsp_payload_last = _zz_system_bmbPeripheral_bmb_rsp_payload_last;
  assign system_bmbPeripheral_bmb_rsp_payload_fragment_opcode = _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_rsp_payload_fragment_data = _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_rsp_payload_fragment_context = _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_context;
  assign system_uart_0_io_txd = system_uart_0_io_logic_io_uart_txd;
  assign system_i2c_0_io_sda_write = system_i2c_0_io_logic_io_i2c_sda_write;
  assign system_i2c_0_io_scl_write = system_i2c_0_io_logic_io_i2c_scl_write;
  assign system_i2c_2_io_sda_write = system_i2c_2_io_logic_io_i2c_sda_write;
  assign system_i2c_2_io_scl_write = system_i2c_2_io_logic_io_i2c_scl_write;
  assign system_i2c_1_io_sda_write = system_i2c_1_io_logic_io_i2c_sda_write;
  assign system_i2c_1_io_scl_write = system_i2c_1_io_logic_io_i2c_scl_write;
  assign system_userTimer_1_interrupts_0 = system_userTimer_1_logic_io_interrupts[0];
  assign system_userTimer_0_interrupts_0 = system_userTimer_0_logic_io_interrupts[0];
  assign system_gpio_0_io_write = system_gpio_0_io_logic_io_gpio_write;
  assign system_gpio_0_io_writeEnable = system_gpio_0_io_logic_io_gpio_writeEnable;
  assign system_gpio_0_io_interrupts_0 = system_gpio_0_io_logic_io_interrupt[0];
  assign system_gpio_0_io_interrupts_1 = system_gpio_0_io_logic_io_interrupt[1];
  assign system_gpio_0_io_interrupts_2 = system_gpio_0_io_logic_io_interrupt[2];
  assign system_gpio_0_io_interrupts_3 = system_gpio_0_io_logic_io_interrupt[3];
  assign _zz_system_watchdog_logic_panics_0_plic_gateway_ip = system_watchdog_logic_logic_io_panics[0];
  assign io_apbSlave_2_PADDR = io_apbSlave_2_logic_io_output_PADDR;
  assign io_apbSlave_2_PSEL = io_apbSlave_2_logic_io_output_PSEL;
  assign io_apbSlave_2_PENABLE = io_apbSlave_2_logic_io_output_PENABLE;
  assign io_apbSlave_2_PWRITE = io_apbSlave_2_logic_io_output_PWRITE;
  assign io_apbSlave_2_PWDATA = io_apbSlave_2_logic_io_output_PWDATA;
  assign io_apbSlave_1_PADDR = io_apbSlave_1_logic_io_output_PADDR;
  assign io_apbSlave_1_PSEL = io_apbSlave_1_logic_io_output_PSEL;
  assign io_apbSlave_1_PENABLE = io_apbSlave_1_logic_io_output_PENABLE;
  assign io_apbSlave_1_PWRITE = io_apbSlave_1_logic_io_output_PWRITE;
  assign io_apbSlave_1_PWDATA = io_apbSlave_1_logic_io_output_PWDATA;
  assign io_apbSlave_4_PADDR = io_apbSlave_4_logic_io_output_PADDR;
  assign io_apbSlave_4_PSEL = io_apbSlave_4_logic_io_output_PSEL;
  assign io_apbSlave_4_PENABLE = io_apbSlave_4_logic_io_output_PENABLE;
  assign io_apbSlave_4_PWRITE = io_apbSlave_4_logic_io_output_PWRITE;
  assign io_apbSlave_4_PWDATA = io_apbSlave_4_logic_io_output_PWDATA;
  assign io_apbSlave_0_PADDR = io_apbSlave_0_logic_io_output_PADDR;
  assign io_apbSlave_0_PSEL = io_apbSlave_0_logic_io_output_PSEL;
  assign io_apbSlave_0_PENABLE = io_apbSlave_0_logic_io_output_PENABLE;
  assign io_apbSlave_0_PWRITE = io_apbSlave_0_logic_io_output_PWRITE;
  assign io_apbSlave_0_PWDATA = io_apbSlave_0_logic_io_output_PWDATA;
  assign io_apbSlave_3_PADDR = io_apbSlave_3_logic_io_output_PADDR;
  assign io_apbSlave_3_PSEL = io_apbSlave_3_logic_io_output_PSEL;
  assign io_apbSlave_3_PENABLE = io_apbSlave_3_logic_io_output_PENABLE;
  assign io_apbSlave_3_PWRITE = io_apbSlave_3_logic_io_output_PWRITE;
  assign io_apbSlave_3_PWDATA = io_apbSlave_3_logic_io_output_PWDATA;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_clint_logic_io_bus_cmd_ready;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_clint_logic_io_bus_rsp_valid;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_clint_logic_io_bus_rsp_payload_last;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_clint_logic_io_bus_rsp_payload_fragment_opcode;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_clint_logic_io_bus_rsp_payload_fragment_data;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_clint_logic_io_bus_rsp_payload_fragment_context;
  assign bufferCC_74_io_dataIn = system_clint_logic_io_timerInterrupt[0];
  assign bufferCC_75_io_dataIn = system_clint_logic_io_softwareInterrupt[0];
  assign bufferCC_76_io_dataIn = system_clint_logic_io_timerInterrupt[1];
  assign bufferCC_77_io_dataIn = system_clint_logic_io_softwareInterrupt[1];
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_uart_0_io_logic_io_bus_cmd_ready;
  assign _zz_io_bus_rsp_ready_1 = (! _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1);
  assign _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_5 = (! system_uart_0_io_interrupt_plic_gateway_waitCompletion);
  assign when_PlicGateway_l21_6 = (! system_spi_0_io_interrupt_plic_gateway_waitCompletion);
  assign system_spi_0_io_sclk_write = system_spi_0_io_logic_io_spi_sclk_write;
  assign system_spi_0_io_data_0_writeEnable = system_spi_0_io_logic_io_spi_data_0_writeEnable;
  assign system_spi_0_io_data_0_write = system_spi_0_io_logic_io_spi_data_0_write;
  assign system_spi_0_io_data_1_writeEnable = system_spi_0_io_logic_io_spi_data_1_writeEnable;
  assign system_spi_0_io_data_1_write = system_spi_0_io_logic_io_spi_data_1_write;
  assign system_spi_0_io_data_2_writeEnable = system_spi_0_io_logic_io_spi_data_2_writeEnable;
  assign system_spi_0_io_data_2_write = system_spi_0_io_logic_io_spi_data_2_write;
  assign system_spi_0_io_data_3_writeEnable = system_spi_0_io_logic_io_spi_data_3_writeEnable;
  assign system_spi_0_io_data_3_write = system_spi_0_io_logic_io_spi_data_3_write;
  assign system_spi_0_io_ss = system_spi_0_io_logic_io_spi_ss;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_spi_0_io_logic_io_ctrl_cmd_ready;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_spi_0_io_logic_io_ctrl_rsp_valid;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_spi_0_io_logic_io_ctrl_rsp_payload_last;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_data;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_spi_0_io_logic_io_ctrl_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_7 = (! system_spi_1_io_interrupt_plic_gateway_waitCompletion);
  assign system_spi_1_io_sclk_write = system_spi_1_io_logic_io_spi_sclk_write;
  assign system_spi_1_io_data_0_writeEnable = system_spi_1_io_logic_io_spi_data_0_writeEnable;
  assign system_spi_1_io_data_0_write = system_spi_1_io_logic_io_spi_data_0_write;
  assign system_spi_1_io_data_1_writeEnable = system_spi_1_io_logic_io_spi_data_1_writeEnable;
  assign system_spi_1_io_data_1_write = system_spi_1_io_logic_io_spi_data_1_write;
  assign system_spi_1_io_data_2_writeEnable = system_spi_1_io_logic_io_spi_data_2_writeEnable;
  assign system_spi_1_io_data_2_write = system_spi_1_io_logic_io_spi_data_2_write;
  assign system_spi_1_io_data_3_writeEnable = system_spi_1_io_logic_io_spi_data_3_writeEnable;
  assign system_spi_1_io_data_3_write = system_spi_1_io_logic_io_spi_data_3_write;
  assign system_spi_1_io_ss = system_spi_1_io_logic_io_spi_ss;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_spi_1_io_logic_io_ctrl_cmd_ready;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_spi_1_io_logic_io_ctrl_rsp_valid;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_spi_1_io_logic_io_ctrl_rsp_payload_last;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_data;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_spi_1_io_logic_io_ctrl_rsp_payload_fragment_context;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_i2c_0_io_logic_io_ctrl_cmd_ready;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_i2c_0_io_logic_io_ctrl_rsp_valid;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_i2c_0_io_logic_io_ctrl_rsp_payload_last;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_data;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_i2c_0_io_logic_io_ctrl_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_8 = (! system_i2c_0_io_interrupt_plic_gateway_waitCompletion);
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_i2c_2_io_logic_io_ctrl_cmd_ready;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_i2c_2_io_logic_io_ctrl_rsp_valid;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_i2c_2_io_logic_io_ctrl_rsp_payload_last;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_data;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_i2c_2_io_logic_io_ctrl_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_9 = (! system_i2c_2_io_interrupt_plic_gateway_waitCompletion);
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_i2c_1_io_logic_io_ctrl_cmd_ready;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_i2c_1_io_logic_io_ctrl_rsp_valid;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_i2c_1_io_logic_io_ctrl_rsp_payload_last;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_opcode;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_data;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_i2c_1_io_logic_io_ctrl_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_10 = (! system_i2c_1_io_interrupt_plic_gateway_waitCompletion);
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_userTimer_1_logic_io_ctrl_cmd_ready;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_userTimer_1_logic_io_ctrl_rsp_valid;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_userTimer_1_logic_io_ctrl_rsp_payload_last;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_opcode;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_data;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_userTimer_1_logic_io_ctrl_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_11 = (! system_userTimer_1_interrupts_0_plic_gateway_waitCompletion);
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire = (system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid && system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready);
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = (! system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid);
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_valid = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_last = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_opcode = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_address = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_length = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_data = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_payload_fragment_context = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_ready = system_userTimer_0_logic_io_ctrl_cmd_ready;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_userTimer_0_logic_io_ctrl_rsp_valid;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_userTimer_0_logic_io_ctrl_rsp_payload_last;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_opcode;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_data;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_userTimer_0_logic_io_ctrl_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_12 = (! system_userTimer_0_interrupts_0_plic_gateway_waitCompletion);
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_gpio_0_io_logic_io_bus_cmd_ready;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_gpio_0_io_logic_io_bus_rsp_valid;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_gpio_0_io_logic_io_bus_rsp_payload_last;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_gpio_0_io_logic_io_bus_rsp_payload_fragment_opcode;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_gpio_0_io_logic_io_bus_rsp_payload_fragment_data;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_gpio_0_io_logic_io_bus_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_13 = (! system_gpio_0_io_interrupts_0_plic_gateway_waitCompletion);
  assign when_PlicGateway_l21_14 = (! system_gpio_0_io_interrupts_1_plic_gateway_waitCompletion);
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_watchdog_logic_logic_io_bus_cmd_ready;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_watchdog_logic_logic_io_bus_rsp_valid;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_watchdog_logic_logic_io_bus_rsp_payload_last;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_watchdog_logic_logic_io_bus_rsp_payload_fragment_opcode;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_watchdog_logic_logic_io_bus_rsp_payload_fragment_data;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_watchdog_logic_logic_io_bus_rsp_payload_fragment_context;
  assign when_PlicGateway_l21_15 = (! system_watchdog_logic_panics_0_plic_gateway_waitCompletion);
  assign system_watchdog_hardPanic = system_watchdog_logic_logic_io_panics[1];
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = io_apbSlave_2_logic_io_input_cmd_ready;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = io_apbSlave_2_logic_io_input_rsp_valid;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = io_apbSlave_2_logic_io_input_rsp_payload_last;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = io_apbSlave_2_logic_io_input_rsp_payload_fragment_opcode;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = io_apbSlave_2_logic_io_input_rsp_payload_fragment_data;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = io_apbSlave_2_logic_io_input_rsp_payload_fragment_context;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = io_apbSlave_1_logic_io_input_cmd_ready;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = io_apbSlave_1_logic_io_input_rsp_valid;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = io_apbSlave_1_logic_io_input_rsp_payload_last;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = io_apbSlave_1_logic_io_input_rsp_payload_fragment_opcode;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = io_apbSlave_1_logic_io_input_rsp_payload_fragment_data;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = io_apbSlave_1_logic_io_input_rsp_payload_fragment_context;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = io_apbSlave_4_logic_io_input_cmd_ready;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = io_apbSlave_4_logic_io_input_rsp_valid;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = io_apbSlave_4_logic_io_input_rsp_payload_last;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = io_apbSlave_4_logic_io_input_rsp_payload_fragment_opcode;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = io_apbSlave_4_logic_io_input_rsp_payload_fragment_data;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = io_apbSlave_4_logic_io_input_rsp_payload_fragment_context;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = io_apbSlave_0_logic_io_input_cmd_ready;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = io_apbSlave_0_logic_io_input_rsp_valid;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = io_apbSlave_0_logic_io_input_rsp_payload_last;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = io_apbSlave_0_logic_io_input_rsp_payload_fragment_opcode;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = io_apbSlave_0_logic_io_input_rsp_payload_fragment_data;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = io_apbSlave_0_logic_io_input_rsp_payload_fragment_context;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = io_apbSlave_3_logic_io_input_cmd_ready;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = io_apbSlave_3_logic_io_input_rsp_valid;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = io_apbSlave_3_logic_io_input_rsp_payload_last;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = io_apbSlave_3_logic_io_input_rsp_payload_fragment_opcode;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = io_apbSlave_3_logic_io_input_rsp_payload_fragment_data;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = io_apbSlave_3_logic_io_input_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid = system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready = system_bmbPeripheral_bmb_decoder_io_outputs_1_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last = system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address = system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length = system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data = system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context = system_bmbPeripheral_bmb_decoder_io_outputs_1_cmd_payload_fragment_context;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready = system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid = system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last = system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address[15:0];
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data;
  assign system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode = system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data = system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context = system_clint_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_1 = system_bmbPeripheral_bmb_decoder_io_outputs_2_cmd_payload_fragment_context;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_1;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_1 = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_1 = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_1;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_1;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_1 = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_1;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_1[5:0];
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_1;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_1;
  assign system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_1;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_1 = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_1 = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_1 = system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_2 = system_bmbPeripheral_bmb_decoder_io_outputs_3_cmd_payload_fragment_context;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_2;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_2 = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_2 = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_2;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_2;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_2 = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_2;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_2[11:0];
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_2;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_2;
  assign system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_2;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_2 = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_2 = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_2 = system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_3 = system_bmbPeripheral_bmb_decoder_io_outputs_4_cmd_payload_fragment_context;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_3;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_3 = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_3 = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_3;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_3;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_3 = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_3;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_3[11:0];
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_3;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_3;
  assign system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_3;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_3 = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_3 = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_3 = system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_4 = system_bmbPeripheral_bmb_decoder_io_outputs_5_cmd_payload_fragment_context;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_4;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_4 = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_4 = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_4;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_4;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_4 = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_4;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_4[7:0];
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_4;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_4;
  assign system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_4;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_4 = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_4 = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_4 = system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_5 = system_bmbPeripheral_bmb_decoder_io_outputs_6_cmd_payload_fragment_context;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_5;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_5 = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_5 = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_5;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_5;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_5 = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_5;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_5[7:0];
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_5;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_5;
  assign system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_5;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_5 = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_5 = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_5 = system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_6 = system_bmbPeripheral_bmb_decoder_io_outputs_7_cmd_payload_fragment_context;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_6;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_6 = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_6 = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_6;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_6;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_6 = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_6;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_6[7:0];
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_6;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_6;
  assign system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_6;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_6 = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_6 = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_6 = system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_7 = system_bmbPeripheral_bmb_decoder_io_outputs_8_cmd_payload_fragment_context;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_7;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_7 = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_7 = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_7;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_7;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_7 = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_7;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_7[7:0];
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_7;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_7;
  assign system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_7;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_7 = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_7 = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_7 = system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_8 = system_bmbPeripheral_bmb_decoder_io_outputs_9_cmd_payload_fragment_context;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_8;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_8 = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_8 = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_8;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_8;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_8 = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_8;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_8[7:0];
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_8;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_8;
  assign system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_8;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_8 = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_8 = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_8 = system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_9 = system_bmbPeripheral_bmb_decoder_io_outputs_10_cmd_payload_fragment_context;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_9;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_9 = system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_9 = system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_9;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_9;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_9 = system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_9;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_9[7:0];
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_9;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_9;
  assign system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_9;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_9 = system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_9 = system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_9 = system_gpio_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_10 = system_bmbPeripheral_bmb_decoder_io_outputs_11_cmd_payload_fragment_context;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_10;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_10 = system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_10 = system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_10;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_10;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_10 = system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_10;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_10[7:0];
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_10;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_10;
  assign system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_10;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_10 = system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_10 = system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_10 = system_watchdog_logic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_plic_logic_bus_readErrorFlag = 1'b0;
  assign system_plic_logic_bus_writeErrorFlag = 1'b0;
  always @(*) begin
    system_plic_logic_bus_readHaltTrigger = 1'b0;
    if(when_PlicMapper_l122) begin
      system_plic_logic_bus_readHaltTrigger = 1'b1;
    end
  end

  assign system_plic_logic_bus_writeHaltTrigger = 1'b0;
  assign _zz_system_plic_logic_bus_rsp_ready = (! (system_plic_logic_bus_readHaltTrigger || system_plic_logic_bus_writeHaltTrigger));
  assign system_plic_logic_bus_rsp_ready = (_zz_system_plic_logic_bus_rsp_ready_1 && _zz_system_plic_logic_bus_rsp_ready);
  always @(*) begin
    _zz_system_plic_logic_bus_rsp_ready_1 = system_plic_logic_bmb_rsp_ready;
    if(when_Stream_l375_58) begin
      _zz_system_plic_logic_bus_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375_58 = (! _zz_system_plic_logic_bmb_rsp_valid);
  assign _zz_system_plic_logic_bmb_rsp_valid = _zz_system_plic_logic_bmb_rsp_valid_1;
  assign system_plic_logic_bmb_rsp_valid = _zz_system_plic_logic_bmb_rsp_valid;
  assign system_plic_logic_bmb_rsp_payload_last = _zz_system_plic_logic_bmb_rsp_payload_last;
  assign system_plic_logic_bmb_rsp_payload_fragment_opcode = _zz_system_plic_logic_bmb_rsp_payload_fragment_opcode;
  assign system_plic_logic_bmb_rsp_payload_fragment_data = _zz_system_plic_logic_bmb_rsp_payload_fragment_data;
  assign system_plic_logic_bmb_rsp_payload_fragment_context = _zz_system_plic_logic_bmb_rsp_payload_fragment_context;
  assign system_plic_logic_bus_askWrite = (system_plic_logic_bmb_cmd_valid && (system_plic_logic_bmb_cmd_payload_fragment_opcode == 1'b1));
  assign system_plic_logic_bus_askRead = (system_plic_logic_bmb_cmd_valid && (system_plic_logic_bmb_cmd_payload_fragment_opcode == 1'b0));
  assign system_plic_logic_bmb_cmd_fire = (system_plic_logic_bmb_cmd_valid && system_plic_logic_bmb_cmd_ready);
  assign system_plic_logic_bus_doWrite = (system_plic_logic_bmb_cmd_fire && (system_plic_logic_bmb_cmd_payload_fragment_opcode == 1'b1));
  assign system_plic_logic_bus_doRead = (system_plic_logic_bmb_cmd_fire && (system_plic_logic_bmb_cmd_payload_fragment_opcode == 1'b0));
  assign system_plic_logic_bus_rsp_valid = system_plic_logic_bmb_cmd_valid;
  assign system_plic_logic_bmb_cmd_ready = system_plic_logic_bus_rsp_ready;
  assign system_plic_logic_bus_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (system_plic_logic_bus_doWrite && system_plic_logic_bus_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      system_plic_logic_bus_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        system_plic_logic_bus_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        system_plic_logic_bus_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (system_plic_logic_bus_doRead && system_plic_logic_bus_readErrorFlag);
  always @(*) begin
    system_plic_logic_bus_rsp_payload_fragment_data = 32'h0;
    case(system_plic_logic_bmb_cmd_payload_fragment_address)
      22'h000040 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = userInterruptA_interrupt_plic_gateway_priority;
      end
      22'h001000 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[16 : 16] = userInterruptA_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[23 : 23] = userInterruptD_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[22 : 22] = userInterruptC_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[17 : 17] = userInterruptB_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[30 : 30] = system_axiA_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 1] = system_uart_0_io_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[4 : 4] = system_spi_0_io_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[5 : 5] = system_spi_1_io_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[8 : 8] = system_i2c_0_io_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[10 : 10] = system_i2c_2_io_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[9 : 9] = system_i2c_1_io_interrupt_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[20 : 20] = system_userTimer_1_interrupts_0_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[19 : 19] = system_userTimer_0_interrupts_0_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[12 : 12] = system_gpio_0_io_interrupts_0_plic_gateway_ip;
        system_plic_logic_bus_rsp_payload_fragment_data[13 : 13] = system_gpio_0_io_interrupts_1_plic_gateway_ip;
      end
      22'h00005c : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = userInterruptD_interrupt_plic_gateway_priority;
      end
      22'h000058 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = userInterruptC_interrupt_plic_gateway_priority;
      end
      22'h000044 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = userInterruptB_interrupt_plic_gateway_priority;
      end
      22'h000078 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_axiA_interrupt_plic_gateway_priority;
      end
      22'h000004 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_uart_0_io_interrupt_plic_gateway_priority;
      end
      22'h000010 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_spi_0_io_interrupt_plic_gateway_priority;
      end
      22'h000014 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_spi_1_io_interrupt_plic_gateway_priority;
      end
      22'h000020 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_i2c_0_io_interrupt_plic_gateway_priority;
      end
      22'h000028 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_i2c_2_io_interrupt_plic_gateway_priority;
      end
      22'h000024 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_i2c_1_io_interrupt_plic_gateway_priority;
      end
      22'h000050 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_userTimer_1_interrupts_0_plic_gateway_priority;
      end
      22'h00004c : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_userTimer_0_interrupts_0_plic_gateway_priority;
      end
      22'h000030 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_gpio_0_io_interrupts_0_plic_gateway_priority;
      end
      22'h000034 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_gpio_0_io_interrupts_1_plic_gateway_priority;
      end
      22'h000080 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_watchdog_logic_panics_0_plic_gateway_priority;
      end
      22'h001004 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[0 : 0] = system_watchdog_logic_panics_0_plic_gateway_ip;
      end
      22'h200000 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_cores_0_externalInterrupt_plic_target_threshold;
      end
      22'h200004 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[5 : 0] = system_cores_0_externalInterrupt_plic_target_claim;
      end
      22'h002000 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[16 : 16] = system_cores_0_externalInterrupt_plic_target_ie_0;
        system_plic_logic_bus_rsp_payload_fragment_data[23 : 23] = system_cores_0_externalInterrupt_plic_target_ie_1;
        system_plic_logic_bus_rsp_payload_fragment_data[22 : 22] = system_cores_0_externalInterrupt_plic_target_ie_2;
        system_plic_logic_bus_rsp_payload_fragment_data[17 : 17] = system_cores_0_externalInterrupt_plic_target_ie_3;
        system_plic_logic_bus_rsp_payload_fragment_data[30 : 30] = system_cores_0_externalInterrupt_plic_target_ie_4;
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 1] = system_cores_0_externalInterrupt_plic_target_ie_5;
        system_plic_logic_bus_rsp_payload_fragment_data[4 : 4] = system_cores_0_externalInterrupt_plic_target_ie_6;
        system_plic_logic_bus_rsp_payload_fragment_data[5 : 5] = system_cores_0_externalInterrupt_plic_target_ie_7;
        system_plic_logic_bus_rsp_payload_fragment_data[8 : 8] = system_cores_0_externalInterrupt_plic_target_ie_8;
        system_plic_logic_bus_rsp_payload_fragment_data[10 : 10] = system_cores_0_externalInterrupt_plic_target_ie_9;
        system_plic_logic_bus_rsp_payload_fragment_data[9 : 9] = system_cores_0_externalInterrupt_plic_target_ie_10;
        system_plic_logic_bus_rsp_payload_fragment_data[20 : 20] = system_cores_0_externalInterrupt_plic_target_ie_11;
        system_plic_logic_bus_rsp_payload_fragment_data[19 : 19] = system_cores_0_externalInterrupt_plic_target_ie_12;
        system_plic_logic_bus_rsp_payload_fragment_data[12 : 12] = system_cores_0_externalInterrupt_plic_target_ie_13;
        system_plic_logic_bus_rsp_payload_fragment_data[13 : 13] = system_cores_0_externalInterrupt_plic_target_ie_14;
      end
      22'h002004 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[0 : 0] = system_cores_0_externalInterrupt_plic_target_ie_15;
      end
      22'h201000 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 0] = system_cores_1_externalInterrupt_plic_target_threshold;
      end
      22'h201004 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[5 : 0] = system_cores_1_externalInterrupt_plic_target_claim;
      end
      22'h002080 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[16 : 16] = system_cores_1_externalInterrupt_plic_target_ie_0;
        system_plic_logic_bus_rsp_payload_fragment_data[23 : 23] = system_cores_1_externalInterrupt_plic_target_ie_1;
        system_plic_logic_bus_rsp_payload_fragment_data[22 : 22] = system_cores_1_externalInterrupt_plic_target_ie_2;
        system_plic_logic_bus_rsp_payload_fragment_data[17 : 17] = system_cores_1_externalInterrupt_plic_target_ie_3;
        system_plic_logic_bus_rsp_payload_fragment_data[30 : 30] = system_cores_1_externalInterrupt_plic_target_ie_4;
        system_plic_logic_bus_rsp_payload_fragment_data[1 : 1] = system_cores_1_externalInterrupt_plic_target_ie_5;
        system_plic_logic_bus_rsp_payload_fragment_data[4 : 4] = system_cores_1_externalInterrupt_plic_target_ie_6;
        system_plic_logic_bus_rsp_payload_fragment_data[5 : 5] = system_cores_1_externalInterrupt_plic_target_ie_7;
        system_plic_logic_bus_rsp_payload_fragment_data[8 : 8] = system_cores_1_externalInterrupt_plic_target_ie_8;
        system_plic_logic_bus_rsp_payload_fragment_data[10 : 10] = system_cores_1_externalInterrupt_plic_target_ie_9;
        system_plic_logic_bus_rsp_payload_fragment_data[9 : 9] = system_cores_1_externalInterrupt_plic_target_ie_10;
        system_plic_logic_bus_rsp_payload_fragment_data[20 : 20] = system_cores_1_externalInterrupt_plic_target_ie_11;
        system_plic_logic_bus_rsp_payload_fragment_data[19 : 19] = system_cores_1_externalInterrupt_plic_target_ie_12;
        system_plic_logic_bus_rsp_payload_fragment_data[12 : 12] = system_cores_1_externalInterrupt_plic_target_ie_13;
        system_plic_logic_bus_rsp_payload_fragment_data[13 : 13] = system_cores_1_externalInterrupt_plic_target_ie_14;
      end
      22'h002084 : begin
        system_plic_logic_bus_rsp_payload_fragment_data[0 : 0] = system_cores_1_externalInterrupt_plic_target_ie_15;
      end
      default : begin
      end
    endcase
  end

  assign system_plic_logic_bus_rsp_payload_fragment_context = system_plic_logic_bmb_cmd_payload_fragment_context;
  assign system_cores_0_externalInterrupt_plic_target_requests_0_priority = 2'b00;
  assign system_cores_0_externalInterrupt_plic_target_requests_0_id = 6'h0;
  assign system_cores_0_externalInterrupt_plic_target_requests_0_valid = 1'b1;
  assign system_cores_0_externalInterrupt_plic_target_requests_1_priority = system_uart_0_io_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_1_id = 6'h01;
  assign system_cores_0_externalInterrupt_plic_target_requests_1_valid = (system_uart_0_io_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_5);
  assign system_cores_0_externalInterrupt_plic_target_requests_2_priority = system_spi_0_io_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_2_id = 6'h04;
  assign system_cores_0_externalInterrupt_plic_target_requests_2_valid = (system_spi_0_io_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_6);
  assign system_cores_0_externalInterrupt_plic_target_requests_3_priority = system_spi_1_io_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_3_id = 6'h05;
  assign system_cores_0_externalInterrupt_plic_target_requests_3_valid = (system_spi_1_io_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_7);
  assign system_cores_0_externalInterrupt_plic_target_requests_4_priority = system_i2c_0_io_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_4_id = 6'h08;
  assign system_cores_0_externalInterrupt_plic_target_requests_4_valid = (system_i2c_0_io_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_8);
  assign system_cores_0_externalInterrupt_plic_target_requests_5_priority = system_i2c_1_io_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_5_id = 6'h09;
  assign system_cores_0_externalInterrupt_plic_target_requests_5_valid = (system_i2c_1_io_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_10);
  assign system_cores_0_externalInterrupt_plic_target_requests_6_priority = system_i2c_2_io_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_6_id = 6'h0a;
  assign system_cores_0_externalInterrupt_plic_target_requests_6_valid = (system_i2c_2_io_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_9);
  assign system_cores_0_externalInterrupt_plic_target_requests_7_priority = system_gpio_0_io_interrupts_0_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_7_id = 6'h0c;
  assign system_cores_0_externalInterrupt_plic_target_requests_7_valid = (system_gpio_0_io_interrupts_0_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_13);
  assign system_cores_0_externalInterrupt_plic_target_requests_8_priority = system_gpio_0_io_interrupts_1_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_8_id = 6'h0d;
  assign system_cores_0_externalInterrupt_plic_target_requests_8_valid = (system_gpio_0_io_interrupts_1_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_14);
  assign system_cores_0_externalInterrupt_plic_target_requests_9_priority = userInterruptA_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_9_id = 6'h10;
  assign system_cores_0_externalInterrupt_plic_target_requests_9_valid = (userInterruptA_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_0);
  assign system_cores_0_externalInterrupt_plic_target_requests_10_priority = userInterruptB_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_10_id = 6'h11;
  assign system_cores_0_externalInterrupt_plic_target_requests_10_valid = (userInterruptB_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_3);
  assign system_cores_0_externalInterrupt_plic_target_requests_11_priority = system_userTimer_0_interrupts_0_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_11_id = 6'h13;
  assign system_cores_0_externalInterrupt_plic_target_requests_11_valid = (system_userTimer_0_interrupts_0_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_12);
  assign system_cores_0_externalInterrupt_plic_target_requests_12_priority = system_userTimer_1_interrupts_0_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_12_id = 6'h14;
  assign system_cores_0_externalInterrupt_plic_target_requests_12_valid = (system_userTimer_1_interrupts_0_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_11);
  assign system_cores_0_externalInterrupt_plic_target_requests_13_priority = userInterruptC_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_13_id = 6'h16;
  assign system_cores_0_externalInterrupt_plic_target_requests_13_valid = (userInterruptC_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_2);
  assign system_cores_0_externalInterrupt_plic_target_requests_14_priority = userInterruptD_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_14_id = 6'h17;
  assign system_cores_0_externalInterrupt_plic_target_requests_14_valid = (userInterruptD_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_1);
  assign system_cores_0_externalInterrupt_plic_target_requests_15_priority = system_axiA_interrupt_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_15_id = 6'h1e;
  assign system_cores_0_externalInterrupt_plic_target_requests_15_valid = (system_axiA_interrupt_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_4);
  assign system_cores_0_externalInterrupt_plic_target_requests_16_priority = system_watchdog_logic_panics_0_plic_gateway_priority;
  assign system_cores_0_externalInterrupt_plic_target_requests_16_id = 6'h20;
  assign system_cores_0_externalInterrupt_plic_target_requests_16_valid = (system_watchdog_logic_panics_0_plic_gateway_ip && system_cores_0_externalInterrupt_plic_target_ie_15);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id = ((! system_cores_0_externalInterrupt_plic_target_requests_1_valid) || (system_cores_0_externalInterrupt_plic_target_requests_0_valid && (system_cores_0_externalInterrupt_plic_target_requests_1_priority <= system_cores_0_externalInterrupt_plic_target_requests_0_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_1 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id ? system_cores_0_externalInterrupt_plic_target_requests_0_priority : system_cores_0_externalInterrupt_plic_target_requests_1_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_2 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id ? system_cores_0_externalInterrupt_plic_target_requests_0_valid : system_cores_0_externalInterrupt_plic_target_requests_1_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_3 = ((! system_cores_0_externalInterrupt_plic_target_requests_3_valid) || (system_cores_0_externalInterrupt_plic_target_requests_2_valid && (system_cores_0_externalInterrupt_plic_target_requests_3_priority <= system_cores_0_externalInterrupt_plic_target_requests_2_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_4 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_3 ? system_cores_0_externalInterrupt_plic_target_requests_2_priority : system_cores_0_externalInterrupt_plic_target_requests_3_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_5 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_3 ? system_cores_0_externalInterrupt_plic_target_requests_2_valid : system_cores_0_externalInterrupt_plic_target_requests_3_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_6 = ((! system_cores_0_externalInterrupt_plic_target_requests_5_valid) || (system_cores_0_externalInterrupt_plic_target_requests_4_valid && (system_cores_0_externalInterrupt_plic_target_requests_5_priority <= system_cores_0_externalInterrupt_plic_target_requests_4_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_7 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_6 ? system_cores_0_externalInterrupt_plic_target_requests_4_priority : system_cores_0_externalInterrupt_plic_target_requests_5_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_8 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_6 ? system_cores_0_externalInterrupt_plic_target_requests_4_valid : system_cores_0_externalInterrupt_plic_target_requests_5_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_9 = ((! system_cores_0_externalInterrupt_plic_target_requests_7_valid) || (system_cores_0_externalInterrupt_plic_target_requests_6_valid && (system_cores_0_externalInterrupt_plic_target_requests_7_priority <= system_cores_0_externalInterrupt_plic_target_requests_6_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_10 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_9 ? system_cores_0_externalInterrupt_plic_target_requests_6_priority : system_cores_0_externalInterrupt_plic_target_requests_7_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_11 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_9 ? system_cores_0_externalInterrupt_plic_target_requests_6_valid : system_cores_0_externalInterrupt_plic_target_requests_7_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_12 = ((! system_cores_0_externalInterrupt_plic_target_requests_9_valid) || (system_cores_0_externalInterrupt_plic_target_requests_8_valid && (system_cores_0_externalInterrupt_plic_target_requests_9_priority <= system_cores_0_externalInterrupt_plic_target_requests_8_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_13 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_12 ? system_cores_0_externalInterrupt_plic_target_requests_8_priority : system_cores_0_externalInterrupt_plic_target_requests_9_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_14 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_12 ? system_cores_0_externalInterrupt_plic_target_requests_8_valid : system_cores_0_externalInterrupt_plic_target_requests_9_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_15 = ((! system_cores_0_externalInterrupt_plic_target_requests_11_valid) || (system_cores_0_externalInterrupt_plic_target_requests_10_valid && (system_cores_0_externalInterrupt_plic_target_requests_11_priority <= system_cores_0_externalInterrupt_plic_target_requests_10_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_16 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_15 ? system_cores_0_externalInterrupt_plic_target_requests_10_priority : system_cores_0_externalInterrupt_plic_target_requests_11_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_17 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_15 ? system_cores_0_externalInterrupt_plic_target_requests_10_valid : system_cores_0_externalInterrupt_plic_target_requests_11_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_18 = ((! system_cores_0_externalInterrupt_plic_target_requests_13_valid) || (system_cores_0_externalInterrupt_plic_target_requests_12_valid && (system_cores_0_externalInterrupt_plic_target_requests_13_priority <= system_cores_0_externalInterrupt_plic_target_requests_12_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_19 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_18 ? system_cores_0_externalInterrupt_plic_target_requests_12_priority : system_cores_0_externalInterrupt_plic_target_requests_13_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_20 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_18 ? system_cores_0_externalInterrupt_plic_target_requests_12_valid : system_cores_0_externalInterrupt_plic_target_requests_13_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_21 = ((! system_cores_0_externalInterrupt_plic_target_requests_15_valid) || (system_cores_0_externalInterrupt_plic_target_requests_14_valid && (system_cores_0_externalInterrupt_plic_target_requests_15_priority <= system_cores_0_externalInterrupt_plic_target_requests_14_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_22 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_21 ? system_cores_0_externalInterrupt_plic_target_requests_14_priority : system_cores_0_externalInterrupt_plic_target_requests_15_priority);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_23 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_21 ? system_cores_0_externalInterrupt_plic_target_requests_14_valid : system_cores_0_externalInterrupt_plic_target_requests_15_valid);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_24 = ((! _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_5) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_2 && (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_4 <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_1)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_25 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_24 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_1 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_4);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_26 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_24 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_2 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_5);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_27 = ((! _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_11) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_8 && (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_10 <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_7)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_28 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_27 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_7 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_10);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_29 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_27 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_8 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_11);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_30 = ((! _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_17) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_14 && (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_16 <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_13)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_31 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_30 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_13 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_16);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_32 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_30 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_14 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_17);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_33 = ((! _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_23) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_20 && (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_22 <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_19)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_34 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_33 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_19 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_22);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_35 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_33 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_20 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_23);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_36 = ((! _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_29) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_26 && (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_28 <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_25)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_36 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_25 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_28);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_37 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_36 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_26 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_29);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_38 = ((! _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_35) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_32 && (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_34 <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_31)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_1 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_38 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_31 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_34);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_39 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_38 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_32 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_35);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_40 = ((! _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_39) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_37 && (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_1 <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority)));
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_2 = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_40 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_1);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_valid = (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_40 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_37 : _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_39);
  assign _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_3 = ((! system_cores_0_externalInterrupt_plic_target_requests_16_valid) || (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_valid && (system_cores_0_externalInterrupt_plic_target_requests_16_priority <= _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_2)));
  assign system_cores_0_externalInterrupt_plic_target_iep = (system_cores_0_externalInterrupt_plic_target_threshold < system_cores_0_externalInterrupt_plic_target_bestRequest_priority);
  assign system_cores_0_externalInterrupt_plic_target_claim = (system_cores_0_externalInterrupt_plic_target_iep ? system_cores_0_externalInterrupt_plic_target_bestRequest_id : 6'h0);
  assign system_cores_1_externalInterrupt_plic_target_requests_0_priority = 2'b00;
  assign system_cores_1_externalInterrupt_plic_target_requests_0_id = 6'h0;
  assign system_cores_1_externalInterrupt_plic_target_requests_0_valid = 1'b1;
  assign system_cores_1_externalInterrupt_plic_target_requests_1_priority = system_uart_0_io_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_1_id = 6'h01;
  assign system_cores_1_externalInterrupt_plic_target_requests_1_valid = (system_uart_0_io_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_5);
  assign system_cores_1_externalInterrupt_plic_target_requests_2_priority = system_spi_0_io_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_2_id = 6'h04;
  assign system_cores_1_externalInterrupt_plic_target_requests_2_valid = (system_spi_0_io_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_6);
  assign system_cores_1_externalInterrupt_plic_target_requests_3_priority = system_spi_1_io_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_3_id = 6'h05;
  assign system_cores_1_externalInterrupt_plic_target_requests_3_valid = (system_spi_1_io_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_7);
  assign system_cores_1_externalInterrupt_plic_target_requests_4_priority = system_i2c_0_io_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_4_id = 6'h08;
  assign system_cores_1_externalInterrupt_plic_target_requests_4_valid = (system_i2c_0_io_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_8);
  assign system_cores_1_externalInterrupt_plic_target_requests_5_priority = system_i2c_1_io_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_5_id = 6'h09;
  assign system_cores_1_externalInterrupt_plic_target_requests_5_valid = (system_i2c_1_io_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_10);
  assign system_cores_1_externalInterrupt_plic_target_requests_6_priority = system_i2c_2_io_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_6_id = 6'h0a;
  assign system_cores_1_externalInterrupt_plic_target_requests_6_valid = (system_i2c_2_io_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_9);
  assign system_cores_1_externalInterrupt_plic_target_requests_7_priority = system_gpio_0_io_interrupts_0_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_7_id = 6'h0c;
  assign system_cores_1_externalInterrupt_plic_target_requests_7_valid = (system_gpio_0_io_interrupts_0_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_13);
  assign system_cores_1_externalInterrupt_plic_target_requests_8_priority = system_gpio_0_io_interrupts_1_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_8_id = 6'h0d;
  assign system_cores_1_externalInterrupt_plic_target_requests_8_valid = (system_gpio_0_io_interrupts_1_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_14);
  assign system_cores_1_externalInterrupt_plic_target_requests_9_priority = userInterruptA_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_9_id = 6'h10;
  assign system_cores_1_externalInterrupt_plic_target_requests_9_valid = (userInterruptA_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_0);
  assign system_cores_1_externalInterrupt_plic_target_requests_10_priority = userInterruptB_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_10_id = 6'h11;
  assign system_cores_1_externalInterrupt_plic_target_requests_10_valid = (userInterruptB_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_3);
  assign system_cores_1_externalInterrupt_plic_target_requests_11_priority = system_userTimer_0_interrupts_0_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_11_id = 6'h13;
  assign system_cores_1_externalInterrupt_plic_target_requests_11_valid = (system_userTimer_0_interrupts_0_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_12);
  assign system_cores_1_externalInterrupt_plic_target_requests_12_priority = system_userTimer_1_interrupts_0_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_12_id = 6'h14;
  assign system_cores_1_externalInterrupt_plic_target_requests_12_valid = (system_userTimer_1_interrupts_0_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_11);
  assign system_cores_1_externalInterrupt_plic_target_requests_13_priority = userInterruptC_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_13_id = 6'h16;
  assign system_cores_1_externalInterrupt_plic_target_requests_13_valid = (userInterruptC_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_2);
  assign system_cores_1_externalInterrupt_plic_target_requests_14_priority = userInterruptD_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_14_id = 6'h17;
  assign system_cores_1_externalInterrupt_plic_target_requests_14_valid = (userInterruptD_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_1);
  assign system_cores_1_externalInterrupt_plic_target_requests_15_priority = system_axiA_interrupt_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_15_id = 6'h1e;
  assign system_cores_1_externalInterrupt_plic_target_requests_15_valid = (system_axiA_interrupt_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_4);
  assign system_cores_1_externalInterrupt_plic_target_requests_16_priority = system_watchdog_logic_panics_0_plic_gateway_priority;
  assign system_cores_1_externalInterrupt_plic_target_requests_16_id = 6'h20;
  assign system_cores_1_externalInterrupt_plic_target_requests_16_valid = (system_watchdog_logic_panics_0_plic_gateway_ip && system_cores_1_externalInterrupt_plic_target_ie_15);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id = ((! system_cores_1_externalInterrupt_plic_target_requests_1_valid) || (system_cores_1_externalInterrupt_plic_target_requests_0_valid && (system_cores_1_externalInterrupt_plic_target_requests_1_priority <= system_cores_1_externalInterrupt_plic_target_requests_0_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_1 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id ? system_cores_1_externalInterrupt_plic_target_requests_0_priority : system_cores_1_externalInterrupt_plic_target_requests_1_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_2 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id ? system_cores_1_externalInterrupt_plic_target_requests_0_valid : system_cores_1_externalInterrupt_plic_target_requests_1_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_3 = ((! system_cores_1_externalInterrupt_plic_target_requests_3_valid) || (system_cores_1_externalInterrupt_plic_target_requests_2_valid && (system_cores_1_externalInterrupt_plic_target_requests_3_priority <= system_cores_1_externalInterrupt_plic_target_requests_2_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_4 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_3 ? system_cores_1_externalInterrupt_plic_target_requests_2_priority : system_cores_1_externalInterrupt_plic_target_requests_3_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_5 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_3 ? system_cores_1_externalInterrupt_plic_target_requests_2_valid : system_cores_1_externalInterrupt_plic_target_requests_3_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_6 = ((! system_cores_1_externalInterrupt_plic_target_requests_5_valid) || (system_cores_1_externalInterrupt_plic_target_requests_4_valid && (system_cores_1_externalInterrupt_plic_target_requests_5_priority <= system_cores_1_externalInterrupt_plic_target_requests_4_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_7 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_6 ? system_cores_1_externalInterrupt_plic_target_requests_4_priority : system_cores_1_externalInterrupt_plic_target_requests_5_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_8 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_6 ? system_cores_1_externalInterrupt_plic_target_requests_4_valid : system_cores_1_externalInterrupt_plic_target_requests_5_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_9 = ((! system_cores_1_externalInterrupt_plic_target_requests_7_valid) || (system_cores_1_externalInterrupt_plic_target_requests_6_valid && (system_cores_1_externalInterrupt_plic_target_requests_7_priority <= system_cores_1_externalInterrupt_plic_target_requests_6_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_10 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_9 ? system_cores_1_externalInterrupt_plic_target_requests_6_priority : system_cores_1_externalInterrupt_plic_target_requests_7_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_11 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_9 ? system_cores_1_externalInterrupt_plic_target_requests_6_valid : system_cores_1_externalInterrupt_plic_target_requests_7_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_12 = ((! system_cores_1_externalInterrupt_plic_target_requests_9_valid) || (system_cores_1_externalInterrupt_plic_target_requests_8_valid && (system_cores_1_externalInterrupt_plic_target_requests_9_priority <= system_cores_1_externalInterrupt_plic_target_requests_8_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_13 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_12 ? system_cores_1_externalInterrupt_plic_target_requests_8_priority : system_cores_1_externalInterrupt_plic_target_requests_9_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_14 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_12 ? system_cores_1_externalInterrupt_plic_target_requests_8_valid : system_cores_1_externalInterrupt_plic_target_requests_9_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_15 = ((! system_cores_1_externalInterrupt_plic_target_requests_11_valid) || (system_cores_1_externalInterrupt_plic_target_requests_10_valid && (system_cores_1_externalInterrupt_plic_target_requests_11_priority <= system_cores_1_externalInterrupt_plic_target_requests_10_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_16 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_15 ? system_cores_1_externalInterrupt_plic_target_requests_10_priority : system_cores_1_externalInterrupt_plic_target_requests_11_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_17 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_15 ? system_cores_1_externalInterrupt_plic_target_requests_10_valid : system_cores_1_externalInterrupt_plic_target_requests_11_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_18 = ((! system_cores_1_externalInterrupt_plic_target_requests_13_valid) || (system_cores_1_externalInterrupt_plic_target_requests_12_valid && (system_cores_1_externalInterrupt_plic_target_requests_13_priority <= system_cores_1_externalInterrupt_plic_target_requests_12_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_19 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_18 ? system_cores_1_externalInterrupt_plic_target_requests_12_priority : system_cores_1_externalInterrupt_plic_target_requests_13_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_20 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_18 ? system_cores_1_externalInterrupt_plic_target_requests_12_valid : system_cores_1_externalInterrupt_plic_target_requests_13_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_21 = ((! system_cores_1_externalInterrupt_plic_target_requests_15_valid) || (system_cores_1_externalInterrupt_plic_target_requests_14_valid && (system_cores_1_externalInterrupt_plic_target_requests_15_priority <= system_cores_1_externalInterrupt_plic_target_requests_14_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_22 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_21 ? system_cores_1_externalInterrupt_plic_target_requests_14_priority : system_cores_1_externalInterrupt_plic_target_requests_15_priority);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_23 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_21 ? system_cores_1_externalInterrupt_plic_target_requests_14_valid : system_cores_1_externalInterrupt_plic_target_requests_15_valid);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_24 = ((! _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_5) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_2 && (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_4 <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_1)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_25 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_24 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_1 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_4);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_26 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_24 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_2 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_5);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_27 = ((! _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_11) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_8 && (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_10 <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_7)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_28 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_27 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_7 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_10);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_29 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_27 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_8 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_11);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_30 = ((! _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_17) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_14 && (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_16 <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_13)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_31 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_30 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_13 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_16);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_32 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_30 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_14 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_17);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_33 = ((! _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_23) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_20 && (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_22 <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_19)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_34 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_33 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_19 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_22);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_35 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_33 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_20 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_23);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_36 = ((! _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_29) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_26 && (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_28 <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_25)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_36 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_25 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_28);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_37 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_36 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_26 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_29);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_38 = ((! _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_35) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_32 && (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_34 <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_31)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_1 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_38 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_31 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_34);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_39 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_38 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_32 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_35);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_40 = ((! _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_39) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_37 && (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_1 <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority)));
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_2 = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_40 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_1);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_valid = (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_40 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_37 : _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_39);
  assign _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_3 = ((! system_cores_1_externalInterrupt_plic_target_requests_16_valid) || (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_valid && (system_cores_1_externalInterrupt_plic_target_requests_16_priority <= _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_2)));
  assign system_cores_1_externalInterrupt_plic_target_iep = (system_cores_1_externalInterrupt_plic_target_threshold < system_cores_1_externalInterrupt_plic_target_bestRequest_priority);
  assign system_cores_1_externalInterrupt_plic_target_claim = (system_cores_1_externalInterrupt_plic_target_iep ? system_cores_1_externalInterrupt_plic_target_bestRequest_id : 6'h0);
  assign userInterruptA_interrupt_plic_gateway_priority = _zz_userInterruptA_interrupt_plic_gateway_priority;
  assign userInterruptD_interrupt_plic_gateway_priority = _zz_userInterruptD_interrupt_plic_gateway_priority;
  assign userInterruptC_interrupt_plic_gateway_priority = _zz_userInterruptC_interrupt_plic_gateway_priority;
  assign userInterruptB_interrupt_plic_gateway_priority = _zz_userInterruptB_interrupt_plic_gateway_priority;
  assign system_axiA_interrupt_plic_gateway_priority = _zz_system_axiA_interrupt_plic_gateway_priority;
  assign system_uart_0_io_interrupt_plic_gateway_priority = _zz_system_uart_0_io_interrupt_plic_gateway_priority;
  assign system_spi_0_io_interrupt_plic_gateway_priority = _zz_system_spi_0_io_interrupt_plic_gateway_priority;
  assign system_spi_1_io_interrupt_plic_gateway_priority = _zz_system_spi_1_io_interrupt_plic_gateway_priority;
  assign system_i2c_0_io_interrupt_plic_gateway_priority = _zz_system_i2c_0_io_interrupt_plic_gateway_priority;
  assign system_i2c_2_io_interrupt_plic_gateway_priority = _zz_system_i2c_2_io_interrupt_plic_gateway_priority;
  assign system_i2c_1_io_interrupt_plic_gateway_priority = _zz_system_i2c_1_io_interrupt_plic_gateway_priority;
  assign system_userTimer_1_interrupts_0_plic_gateway_priority = _zz_system_userTimer_1_interrupts_0_plic_gateway_priority;
  assign system_userTimer_0_interrupts_0_plic_gateway_priority = _zz_system_userTimer_0_interrupts_0_plic_gateway_priority;
  assign system_gpio_0_io_interrupts_0_plic_gateway_priority = _zz_system_gpio_0_io_interrupts_0_plic_gateway_priority;
  assign system_gpio_0_io_interrupts_1_plic_gateway_priority = _zz_system_gpio_0_io_interrupts_1_plic_gateway_priority;
  assign system_watchdog_logic_panics_0_plic_gateway_priority = _zz_system_watchdog_logic_panics_0_plic_gateway_priority;
  always @(*) begin
    system_plic_logic_bridge_claim_valid = 1'b0;
    case(system_plic_logic_bmb_cmd_payload_fragment_address)
      22'h200004 : begin
        if(system_plic_logic_bus_doRead) begin
          system_plic_logic_bridge_claim_valid = 1'b1;
        end
      end
      22'h201004 : begin
        if(system_plic_logic_bus_doRead) begin
          system_plic_logic_bridge_claim_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    system_plic_logic_bridge_claim_payload = 6'bxxxxxx;
    case(system_plic_logic_bmb_cmd_payload_fragment_address)
      22'h200004 : begin
        if(system_plic_logic_bus_doRead) begin
          system_plic_logic_bridge_claim_payload = system_cores_0_externalInterrupt_plic_target_claim;
        end
      end
      22'h201004 : begin
        if(system_plic_logic_bus_doRead) begin
          system_plic_logic_bridge_claim_payload = system_cores_1_externalInterrupt_plic_target_claim;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    system_plic_logic_bridge_completion_valid = 1'b0;
    if(system_plic_logic_bridge_targetMapping_0_targetCompletion_valid) begin
      system_plic_logic_bridge_completion_valid = 1'b1;
    end
    if(system_plic_logic_bridge_targetMapping_1_targetCompletion_valid) begin
      system_plic_logic_bridge_completion_valid = 1'b1;
    end
  end

  always @(*) begin
    system_plic_logic_bridge_completion_payload = 6'bxxxxxx;
    if(system_plic_logic_bridge_targetMapping_0_targetCompletion_valid) begin
      system_plic_logic_bridge_completion_payload = system_plic_logic_bridge_targetMapping_0_targetCompletion_payload;
    end
    if(system_plic_logic_bridge_targetMapping_1_targetCompletion_valid) begin
      system_plic_logic_bridge_completion_payload = system_plic_logic_bridge_targetMapping_1_targetCompletion_payload;
    end
  end

  always @(*) begin
    system_plic_logic_bridge_coherencyStall_willIncrement = 1'b0;
    if(when_PlicMapper_l122) begin
      system_plic_logic_bridge_coherencyStall_willIncrement = 1'b1;
    end
    if(when_BmbSlaveFactory_l77) begin
      if(system_plic_logic_bus_askWrite) begin
        system_plic_logic_bridge_coherencyStall_willIncrement = 1'b1;
      end
      if(system_plic_logic_bus_askRead) begin
        system_plic_logic_bridge_coherencyStall_willIncrement = 1'b1;
      end
    end
  end

  assign system_plic_logic_bridge_coherencyStall_willClear = 1'b0;
  assign system_plic_logic_bridge_coherencyStall_willOverflowIfInc = (system_plic_logic_bridge_coherencyStall_value == 1'b1);
  assign system_plic_logic_bridge_coherencyStall_willOverflow = (system_plic_logic_bridge_coherencyStall_willOverflowIfInc && system_plic_logic_bridge_coherencyStall_willIncrement);
  always @(*) begin
    system_plic_logic_bridge_coherencyStall_valueNext = (system_plic_logic_bridge_coherencyStall_value + system_plic_logic_bridge_coherencyStall_willIncrement);
    if(system_plic_logic_bridge_coherencyStall_willClear) begin
      system_plic_logic_bridge_coherencyStall_valueNext = 1'b0;
    end
  end

  assign when_PlicMapper_l122 = (system_plic_logic_bridge_coherencyStall_value != 1'b0);
  assign system_cores_0_externalInterrupt_plic_target_threshold = _zz_system_cores_0_externalInterrupt_plic_target_threshold;
  always @(*) begin
    system_plic_logic_bridge_targetMapping_0_targetCompletion_valid = 1'b0;
    case(system_plic_logic_bmb_cmd_payload_fragment_address)
      22'h200004 : begin
        if(system_plic_logic_bus_doWrite) begin
          system_plic_logic_bridge_targetMapping_0_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign system_cores_0_externalInterrupt_plic_target_ie_0 = _zz_system_cores_0_externalInterrupt_plic_target_ie_0;
  assign system_cores_0_externalInterrupt_plic_target_ie_1 = _zz_system_cores_0_externalInterrupt_plic_target_ie_1;
  assign system_cores_0_externalInterrupt_plic_target_ie_2 = _zz_system_cores_0_externalInterrupt_plic_target_ie_2;
  assign system_cores_0_externalInterrupt_plic_target_ie_3 = _zz_system_cores_0_externalInterrupt_plic_target_ie_3;
  assign system_cores_0_externalInterrupt_plic_target_ie_4 = _zz_system_cores_0_externalInterrupt_plic_target_ie_4;
  assign system_cores_0_externalInterrupt_plic_target_ie_5 = _zz_system_cores_0_externalInterrupt_plic_target_ie_5;
  assign system_cores_0_externalInterrupt_plic_target_ie_6 = _zz_system_cores_0_externalInterrupt_plic_target_ie_6;
  assign system_cores_0_externalInterrupt_plic_target_ie_7 = _zz_system_cores_0_externalInterrupt_plic_target_ie_7;
  assign system_cores_0_externalInterrupt_plic_target_ie_8 = _zz_system_cores_0_externalInterrupt_plic_target_ie_8;
  assign system_cores_0_externalInterrupt_plic_target_ie_9 = _zz_system_cores_0_externalInterrupt_plic_target_ie_9;
  assign system_cores_0_externalInterrupt_plic_target_ie_10 = _zz_system_cores_0_externalInterrupt_plic_target_ie_10;
  assign system_cores_0_externalInterrupt_plic_target_ie_11 = _zz_system_cores_0_externalInterrupt_plic_target_ie_11;
  assign system_cores_0_externalInterrupt_plic_target_ie_12 = _zz_system_cores_0_externalInterrupt_plic_target_ie_12;
  assign system_cores_0_externalInterrupt_plic_target_ie_13 = _zz_system_cores_0_externalInterrupt_plic_target_ie_13;
  assign system_cores_0_externalInterrupt_plic_target_ie_14 = _zz_system_cores_0_externalInterrupt_plic_target_ie_14;
  assign system_cores_0_externalInterrupt_plic_target_ie_15 = _zz_system_cores_0_externalInterrupt_plic_target_ie_15;
  assign system_cores_1_externalInterrupt_plic_target_threshold = _zz_system_cores_1_externalInterrupt_plic_target_threshold;
  always @(*) begin
    system_plic_logic_bridge_targetMapping_1_targetCompletion_valid = 1'b0;
    case(system_plic_logic_bmb_cmd_payload_fragment_address)
      22'h201004 : begin
        if(system_plic_logic_bus_doWrite) begin
          system_plic_logic_bridge_targetMapping_1_targetCompletion_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign system_cores_1_externalInterrupt_plic_target_ie_0 = _zz_system_cores_1_externalInterrupt_plic_target_ie_0;
  assign system_cores_1_externalInterrupt_plic_target_ie_1 = _zz_system_cores_1_externalInterrupt_plic_target_ie_1;
  assign system_cores_1_externalInterrupt_plic_target_ie_2 = _zz_system_cores_1_externalInterrupt_plic_target_ie_2;
  assign system_cores_1_externalInterrupt_plic_target_ie_3 = _zz_system_cores_1_externalInterrupt_plic_target_ie_3;
  assign system_cores_1_externalInterrupt_plic_target_ie_4 = _zz_system_cores_1_externalInterrupt_plic_target_ie_4;
  assign system_cores_1_externalInterrupt_plic_target_ie_5 = _zz_system_cores_1_externalInterrupt_plic_target_ie_5;
  assign system_cores_1_externalInterrupt_plic_target_ie_6 = _zz_system_cores_1_externalInterrupt_plic_target_ie_6;
  assign system_cores_1_externalInterrupt_plic_target_ie_7 = _zz_system_cores_1_externalInterrupt_plic_target_ie_7;
  assign system_cores_1_externalInterrupt_plic_target_ie_8 = _zz_system_cores_1_externalInterrupt_plic_target_ie_8;
  assign system_cores_1_externalInterrupt_plic_target_ie_9 = _zz_system_cores_1_externalInterrupt_plic_target_ie_9;
  assign system_cores_1_externalInterrupt_plic_target_ie_10 = _zz_system_cores_1_externalInterrupt_plic_target_ie_10;
  assign system_cores_1_externalInterrupt_plic_target_ie_11 = _zz_system_cores_1_externalInterrupt_plic_target_ie_11;
  assign system_cores_1_externalInterrupt_plic_target_ie_12 = _zz_system_cores_1_externalInterrupt_plic_target_ie_12;
  assign system_cores_1_externalInterrupt_plic_target_ie_13 = _zz_system_cores_1_externalInterrupt_plic_target_ie_13;
  assign system_cores_1_externalInterrupt_plic_target_ie_14 = _zz_system_cores_1_externalInterrupt_plic_target_ie_14;
  assign system_cores_1_externalInterrupt_plic_target_ie_15 = _zz_system_cores_1_externalInterrupt_plic_target_ie_15;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_11 = system_bmbPeripheral_bmb_decoder_io_outputs_12_cmd_payload_fragment_context;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_11;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_11 = io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_11 = io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_11;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_11;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_11 = io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_11;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_11[15:0];
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_11;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_11;
  assign io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_11;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_11 = io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_11 = io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_11 = io_apbSlave_2_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_12 = system_bmbPeripheral_bmb_decoder_io_outputs_13_cmd_payload_fragment_context;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_12;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_12 = io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_12 = io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_12;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_12;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_12 = io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_12;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_12[15:0];
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_12;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_12;
  assign io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_12;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_12 = io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_12 = io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_12 = io_apbSlave_1_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_13 = system_bmbPeripheral_bmb_decoder_io_outputs_14_cmd_payload_fragment_context;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_13;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_13 = io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_13 = io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_13;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_13;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_13 = io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_13;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_13[15:0];
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_13;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_13;
  assign io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_13;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_13 = io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_13 = io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_13 = io_apbSlave_4_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_14 = system_bmbPeripheral_bmb_decoder_io_outputs_15_cmd_payload_fragment_context;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_14;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_14 = io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_14 = io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_14;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_14;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_14 = io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_14;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_14[15:0];
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_14;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_14;
  assign io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_14;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_14 = io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_14 = io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_14 = io_apbSlave_0_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_15 = system_bmbPeripheral_bmb_decoder_io_outputs_16_cmd_payload_fragment_context;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_15;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_15 = io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_15 = io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_15;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_15;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_15 = io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_15;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_15[15:0];
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_15;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_15;
  assign io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_15;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_15 = io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_15 = io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_15 = io_apbSlave_3_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign jtagCtrl_tdo = system_riscvJtag_hard_noTap_tunnel_io_instruction_tdo;
  assign system_plic_logic_bmb_cmd_valid = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready = system_plic_logic_bmb_cmd_ready;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid = system_plic_logic_bmb_rsp_valid;
  assign system_plic_logic_bmb_rsp_ready = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready;
  assign system_plic_logic_bmb_cmd_payload_last = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last = system_plic_logic_bmb_rsp_payload_last;
  assign system_plic_logic_bmb_cmd_payload_fragment_opcode = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
  assign system_plic_logic_bmb_cmd_payload_fragment_address = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
  assign system_plic_logic_bmb_cmd_payload_fragment_length = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
  assign system_plic_logic_bmb_cmd_payload_fragment_data = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
  assign system_plic_logic_bmb_cmd_payload_fragment_context = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode = system_plic_logic_bmb_rsp_payload_fragment_opcode;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data = system_plic_logic_bmb_rsp_payload_fragment_data;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context = system_plic_logic_bmb_rsp_payload_fragment_context;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_valid_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_valid;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_ready_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_rsp_ready;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_last;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_address;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_length;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_16 = system_bmbPeripheral_bmb_decoder_io_outputs_0_cmd_payload_fragment_context;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid = system_bmbPeripheral_bmb_withoutMask_cmd_valid_16;
  assign system_bmbPeripheral_bmb_withoutMask_cmd_ready_16 = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_valid_16 = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready = system_bmbPeripheral_bmb_withoutMask_rsp_ready_16;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last = system_bmbPeripheral_bmb_withoutMask_cmd_payload_last_16;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_last_16 = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_opcode_16;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_address_16[21:0];
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_length_16;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_data_16;
  assign system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context = system_bmbPeripheral_bmb_withoutMask_cmd_payload_fragment_context_16;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_opcode_16 = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_data_16 = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
  assign system_bmbPeripheral_bmb_withoutMask_rsp_payload_fragment_context_16 = system_plic_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
  assign system_plic_logic_bridge_targetMapping_0_targetCompletion_payload = system_plic_logic_bmb_cmd_payload_fragment_data[5 : 0];
  assign system_plic_logic_bridge_targetMapping_1_targetCompletion_payload = system_plic_logic_bmb_cmd_payload_fragment_data[5 : 0];
  assign when_BmbSlaveFactory_l77 = 1'b1;
  always @(posedge io_systemClk) begin
    if(when_ClockDomainGenerator_l222) begin
      debugCd_logic_holdingLogic_resetCounter <= (debugCd_logic_holdingLogic_resetCounter + 12'h001);
    end
    if(debugCd_logic_inputResetTrigger) begin
      debugCd_logic_holdingLogic_resetCounter <= 12'h0;
    end
    debugCd_logic_outputReset <= debugCd_logic_outputResetUnbuffered;
  end

  always @(posedge io_memoryClk) begin
    if(when_ClockDomainGenerator_l222_1) begin
      ddrCd_logic_holdingLogic_resetCounter <= (ddrCd_logic_holdingLogic_resetCounter + 6'h01);
    end
    if(ddrCd_logic_inputResetTrigger) begin
      ddrCd_logic_holdingLogic_resetCounter <= 6'h0;
    end
    ddrCd_logic_outputReset <= ddrCd_logic_outputResetUnbuffered;
  end

  always @(posedge io_peripheralClk) begin
    if(when_ClockDomainGenerator_l222_2) begin
      peripheralCd_logic_holdingLogic_resetCounter <= (peripheralCd_logic_holdingLogic_resetCounter + 6'h01);
    end
    if(peripheralCd_logic_inputResetTrigger) begin
      peripheralCd_logic_holdingLogic_resetCounter <= 6'h0;
    end
    peripheralCd_logic_outputReset <= peripheralCd_logic_outputResetUnbuffered;
  end

  always @(posedge io_systemClk) begin
    if(when_ClockDomainGenerator_l222_3) begin
      systemCd_logic_holdingLogic_resetCounter <= (systemCd_logic_holdingLogic_resetCounter + 6'h01);
    end
    if(systemCd_logic_inputResetTrigger) begin
      systemCd_logic_holdingLogic_resetCounter <= 6'h0;
    end
    systemCd_logic_outputReset <= systemCd_logic_outputResetUnbuffered;
  end

  always @(posedge io_memoryClk) begin
    io_memoryReset <= ddrCd_logic_outputReset;
    if(system_ddr_ddrLogic_cc_fifo_io_output_cmd_ready) begin
      io_output_cmd_rData_last_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_last;
      io_output_cmd_rData_fragment_source_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_source;
      io_output_cmd_rData_fragment_opcode_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_opcode;
      io_output_cmd_rData_fragment_address_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_address;
      io_output_cmd_rData_fragment_length_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_length;
      io_output_cmd_rData_fragment_data_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_data;
      io_output_cmd_rData_fragment_mask_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_mask;
      io_output_cmd_rData_fragment_context_1 <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_payload_fragment_context;
    end
    if(_zz_io_input_rsp_ready_1) begin
      _zz_io_output_rsp_payload_last_1 <= system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_last;
      _zz_io_output_rsp_payload_fragment_source_1 <= system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_source;
      _zz_io_output_rsp_payload_fragment_opcode_1 <= system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_opcode;
      _zz_io_output_rsp_payload_fragment_data_1 <= system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_data;
      _zz_io_output_rsp_payload_fragment_context_1 <= system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_payload_fragment_context;
    end
    if(io_output_arw_rValidN) begin
      io_output_arw_rData_addr <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_addr;
      io_output_arw_rData_len <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_len;
      io_output_arw_rData_size <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_size;
      io_output_arw_rData_cache <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_cache;
      io_output_arw_rData_prot <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_prot;
      io_output_arw_rData_write <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_payload_write;
    end
    if(io_output_arw_s2mPipe_ready) begin
      io_output_arw_s2mPipe_rData_addr <= io_output_arw_s2mPipe_payload_addr;
      io_output_arw_s2mPipe_rData_len <= io_output_arw_s2mPipe_payload_len;
      io_output_arw_s2mPipe_rData_size <= io_output_arw_s2mPipe_payload_size;
      io_output_arw_s2mPipe_rData_cache <= io_output_arw_s2mPipe_payload_cache;
      io_output_arw_s2mPipe_rData_prot <= io_output_arw_s2mPipe_payload_prot;
      io_output_arw_s2mPipe_rData_write <= io_output_arw_s2mPipe_payload_write;
    end
    if(io_output_arw_s2mPipe_m2sPipe_ready) begin
      io_output_arw_s2mPipe_m2sPipe_rData_addr <= io_output_arw_s2mPipe_m2sPipe_payload_addr;
      io_output_arw_s2mPipe_m2sPipe_rData_len <= io_output_arw_s2mPipe_m2sPipe_payload_len;
      io_output_arw_s2mPipe_m2sPipe_rData_size <= io_output_arw_s2mPipe_m2sPipe_payload_size;
      io_output_arw_s2mPipe_m2sPipe_rData_cache <= io_output_arw_s2mPipe_m2sPipe_payload_cache;
      io_output_arw_s2mPipe_m2sPipe_rData_prot <= io_output_arw_s2mPipe_m2sPipe_payload_prot;
      io_output_arw_s2mPipe_m2sPipe_rData_write <= io_output_arw_s2mPipe_m2sPipe_payload_write;
    end
    if(io_output_w_rValidN) begin
      io_output_w_rData_data <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_data;
      io_output_w_rData_strb <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_strb;
      io_output_w_rData_last <= system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_payload_last;
    end
    if(io_output_w_s2mPipe_ready) begin
      io_output_w_s2mPipe_rData_data <= io_output_w_s2mPipe_payload_data;
      io_output_w_s2mPipe_rData_strb <= io_output_w_s2mPipe_payload_strb;
      io_output_w_s2mPipe_rData_last <= io_output_w_s2mPipe_payload_last;
    end
    if(io_output_w_s2mPipe_m2sPipe_ready) begin
      io_output_w_s2mPipe_m2sPipe_rData_data <= io_output_w_s2mPipe_m2sPipe_payload_data;
      io_output_w_s2mPipe_m2sPipe_rData_strb <= io_output_w_s2mPipe_m2sPipe_payload_strb;
      io_output_w_s2mPipe_m2sPipe_rData_last <= io_output_w_s2mPipe_m2sPipe_payload_last;
    end
    if(system_ddr_ddrLogic_cpuAccess_b_ready) begin
      system_ddr_ddrLogic_cpuAccess_b_rData_resp <= system_ddr_ddrLogic_cpuAccess_b_payload_resp;
    end
    if(system_ddr_ddrLogic_cpuAccess_b_s2mPipe_ready) begin
      system_ddr_ddrLogic_cpuAccess_b_s2mPipe_rData_resp <= system_ddr_ddrLogic_cpuAccess_b_s2mPipe_payload_resp;
    end
    if(system_ddr_ddrLogic_cpuAccess_r_ready) begin
      system_ddr_ddrLogic_cpuAccess_r_rData_data <= system_ddr_ddrLogic_cpuAccess_r_payload_data;
      system_ddr_ddrLogic_cpuAccess_r_rData_resp <= system_ddr_ddrLogic_cpuAccess_r_payload_resp;
      system_ddr_ddrLogic_cpuAccess_r_rData_last <= system_ddr_ddrLogic_cpuAccess_r_payload_last;
    end
    if(system_ddr_ddrLogic_cpuAccess_r_s2mPipe_ready) begin
      system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_data <= system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_data;
      system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_resp <= system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_resp;
      system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rData_last <= system_ddr_ddrLogic_cpuAccess_r_s2mPipe_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_ready) begin
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_addr <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_addr;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_id <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_id;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_region <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_region;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_len <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_len;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_size <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_size;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_burst <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_burst;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_lock <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_lock;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_cache <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_cache;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_qos <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_qos;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rData_prot <= system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_payload_prot;
    end
    if(system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_ready) begin
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_addr <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_addr;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_id <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_id;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_region <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_region;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_len <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_len;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_size <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_size;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_burst <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_burst;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_lock <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_lock;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_cache <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_cache;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_qos <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_qos;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rData_prot <= system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_payload_prot;
    end
    if(system_ddr_ddrLogic_userAdapters_0_userAxi4_w_ready) begin
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_data <= system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_data;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_strb <= system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_strb;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rData_last <= system_ddr_ddrLogic_userAdapters_0_userAxi4_w_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_ready) begin
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_data <= system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_data;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_strb <= system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_strb;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rData_last <= system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_ready) begin
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_data <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_data;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_id <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_id;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_resp <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_resp;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rData_last <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_ready) begin
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_data <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_data;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_id <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_id;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_resp <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_resp;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rData_last <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_ready) begin
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rData_id <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_payload_id;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rData_resp <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_payload_resp;
    end
    if(system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_ready) begin
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_addr <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_addr;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_id <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_id;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_region <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_region;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_len <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_len;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_size <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_size;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_burst <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_burst;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_lock <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_lock;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_cache <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_cache;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_qos <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_qos;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rData_prot <= system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_payload_prot;
    end
    if(system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_ready) begin
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_addr <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_addr;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_id <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_id;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_region <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_region;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_len <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_len;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_size <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_size;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_burst <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_burst;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_lock <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_lock;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_cache <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_cache;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_qos <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_qos;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rData_prot <= system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_payload_prot;
    end
    if(system_ddr_ddrLogic_userAdapters_1_userAxi4_w_ready) begin
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_data <= system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_data;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_strb <= system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_strb;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rData_last <= system_ddr_ddrLogic_userAdapters_1_userAxi4_w_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_ready) begin
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_data <= system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_data;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_strb <= system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_strb;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rData_last <= system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_ready) begin
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_data <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_data;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_id <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_id;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_resp <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_resp;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rData_last <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_ready) begin
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_data <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_data;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_id <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_id;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_resp <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_resp;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rData_last <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_ready) begin
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rData_id <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_payload_id;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rData_resp <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_payload_resp;
    end
    if(io_output_aw_rValidN) begin
      io_output_aw_rData_addr <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_addr;
      io_output_aw_rData_id <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_id;
      io_output_aw_rData_region <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_region;
      io_output_aw_rData_len <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_len;
      io_output_aw_rData_size <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_size;
      io_output_aw_rData_burst <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_burst;
      io_output_aw_rData_lock <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_lock;
      io_output_aw_rData_cache <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_cache;
      io_output_aw_rData_qos <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_qos;
      io_output_aw_rData_prot <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_payload_prot;
    end
    if(io_output_aw_s2mPipe_ready) begin
      io_output_aw_s2mPipe_rData_addr <= io_output_aw_s2mPipe_payload_addr;
      io_output_aw_s2mPipe_rData_id <= io_output_aw_s2mPipe_payload_id;
      io_output_aw_s2mPipe_rData_region <= io_output_aw_s2mPipe_payload_region;
      io_output_aw_s2mPipe_rData_len <= io_output_aw_s2mPipe_payload_len;
      io_output_aw_s2mPipe_rData_size <= io_output_aw_s2mPipe_payload_size;
      io_output_aw_s2mPipe_rData_burst <= io_output_aw_s2mPipe_payload_burst;
      io_output_aw_s2mPipe_rData_lock <= io_output_aw_s2mPipe_payload_lock;
      io_output_aw_s2mPipe_rData_cache <= io_output_aw_s2mPipe_payload_cache;
      io_output_aw_s2mPipe_rData_qos <= io_output_aw_s2mPipe_payload_qos;
      io_output_aw_s2mPipe_rData_prot <= io_output_aw_s2mPipe_payload_prot;
    end
    if(io_output_ar_rValidN) begin
      io_output_ar_rData_addr <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_addr;
      io_output_ar_rData_id <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_id;
      io_output_ar_rData_region <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_region;
      io_output_ar_rData_len <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_len;
      io_output_ar_rData_size <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_size;
      io_output_ar_rData_burst <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_burst;
      io_output_ar_rData_lock <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_lock;
      io_output_ar_rData_cache <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_cache;
      io_output_ar_rData_qos <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_qos;
      io_output_ar_rData_prot <= system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_payload_prot;
    end
    if(io_output_ar_s2mPipe_ready) begin
      io_output_ar_s2mPipe_rData_addr <= io_output_ar_s2mPipe_payload_addr;
      io_output_ar_s2mPipe_rData_id <= io_output_ar_s2mPipe_payload_id;
      io_output_ar_s2mPipe_rData_region <= io_output_ar_s2mPipe_payload_region;
      io_output_ar_s2mPipe_rData_len <= io_output_ar_s2mPipe_payload_len;
      io_output_ar_s2mPipe_rData_size <= io_output_ar_s2mPipe_payload_size;
      io_output_ar_s2mPipe_rData_burst <= io_output_ar_s2mPipe_payload_burst;
      io_output_ar_s2mPipe_rData_lock <= io_output_ar_s2mPipe_payload_lock;
      io_output_ar_s2mPipe_rData_cache <= io_output_ar_s2mPipe_payload_cache;
      io_output_ar_s2mPipe_rData_qos <= io_output_ar_s2mPipe_payload_qos;
      io_output_ar_s2mPipe_rData_prot <= io_output_ar_s2mPipe_payload_prot;
    end
    if(system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_ready) begin
      io_output_w_rData_data_1 <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_data;
      io_output_w_rData_strb_1 <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_strb;
      io_output_w_rData_last_1 <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_payload_last;
    end
    if(system_ddr_ddrLogic_ddrAAxi4_b_ready) begin
      system_ddr_ddrLogic_ddrAAxi4_b_rData_id <= system_ddr_ddrLogic_ddrAAxi4_b_payload_id;
      system_ddr_ddrLogic_ddrAAxi4_b_rData_resp <= system_ddr_ddrLogic_ddrAAxi4_b_payload_resp;
    end
    if(system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_ready) begin
      system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rData_id <= system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_payload_id;
      system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rData_resp <= system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_payload_resp;
    end
  end

  always @(posedge io_peripheralClk) begin
    io_peripheralReset <= peripheralCd_logic_outputReset;
    if(axiA_rready) begin
      axiA_r_rData_data <= axiA_rdata;
      axiA_r_rData_id <= axiA_rid;
      axiA_r_rData_resp <= axiA_rresp;
      axiA_r_rData_last <= axiA_rlast;
    end
    if(system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context;
    end
    if(_zz_io_input_rsp_ready_3) begin
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_2 <= _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last;
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source_1 <= _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source;
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode_1 <= _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode;
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data_1 <= _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data;
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context_1 <= _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context;
    end
    if(_zz_2) begin
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_3 <= (_zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 ? _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last : _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_2);
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source_2 <= (_zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 ? _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source : _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source_1);
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode_2 <= (_zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 ? _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode : _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode_1);
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data_2 <= (_zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 ? _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data : _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data_1);
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context_2 <= (_zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 ? _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context : _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context_1);
    end
    if(_zz_io_input_rsp_ready_4) begin
      _zz_system_bmbPeripheral_bmb_rsp_payload_last <= system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_last;
      _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_opcode <= system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_opcode;
      _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_data <= system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_data;
      _zz_system_bmbPeripheral_bmb_rsp_payload_fragment_context <= system_bmbPeripheral_bmb_decoder_io_input_rsp_payload_fragment_context;
    end
    if(system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(_zz_io_bus_rsp_ready_1) begin
      _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last <= system_uart_0_io_logic_io_bus_rsp_payload_last;
      _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode <= system_uart_0_io_logic_io_bus_rsp_payload_fragment_opcode;
      _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data <= system_uart_0_io_logic_io_bus_rsp_payload_fragment_data;
      _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context <= system_uart_0_io_logic_io_bus_rsp_payload_fragment_context;
    end
    if(system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(_zz_system_plic_logic_bus_rsp_ready_1) begin
      _zz_system_plic_logic_bmb_rsp_payload_last <= system_plic_logic_bus_rsp_payload_last;
      _zz_system_plic_logic_bmb_rsp_payload_fragment_opcode <= system_plic_logic_bus_rsp_payload_fragment_opcode;
      _zz_system_plic_logic_bmb_rsp_payload_fragment_data <= system_plic_logic_bus_rsp_payload_fragment_data;
      _zz_system_plic_logic_bmb_rsp_payload_fragment_context <= system_plic_logic_bus_rsp_payload_fragment_context;
    end
    system_cores_0_externalInterrupt_plic_target_bestRequest_priority <= (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_3 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_2 : system_cores_0_externalInterrupt_plic_target_requests_16_priority);
    system_cores_0_externalInterrupt_plic_target_bestRequest_id <= (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_3 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_40 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_36 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_24 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id ? system_cores_0_externalInterrupt_plic_target_requests_0_id : system_cores_0_externalInterrupt_plic_target_requests_1_id) : (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_3 ? system_cores_0_externalInterrupt_plic_target_requests_2_id : system_cores_0_externalInterrupt_plic_target_requests_3_id)) : (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_27 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_6 ? system_cores_0_externalInterrupt_plic_target_requests_4_id : system_cores_0_externalInterrupt_plic_target_requests_5_id) : (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_9 ? system_cores_0_externalInterrupt_plic_target_requests_6_id : system_cores_0_externalInterrupt_plic_target_requests_7_id))) : (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_38 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_30 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_12 ? system_cores_0_externalInterrupt_plic_target_requests_8_id : system_cores_0_externalInterrupt_plic_target_requests_9_id) : (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_15 ? system_cores_0_externalInterrupt_plic_target_requests_10_id : system_cores_0_externalInterrupt_plic_target_requests_11_id)) : (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_33 ? (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_18 ? system_cores_0_externalInterrupt_plic_target_requests_12_id : system_cores_0_externalInterrupt_plic_target_requests_13_id) : (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_id_21 ? system_cores_0_externalInterrupt_plic_target_requests_14_id : system_cores_0_externalInterrupt_plic_target_requests_15_id)))) : system_cores_0_externalInterrupt_plic_target_requests_16_id);
    system_cores_0_externalInterrupt_plic_target_bestRequest_valid <= (_zz_system_cores_0_externalInterrupt_plic_target_bestRequest_priority_3 ? _zz_system_cores_0_externalInterrupt_plic_target_bestRequest_valid : system_cores_0_externalInterrupt_plic_target_requests_16_valid);
    system_cores_1_externalInterrupt_plic_target_bestRequest_priority <= (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_3 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_2 : system_cores_1_externalInterrupt_plic_target_requests_16_priority);
    system_cores_1_externalInterrupt_plic_target_bestRequest_id <= (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_3 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_40 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_36 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_24 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id ? system_cores_1_externalInterrupt_plic_target_requests_0_id : system_cores_1_externalInterrupt_plic_target_requests_1_id) : (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_3 ? system_cores_1_externalInterrupt_plic_target_requests_2_id : system_cores_1_externalInterrupt_plic_target_requests_3_id)) : (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_27 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_6 ? system_cores_1_externalInterrupt_plic_target_requests_4_id : system_cores_1_externalInterrupt_plic_target_requests_5_id) : (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_9 ? system_cores_1_externalInterrupt_plic_target_requests_6_id : system_cores_1_externalInterrupt_plic_target_requests_7_id))) : (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_38 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_30 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_12 ? system_cores_1_externalInterrupt_plic_target_requests_8_id : system_cores_1_externalInterrupt_plic_target_requests_9_id) : (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_15 ? system_cores_1_externalInterrupt_plic_target_requests_10_id : system_cores_1_externalInterrupt_plic_target_requests_11_id)) : (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_33 ? (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_18 ? system_cores_1_externalInterrupt_plic_target_requests_12_id : system_cores_1_externalInterrupt_plic_target_requests_13_id) : (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_id_21 ? system_cores_1_externalInterrupt_plic_target_requests_14_id : system_cores_1_externalInterrupt_plic_target_requests_15_id)))) : system_cores_1_externalInterrupt_plic_target_requests_16_id);
    system_cores_1_externalInterrupt_plic_target_bestRequest_valid <= (_zz_system_cores_1_externalInterrupt_plic_target_bestRequest_priority_3 ? _zz_system_cores_1_externalInterrupt_plic_target_bestRequest_valid : system_cores_1_externalInterrupt_plic_target_requests_16_valid);
    system_cores_0_externalInterrupt_plic_target_iep_regNext <= system_cores_0_externalInterrupt_plic_target_iep;
    system_cores_1_externalInterrupt_plic_target_iep_regNext <= system_cores_1_externalInterrupt_plic_target_iep;
  end

  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      userInterruptA_interrupt_plic_gateway_ip <= 1'b0;
      userInterruptA_interrupt_plic_gateway_waitCompletion <= 1'b0;
      userInterruptD_interrupt_plic_gateway_ip <= 1'b0;
      userInterruptD_interrupt_plic_gateway_waitCompletion <= 1'b0;
      userInterruptC_interrupt_plic_gateway_ip <= 1'b0;
      userInterruptC_interrupt_plic_gateway_waitCompletion <= 1'b0;
      userInterruptB_interrupt_plic_gateway_ip <= 1'b0;
      userInterruptB_interrupt_plic_gateway_waitCompletion <= 1'b0;
      axiA_r_rValid <= 1'b0;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b1;
      system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid <= 1'b0;
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 <= 1'b1;
      _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_2 <= 1'b0;
      system_axiA_interrupt_plic_gateway_ip <= 1'b0;
      system_axiA_interrupt_plic_gateway_waitCompletion <= 1'b0;
      _zz_system_bmbPeripheral_bmb_rsp_valid_1 <= 1'b0;
      system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= 1'b0;
      system_uart_0_io_interrupt_plic_gateway_ip <= 1'b0;
      system_uart_0_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
      system_spi_0_io_interrupt_plic_gateway_ip <= 1'b0;
      system_spi_0_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
      system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      system_spi_1_io_interrupt_plic_gateway_ip <= 1'b0;
      system_spi_1_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
      system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      system_i2c_0_io_interrupt_plic_gateway_ip <= 1'b0;
      system_i2c_0_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
      system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      system_i2c_2_io_interrupt_plic_gateway_ip <= 1'b0;
      system_i2c_2_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
      system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      system_i2c_1_io_interrupt_plic_gateway_ip <= 1'b0;
      system_i2c_1_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
      system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      system_userTimer_1_interrupts_0_plic_gateway_ip <= 1'b0;
      system_userTimer_1_interrupts_0_plic_gateway_waitCompletion <= 1'b0;
      system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      system_userTimer_0_interrupts_0_plic_gateway_ip <= 1'b0;
      system_userTimer_0_interrupts_0_plic_gateway_waitCompletion <= 1'b0;
      system_gpio_0_io_interrupts_0_plic_gateway_ip <= 1'b0;
      system_gpio_0_io_interrupts_0_plic_gateway_waitCompletion <= 1'b0;
      system_gpio_0_io_interrupts_1_plic_gateway_ip <= 1'b0;
      system_gpio_0_io_interrupts_1_plic_gateway_waitCompletion <= 1'b0;
      system_watchdog_logic_panics_0_plic_gateway_ip <= 1'b0;
      system_watchdog_logic_panics_0_plic_gateway_waitCompletion <= 1'b0;
      _zz_system_plic_logic_bmb_rsp_valid_1 <= 1'b0;
      _zz_userInterruptA_interrupt_plic_gateway_priority <= 2'b00;
      _zz_userInterruptD_interrupt_plic_gateway_priority <= 2'b00;
      _zz_userInterruptC_interrupt_plic_gateway_priority <= 2'b00;
      _zz_userInterruptB_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_axiA_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_uart_0_io_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_spi_0_io_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_spi_1_io_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_i2c_0_io_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_i2c_2_io_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_i2c_1_io_interrupt_plic_gateway_priority <= 2'b00;
      _zz_system_userTimer_1_interrupts_0_plic_gateway_priority <= 2'b00;
      _zz_system_userTimer_0_interrupts_0_plic_gateway_priority <= 2'b00;
      _zz_system_gpio_0_io_interrupts_0_plic_gateway_priority <= 2'b00;
      _zz_system_gpio_0_io_interrupts_1_plic_gateway_priority <= 2'b00;
      _zz_system_watchdog_logic_panics_0_plic_gateway_priority <= 2'b00;
      system_plic_logic_bridge_coherencyStall_value <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_threshold <= 2'b00;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_0 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_1 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_2 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_3 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_4 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_5 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_6 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_7 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_8 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_9 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_10 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_11 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_12 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_13 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_14 <= 1'b0;
      _zz_system_cores_0_externalInterrupt_plic_target_ie_15 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_threshold <= 2'b00;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_0 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_1 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_2 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_3 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_4 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_5 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_6 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_7 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_8 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_9 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_10 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_11 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_12 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_13 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_14 <= 1'b0;
      _zz_system_cores_1_externalInterrupt_plic_target_ie_15 <= 1'b0;
    end else begin
      if(when_PlicGateway_l21) begin
        userInterruptA_interrupt_plic_gateway_ip <= userInterruptA_interrupt;
        userInterruptA_interrupt_plic_gateway_waitCompletion <= userInterruptA_interrupt;
      end
      if(when_PlicGateway_l21_1) begin
        userInterruptD_interrupt_plic_gateway_ip <= userInterruptD_interrupt;
        userInterruptD_interrupt_plic_gateway_waitCompletion <= userInterruptD_interrupt;
      end
      if(when_PlicGateway_l21_2) begin
        userInterruptC_interrupt_plic_gateway_ip <= userInterruptC_interrupt;
        userInterruptC_interrupt_plic_gateway_waitCompletion <= userInterruptC_interrupt;
      end
      if(when_PlicGateway_l21_3) begin
        userInterruptB_interrupt_plic_gateway_ip <= userInterruptB_interrupt;
        userInterruptB_interrupt_plic_gateway_waitCompletion <= userInterruptB_interrupt;
      end
      if(axiA_rready) begin
        axiA_r_rValid <= axiA_rvalid;
      end
      if(system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b0;
      end
      if(system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
        system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b1;
      end
      if(system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
        system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid <= system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid;
      end
      if(_zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid) begin
        _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 <= 1'b0;
      end
      if(_zz_2) begin
        _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1 <= 1'b1;
      end
      if(_zz_2) begin
        _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_2 <= (_zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid || (! _zz_system_axiA_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last_1));
      end
      if(when_PlicGateway_l21_4) begin
        system_axiA_interrupt_plic_gateway_ip <= axiAInterrupt;
        system_axiA_interrupt_plic_gateway_waitCompletion <= axiAInterrupt;
      end
      if(system_bmbPeripheral_bmb_decoder_io_input_rsp_valid) begin
        _zz_system_bmbPeripheral_bmb_rsp_valid_1 <= 1'b1;
      end
      if((_zz_system_bmbPeripheral_bmb_rsp_valid && system_bmbPeripheral_bmb_rsp_ready)) begin
        _zz_system_bmbPeripheral_bmb_rsp_valid_1 <= 1'b0;
      end
      if(system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(system_uart_0_io_logic_io_bus_rsp_valid) begin
        _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= 1'b1;
      end
      if((_zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid && system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_ready)) begin
        _zz_system_uart_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= 1'b0;
      end
      if(when_PlicGateway_l21_5) begin
        system_uart_0_io_interrupt_plic_gateway_ip <= system_uart_0_io_logic_io_interrupt;
        system_uart_0_io_interrupt_plic_gateway_waitCompletion <= system_uart_0_io_logic_io_interrupt;
      end
      if(when_PlicGateway_l21_6) begin
        system_spi_0_io_interrupt_plic_gateway_ip <= system_spi_0_io_logic_io_interrupt;
        system_spi_0_io_interrupt_plic_gateway_waitCompletion <= system_spi_0_io_logic_io_interrupt;
      end
      if(system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_spi_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(when_PlicGateway_l21_7) begin
        system_spi_1_io_interrupt_plic_gateway_ip <= system_spi_1_io_logic_io_interrupt;
        system_spi_1_io_interrupt_plic_gateway_waitCompletion <= system_spi_1_io_logic_io_interrupt;
      end
      if(system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_spi_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_i2c_0_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(when_PlicGateway_l21_8) begin
        system_i2c_0_io_interrupt_plic_gateway_ip <= system_i2c_0_io_logic_io_interrupt;
        system_i2c_0_io_interrupt_plic_gateway_waitCompletion <= system_i2c_0_io_logic_io_interrupt;
      end
      if(system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_i2c_2_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(when_PlicGateway_l21_9) begin
        system_i2c_2_io_interrupt_plic_gateway_ip <= system_i2c_2_io_logic_io_interrupt;
        system_i2c_2_io_interrupt_plic_gateway_waitCompletion <= system_i2c_2_io_logic_io_interrupt;
      end
      if(system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_i2c_1_io_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(when_PlicGateway_l21_10) begin
        system_i2c_1_io_interrupt_plic_gateway_ip <= system_i2c_1_io_logic_io_interrupt;
        system_i2c_1_io_interrupt_plic_gateway_waitCompletion <= system_i2c_1_io_logic_io_interrupt;
      end
      if(system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_userTimer_1_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(when_PlicGateway_l21_11) begin
        system_userTimer_1_interrupts_0_plic_gateway_ip <= system_userTimer_1_interrupts_0;
        system_userTimer_1_interrupts_0_plic_gateway_waitCompletion <= system_userTimer_1_interrupts_0;
      end
      if(system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b1;
      end
      if(system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_halfPipe_fire) begin
        system_userTimer_0_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValid <= 1'b0;
      end
      if(when_PlicGateway_l21_12) begin
        system_userTimer_0_interrupts_0_plic_gateway_ip <= system_userTimer_0_interrupts_0;
        system_userTimer_0_interrupts_0_plic_gateway_waitCompletion <= system_userTimer_0_interrupts_0;
      end
      if(when_PlicGateway_l21_13) begin
        system_gpio_0_io_interrupts_0_plic_gateway_ip <= system_gpio_0_io_interrupts_0;
        system_gpio_0_io_interrupts_0_plic_gateway_waitCompletion <= system_gpio_0_io_interrupts_0;
      end
      if(when_PlicGateway_l21_14) begin
        system_gpio_0_io_interrupts_1_plic_gateway_ip <= system_gpio_0_io_interrupts_1;
        system_gpio_0_io_interrupts_1_plic_gateway_waitCompletion <= system_gpio_0_io_interrupts_1;
      end
      if(when_PlicGateway_l21_15) begin
        system_watchdog_logic_panics_0_plic_gateway_ip <= _zz_system_watchdog_logic_panics_0_plic_gateway_ip;
        system_watchdog_logic_panics_0_plic_gateway_waitCompletion <= _zz_system_watchdog_logic_panics_0_plic_gateway_ip;
      end
      if(_zz_system_plic_logic_bus_rsp_ready_1) begin
        _zz_system_plic_logic_bmb_rsp_valid_1 <= (system_plic_logic_bus_rsp_valid && _zz_system_plic_logic_bus_rsp_ready);
      end
      if(system_plic_logic_bridge_claim_valid) begin
        case(system_plic_logic_bridge_claim_payload)
          6'h10 : begin
            userInterruptA_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h17 : begin
            userInterruptD_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h16 : begin
            userInterruptC_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h11 : begin
            userInterruptB_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h1e : begin
            system_axiA_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h01 : begin
            system_uart_0_io_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h04 : begin
            system_spi_0_io_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h05 : begin
            system_spi_1_io_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h08 : begin
            system_i2c_0_io_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h0a : begin
            system_i2c_2_io_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h09 : begin
            system_i2c_1_io_interrupt_plic_gateway_ip <= 1'b0;
          end
          6'h14 : begin
            system_userTimer_1_interrupts_0_plic_gateway_ip <= 1'b0;
          end
          6'h13 : begin
            system_userTimer_0_interrupts_0_plic_gateway_ip <= 1'b0;
          end
          6'h0c : begin
            system_gpio_0_io_interrupts_0_plic_gateway_ip <= 1'b0;
          end
          6'h0d : begin
            system_gpio_0_io_interrupts_1_plic_gateway_ip <= 1'b0;
          end
          6'h20 : begin
            system_watchdog_logic_panics_0_plic_gateway_ip <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      if(system_plic_logic_bridge_completion_valid) begin
        case(system_plic_logic_bridge_completion_payload)
          6'h10 : begin
            userInterruptA_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h17 : begin
            userInterruptD_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h16 : begin
            userInterruptC_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h11 : begin
            userInterruptB_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h1e : begin
            system_axiA_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h01 : begin
            system_uart_0_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h04 : begin
            system_spi_0_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h05 : begin
            system_spi_1_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h08 : begin
            system_i2c_0_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h0a : begin
            system_i2c_2_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h09 : begin
            system_i2c_1_io_interrupt_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h14 : begin
            system_userTimer_1_interrupts_0_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h13 : begin
            system_userTimer_0_interrupts_0_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h0c : begin
            system_gpio_0_io_interrupts_0_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h0d : begin
            system_gpio_0_io_interrupts_1_plic_gateway_waitCompletion <= 1'b0;
          end
          6'h20 : begin
            system_watchdog_logic_panics_0_plic_gateway_waitCompletion <= 1'b0;
          end
          default : begin
          end
        endcase
      end
      system_plic_logic_bridge_coherencyStall_value <= system_plic_logic_bridge_coherencyStall_valueNext;
      case(system_plic_logic_bmb_cmd_payload_fragment_address)
        22'h000040 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_userInterruptA_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h00005c : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_userInterruptD_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000058 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_userInterruptC_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000044 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_userInterruptB_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000078 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_axiA_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000004 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_uart_0_io_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000010 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_spi_0_io_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000014 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_spi_1_io_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000020 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_i2c_0_io_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000028 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_i2c_2_io_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000024 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_i2c_1_io_interrupt_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000050 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_userTimer_1_interrupts_0_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h00004c : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_userTimer_0_interrupts_0_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000030 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_gpio_0_io_interrupts_0_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000034 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_gpio_0_io_interrupts_1_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h000080 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_watchdog_logic_panics_0_plic_gateway_priority <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h200000 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_cores_0_externalInterrupt_plic_target_threshold <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h002000 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_cores_0_externalInterrupt_plic_target_ie_0 <= system_plic_logic_bmb_cmd_payload_fragment_data[16];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_1 <= system_plic_logic_bmb_cmd_payload_fragment_data[23];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_2 <= system_plic_logic_bmb_cmd_payload_fragment_data[22];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_3 <= system_plic_logic_bmb_cmd_payload_fragment_data[17];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_4 <= system_plic_logic_bmb_cmd_payload_fragment_data[30];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_5 <= system_plic_logic_bmb_cmd_payload_fragment_data[1];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_6 <= system_plic_logic_bmb_cmd_payload_fragment_data[4];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_7 <= system_plic_logic_bmb_cmd_payload_fragment_data[5];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_8 <= system_plic_logic_bmb_cmd_payload_fragment_data[8];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_9 <= system_plic_logic_bmb_cmd_payload_fragment_data[10];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_10 <= system_plic_logic_bmb_cmd_payload_fragment_data[9];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_11 <= system_plic_logic_bmb_cmd_payload_fragment_data[20];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_12 <= system_plic_logic_bmb_cmd_payload_fragment_data[19];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_13 <= system_plic_logic_bmb_cmd_payload_fragment_data[12];
            _zz_system_cores_0_externalInterrupt_plic_target_ie_14 <= system_plic_logic_bmb_cmd_payload_fragment_data[13];
          end
        end
        22'h002004 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_cores_0_externalInterrupt_plic_target_ie_15 <= system_plic_logic_bmb_cmd_payload_fragment_data[0];
          end
        end
        22'h201000 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_cores_1_externalInterrupt_plic_target_threshold <= system_plic_logic_bmb_cmd_payload_fragment_data[1 : 0];
          end
        end
        22'h002080 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_cores_1_externalInterrupt_plic_target_ie_0 <= system_plic_logic_bmb_cmd_payload_fragment_data[16];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_1 <= system_plic_logic_bmb_cmd_payload_fragment_data[23];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_2 <= system_plic_logic_bmb_cmd_payload_fragment_data[22];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_3 <= system_plic_logic_bmb_cmd_payload_fragment_data[17];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_4 <= system_plic_logic_bmb_cmd_payload_fragment_data[30];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_5 <= system_plic_logic_bmb_cmd_payload_fragment_data[1];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_6 <= system_plic_logic_bmb_cmd_payload_fragment_data[4];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_7 <= system_plic_logic_bmb_cmd_payload_fragment_data[5];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_8 <= system_plic_logic_bmb_cmd_payload_fragment_data[8];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_9 <= system_plic_logic_bmb_cmd_payload_fragment_data[10];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_10 <= system_plic_logic_bmb_cmd_payload_fragment_data[9];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_11 <= system_plic_logic_bmb_cmd_payload_fragment_data[20];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_12 <= system_plic_logic_bmb_cmd_payload_fragment_data[19];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_13 <= system_plic_logic_bmb_cmd_payload_fragment_data[12];
            _zz_system_cores_1_externalInterrupt_plic_target_ie_14 <= system_plic_logic_bmb_cmd_payload_fragment_data[13];
          end
        end
        22'h002084 : begin
          if(system_plic_logic_bus_doWrite) begin
            _zz_system_cores_1_externalInterrupt_plic_target_ie_15 <= system_plic_logic_bmb_cmd_payload_fragment_data[0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid <= 1'b0;
      dBus_Bridge_withWriteBuffer_buffer_mask <= 8'h0;
      dBus_Bridge_withWriteBuffer_aggregationCounter <= 4'b0000;
      dBus_Bridge_withWriteBuffer_timer <= 6'h0;
      io_pop_rValidN <= 1'b1;
      io_pop_s2mPipe_rValid <= 1'b0;
      _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid_1 <= 1'b0;
      dBus_Bridge_withWriteBuffer_buffer_mask_1 <= 8'h0;
      dBus_Bridge_withWriteBuffer_aggregationCounter_1 <= 4'b0000;
      dBus_Bridge_withWriteBuffer_timer_1 <= 6'h0;
      io_pop_rValidN_1 <= 1'b1;
      io_pop_s2mPipe_rValid_1 <= 1'b0;
      _zz_system_cores_0_iBus_rsp_valid_1 <= 1'b0;
      _zz_system_cores_1_iBus_rsp_valid_1 <= 1'b0;
      dBus_Bridge_bus_cmd_rValid <= 1'b0;
      _zz_dBus_Bridge_bus_inv_valid_1 <= 1'b0;
      dBus_Bridge_bus_ack_rValid <= 1'b0;
      _zz_dBus_Bridge_bus_sync_valid_1 <= 1'b0;
      dBus_Bridge_bus_cmd_rValid_1 <= 1'b0;
      _zz_dBus_Bridge_bus_inv_valid_3 <= 1'b0;
      dBus_Bridge_bus_ack_rValid_1 <= 1'b0;
      _zz_dBus_Bridge_bus_sync_valid_3 <= 1'b0;
      FpuPlugin_port_commit_rValid <= 1'b0;
      io_port_0_completion_regNext_valid <= 1'b0;
      io_port_0_rsp_rValidN <= 1'b1;
      FpuPlugin_port_commit_rValid_1 <= 1'b0;
      io_port_1_completion_regNext_valid <= 1'b0;
      io_port_1_rsp_rValidN <= 1'b1;
      _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1 <= 1'b1;
      system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_rValid <= 1'b0;
      io_output_cmd_rValidN <= 1'b1;
      io_output_cmd_s2mPipe_rValid <= 1'b0;
      _zz_when_Stream_l375_1 <= 1'b0;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b1;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid <= 1'b0;
      _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= 1'b0;
      system_fabric_iBus_bmb_cmd_rValid <= 1'b0;
      system_bridge_bmb_cmd_rValidN <= 1'b1;
      system_bridge_bmb_cmd_s2mPipe_rValid <= 1'b0;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b1;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid <= 1'b0;
      _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= 1'b0;
      _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= 1'b0;
    end else begin
      if(_zz_dBus_cmd_ready) begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid <= system_cores_0_logic_cpu_dBus_cmd_valid;
      end
      if(dBus_cmd_fire) begin
        dBus_Bridge_withWriteBuffer_aggregationCounter <= (dBus_Bridge_withWriteBuffer_aggregationCounter + 4'b0001);
      end
      if(when_DataCache_l465) begin
        dBus_Bridge_withWriteBuffer_timer <= (dBus_Bridge_withWriteBuffer_timer + 6'h01);
      end
      if(when_DataCache_l468) begin
        dBus_Bridge_withWriteBuffer_buffer_mask <= 8'h0;
        dBus_Bridge_withWriteBuffer_aggregationCounter <= 4'b0000;
        dBus_Bridge_withWriteBuffer_timer <= 6'h0;
      end
      if(dBus_cmd_fire) begin
        if(when_DataCache_l493) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[0] <= 1'b1;
        end
        if(when_DataCache_l493_1) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[1] <= 1'b1;
        end
        if(when_DataCache_l493_2) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[2] <= 1'b1;
        end
        if(when_DataCache_l493_3) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[3] <= 1'b1;
        end
        if(when_DataCache_l493_4) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[4] <= 1'b1;
        end
        if(when_DataCache_l493_5) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[5] <= 1'b1;
        end
        if(when_DataCache_l493_6) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[6] <= 1'b1;
        end
        if(when_DataCache_l493_7) begin
          dBus_Bridge_withWriteBuffer_buffer_mask[7] <= 1'b1;
        end
      end
      if(dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_valid) begin
        io_pop_rValidN <= 1'b0;
      end
      if(io_pop_s2mPipe_ready) begin
        io_pop_rValidN <= 1'b1;
      end
      if(io_pop_s2mPipe_ready) begin
        io_pop_s2mPipe_rValid <= io_pop_s2mPipe_valid;
      end
      if(_zz_dBus_cmd_ready_1) begin
        _zz_dBus_Bridge_withWriteBuffer_buffer_stream_valid_1 <= system_cores_1_logic_cpu_dBus_cmd_valid;
      end
      if(dBus_cmd_fire_1) begin
        dBus_Bridge_withWriteBuffer_aggregationCounter_1 <= (dBus_Bridge_withWriteBuffer_aggregationCounter_1 + 4'b0001);
      end
      if(when_DataCache_l465_1) begin
        dBus_Bridge_withWriteBuffer_timer_1 <= (dBus_Bridge_withWriteBuffer_timer_1 + 6'h01);
      end
      if(when_DataCache_l468_1) begin
        dBus_Bridge_withWriteBuffer_buffer_mask_1 <= 8'h0;
        dBus_Bridge_withWriteBuffer_aggregationCounter_1 <= 4'b0000;
        dBus_Bridge_withWriteBuffer_timer_1 <= 6'h0;
      end
      if(dBus_cmd_fire_1) begin
        if(when_DataCache_l493_8) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[0] <= 1'b1;
        end
        if(when_DataCache_l493_9) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[1] <= 1'b1;
        end
        if(when_DataCache_l493_10) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[2] <= 1'b1;
        end
        if(when_DataCache_l493_11) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[3] <= 1'b1;
        end
        if(when_DataCache_l493_12) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[4] <= 1'b1;
        end
        if(when_DataCache_l493_13) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[5] <= 1'b1;
        end
        if(when_DataCache_l493_14) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[6] <= 1'b1;
        end
        if(when_DataCache_l493_15) begin
          dBus_Bridge_withWriteBuffer_buffer_mask_1[7] <= 1'b1;
        end
      end
      if(dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_valid) begin
        io_pop_rValidN_1 <= 1'b0;
      end
      if(io_pop_s2mPipe_ready_1) begin
        io_pop_rValidN_1 <= 1'b1;
      end
      if(io_pop_s2mPipe_ready_1) begin
        io_pop_s2mPipe_rValid_1 <= io_pop_s2mPipe_valid_1;
      end
      if(_zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready) begin
        _zz_system_cores_0_iBus_rsp_valid_1 <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_valid;
      end
      if(_zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready) begin
        _zz_system_cores_1_iBus_rsp_valid_1 <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_valid;
      end
      if(dBus_Bridge_bus_cmd_ready) begin
        dBus_Bridge_bus_cmd_rValid <= dBus_Bridge_bus_cmd_valid;
      end
      if(_zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready) begin
        _zz_dBus_Bridge_bus_inv_valid_1 <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_valid;
      end
      if(dBus_Bridge_bus_ack_ready) begin
        dBus_Bridge_bus_ack_rValid <= dBus_Bridge_bus_ack_valid;
      end
      if(_zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_ready) begin
        _zz_dBus_Bridge_bus_sync_valid_1 <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_sync_valid;
      end
      if(dBus_Bridge_bus_cmd_ready_1) begin
        dBus_Bridge_bus_cmd_rValid_1 <= dBus_Bridge_bus_cmd_valid_1;
      end
      if(_zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready) begin
        _zz_dBus_Bridge_bus_inv_valid_3 <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_valid;
      end
      if(dBus_Bridge_bus_ack_ready_1) begin
        dBus_Bridge_bus_ack_rValid_1 <= dBus_Bridge_bus_ack_valid_1;
      end
      if(_zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_ready) begin
        _zz_dBus_Bridge_bus_sync_valid_3 <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_sync_valid;
      end
      if(system_cores_0_logic_cpu_FpuPlugin_port_commit_ready) begin
        FpuPlugin_port_commit_rValid <= system_cores_0_logic_cpu_FpuPlugin_port_commit_valid;
      end
      io_port_0_completion_regNext_valid <= system_fpu_logic_io_port_0_completion_valid;
      if(system_fpu_logic_io_port_0_rsp_valid) begin
        io_port_0_rsp_rValidN <= 1'b0;
      end
      if(io_port_0_rsp_s2mPipe_ready) begin
        io_port_0_rsp_rValidN <= 1'b1;
      end
      if(system_cores_1_logic_cpu_FpuPlugin_port_commit_ready) begin
        FpuPlugin_port_commit_rValid_1 <= system_cores_1_logic_cpu_FpuPlugin_port_commit_valid;
      end
      io_port_1_completion_regNext_valid <= system_fpu_logic_io_port_1_completion_valid;
      if(system_fpu_logic_io_port_1_rsp_valid) begin
        io_port_1_rsp_rValidN <= 1'b0;
      end
      if(io_port_1_rsp_s2mPipe_ready) begin
        io_port_1_rsp_rValidN <= 1'b1;
      end
      if(_zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid) begin
        _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1 <= 1'b0;
      end
      if(system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_ready) begin
        _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_valid_1 <= 1'b1;
      end
      if(system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_ready) begin
        system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_rValid <= system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_ack_valid;
      end
      if(system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_valid) begin
        io_output_cmd_rValidN <= 1'b0;
      end
      if(io_output_cmd_s2mPipe_ready) begin
        io_output_cmd_rValidN <= 1'b1;
      end
      if(io_output_cmd_s2mPipe_ready) begin
        io_output_cmd_s2mPipe_rValid <= io_output_cmd_s2mPipe_valid;
      end
      if(_zz_system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready) begin
        _zz_when_Stream_l375_1 <= system_fabric_invalidationMonitor_output_connector_decoder_rsp_valid;
      end
      if(system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b0;
      end
      if(system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
        system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b1;
      end
      if(system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
        system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid;
      end
      if(_zz_io_input_rsp_ready) begin
        _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= system_fabric_exclusiveMonitor_logic_io_input_rsp_valid;
      end
      if(system_fabric_iBus_bmb_cmd_ready) begin
        system_fabric_iBus_bmb_cmd_rValid <= system_fabric_iBus_bmb_cmd_valid;
      end
      if(system_bridge_bmb_cmd_valid) begin
        system_bridge_bmb_cmd_rValidN <= 1'b0;
      end
      if(system_bridge_bmb_cmd_s2mPipe_ready) begin
        system_bridge_bmb_cmd_rValidN <= 1'b1;
      end
      if(system_bridge_bmb_cmd_s2mPipe_ready) begin
        system_bridge_bmb_cmd_s2mPipe_rValid <= system_bridge_bmb_cmd_s2mPipe_valid;
      end
      if(system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_valid) begin
        system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b0;
      end
      if(system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
        system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rValidN <= 1'b1;
      end
      if(system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
        system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rValid <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_valid;
      end
      if(_zz_io_input_rsp_ready_2) begin
        _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= system_ddr_ddrLogic_cc_fifo_io_input_rsp_valid;
      end
      if(_zz_io_bus_rsp_ready) begin
        _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_valid_1 <= system_ramA_logic_io_bus_rsp_valid;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(dBus_cmd_fire) begin
      if(when_DataCache_l493) begin
        dBus_Bridge_withWriteBuffer_buffer_data[7 : 0] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[7 : 0];
      end
      if(when_DataCache_l493_1) begin
        dBus_Bridge_withWriteBuffer_buffer_data[15 : 8] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[15 : 8];
      end
      if(when_DataCache_l493_2) begin
        dBus_Bridge_withWriteBuffer_buffer_data[23 : 16] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[23 : 16];
      end
      if(when_DataCache_l493_3) begin
        dBus_Bridge_withWriteBuffer_buffer_data[31 : 24] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[31 : 24];
      end
      if(when_DataCache_l493_4) begin
        dBus_Bridge_withWriteBuffer_buffer_data[39 : 32] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[39 : 32];
      end
      if(when_DataCache_l493_5) begin
        dBus_Bridge_withWriteBuffer_buffer_data[47 : 40] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[47 : 40];
      end
      if(when_DataCache_l493_6) begin
        dBus_Bridge_withWriteBuffer_buffer_data[55 : 48] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[55 : 48];
      end
      if(when_DataCache_l493_7) begin
        dBus_Bridge_withWriteBuffer_buffer_data[63 : 56] <= system_cores_0_logic_cpu_dBus_cmd_payload_data[63 : 56];
      end
    end
    if(dBus_cmd_fire) begin
      dBus_Bridge_withWriteBuffer_buffer_write <= system_cores_0_logic_cpu_dBus_cmd_payload_wr;
      dBus_Bridge_withWriteBuffer_buffer_address <= system_cores_0_logic_cpu_dBus_cmd_payload_address;
      dBus_Bridge_withWriteBuffer_buffer_length <= _zz_dBus_Bridge_withWriteBuffer_buffer_length;
      dBus_Bridge_withWriteBuffer_buffer_exclusive <= system_cores_0_logic_cpu_dBus_cmd_payload_exclusive;
      if(when_DataCache_l506) begin
        dBus_Bridge_withWriteBuffer_aggregationEnabled <= 1'b1;
        dBus_Bridge_withWriteBuffer_buffer_address[2 : 0] <= 3'b000;
        dBus_Bridge_withWriteBuffer_buffer_length <= 6'h07;
      end else begin
        dBus_Bridge_withWriteBuffer_aggregationEnabled <= 1'b0;
      end
    end
    if(io_pop_rValidN) begin
      io_pop_rData <= dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_io_pop_payload;
    end
    if(io_pop_s2mPipe_ready) begin
      io_pop_s2mPipe_rData <= io_pop_s2mPipe_payload;
    end
    if(dBus_cmd_fire_1) begin
      if(when_DataCache_l493_8) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[7 : 0] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[7 : 0];
      end
      if(when_DataCache_l493_9) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[15 : 8] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[15 : 8];
      end
      if(when_DataCache_l493_10) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[23 : 16] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[23 : 16];
      end
      if(when_DataCache_l493_11) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[31 : 24] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[31 : 24];
      end
      if(when_DataCache_l493_12) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[39 : 32] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[39 : 32];
      end
      if(when_DataCache_l493_13) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[47 : 40] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[47 : 40];
      end
      if(when_DataCache_l493_14) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[55 : 48] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[55 : 48];
      end
      if(when_DataCache_l493_15) begin
        dBus_Bridge_withWriteBuffer_buffer_data_1[63 : 56] <= system_cores_1_logic_cpu_dBus_cmd_payload_data[63 : 56];
      end
    end
    if(dBus_cmd_fire_1) begin
      dBus_Bridge_withWriteBuffer_buffer_write_1 <= system_cores_1_logic_cpu_dBus_cmd_payload_wr;
      dBus_Bridge_withWriteBuffer_buffer_address_1 <= system_cores_1_logic_cpu_dBus_cmd_payload_address;
      dBus_Bridge_withWriteBuffer_buffer_length_1 <= _zz_dBus_Bridge_withWriteBuffer_buffer_length_1;
      dBus_Bridge_withWriteBuffer_buffer_exclusive_1 <= system_cores_1_logic_cpu_dBus_cmd_payload_exclusive;
      if(when_DataCache_l506_1) begin
        dBus_Bridge_withWriteBuffer_aggregationEnabled_1 <= 1'b1;
        dBus_Bridge_withWriteBuffer_buffer_address_1[2 : 0] <= 3'b000;
        dBus_Bridge_withWriteBuffer_buffer_length_1 <= 6'h07;
      end else begin
        dBus_Bridge_withWriteBuffer_aggregationEnabled_1 <= 1'b0;
      end
    end
    if(io_pop_rValidN_1) begin
      io_pop_rData_1 <= dBus_Bridge_withWriteBuffer_syncLogic_cmdCtx_fifo_1_io_pop_payload;
    end
    if(io_pop_s2mPipe_ready_1) begin
      io_pop_s2mPipe_rData_1 <= io_pop_s2mPipe_payload_1;
    end
    io_systemReset <= systemCd_logic_outputReset;
    if(_zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_ready) begin
      _zz_system_cores_0_iBus_rsp_payload_last <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_last;
      _zz_system_cores_0_iBus_rsp_payload_fragment_opcode <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_opcode;
      _zz_system_cores_0_iBus_rsp_payload_fragment_data <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_rsp_payload_fragment_data;
    end
    if(_zz_system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_ready) begin
      _zz_system_cores_1_iBus_rsp_payload_last <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_last;
      _zz_system_cores_1_iBus_rsp_payload_fragment_opcode <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_opcode;
      _zz_system_cores_1_iBus_rsp_payload_fragment_data <= system_fabric_iBus_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_rsp_payload_fragment_data;
    end
    if(dBus_Bridge_bus_cmd_ready) begin
      dBus_Bridge_bus_cmd_rData_last <= dBus_Bridge_bus_cmd_payload_last;
      dBus_Bridge_bus_cmd_rData_fragment_opcode <= dBus_Bridge_bus_cmd_payload_fragment_opcode;
      dBus_Bridge_bus_cmd_rData_fragment_exclusive <= dBus_Bridge_bus_cmd_payload_fragment_exclusive;
      dBus_Bridge_bus_cmd_rData_fragment_address <= dBus_Bridge_bus_cmd_payload_fragment_address;
      dBus_Bridge_bus_cmd_rData_fragment_length <= dBus_Bridge_bus_cmd_payload_fragment_length;
      dBus_Bridge_bus_cmd_rData_fragment_data <= dBus_Bridge_bus_cmd_payload_fragment_data;
      dBus_Bridge_bus_cmd_rData_fragment_mask <= dBus_Bridge_bus_cmd_payload_fragment_mask;
      dBus_Bridge_bus_cmd_rData_fragment_context <= dBus_Bridge_bus_cmd_payload_fragment_context;
    end
    if(_zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_ready) begin
      _zz_dBus_Bridge_bus_inv_payload_all <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_all;
      _zz_dBus_Bridge_bus_inv_payload_address <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_address;
      _zz_dBus_Bridge_bus_inv_payload_length <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_1_decoder_inv_payload_length;
    end
    if(dBus_Bridge_bus_cmd_ready_1) begin
      dBus_Bridge_bus_cmd_rData_last_1 <= dBus_Bridge_bus_cmd_payload_last_1;
      dBus_Bridge_bus_cmd_rData_fragment_opcode_1 <= dBus_Bridge_bus_cmd_payload_fragment_opcode_1;
      dBus_Bridge_bus_cmd_rData_fragment_exclusive_1 <= dBus_Bridge_bus_cmd_payload_fragment_exclusive_1;
      dBus_Bridge_bus_cmd_rData_fragment_address_1 <= dBus_Bridge_bus_cmd_payload_fragment_address_1;
      dBus_Bridge_bus_cmd_rData_fragment_length_1 <= dBus_Bridge_bus_cmd_payload_fragment_length_1;
      dBus_Bridge_bus_cmd_rData_fragment_data_1 <= dBus_Bridge_bus_cmd_payload_fragment_data_1;
      dBus_Bridge_bus_cmd_rData_fragment_mask_1 <= dBus_Bridge_bus_cmd_payload_fragment_mask_1;
      dBus_Bridge_bus_cmd_rData_fragment_context_1 <= dBus_Bridge_bus_cmd_payload_fragment_context_1;
    end
    if(_zz_system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_ready) begin
      _zz_dBus_Bridge_bus_inv_payload_all_1 <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_all;
      _zz_dBus_Bridge_bus_inv_payload_address_1 <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_address;
      _zz_dBus_Bridge_bus_inv_payload_length_1 <= system_fabric_dBusCoherent_bmb_slaveModel_arbiterGen_logic_sorted_0_decoder_inv_payload_length;
    end
    if(system_cores_0_logic_cpu_FpuPlugin_port_commit_ready) begin
      FpuPlugin_port_commit_rData_opcode <= system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_opcode;
      FpuPlugin_port_commit_rData_rd <= system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_rd;
      FpuPlugin_port_commit_rData_write <= system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_write;
      FpuPlugin_port_commit_rData_value <= system_cores_0_logic_cpu_FpuPlugin_port_commit_payload_value;
    end
    io_port_0_completion_regNext_payload_flags_NX <= system_fpu_logic_io_port_0_completion_payload_flags_NX;
    io_port_0_completion_regNext_payload_flags_UF <= system_fpu_logic_io_port_0_completion_payload_flags_UF;
    io_port_0_completion_regNext_payload_flags_OF <= system_fpu_logic_io_port_0_completion_payload_flags_OF;
    io_port_0_completion_regNext_payload_flags_DZ <= system_fpu_logic_io_port_0_completion_payload_flags_DZ;
    io_port_0_completion_regNext_payload_flags_NV <= system_fpu_logic_io_port_0_completion_payload_flags_NV;
    io_port_0_completion_regNext_payload_written <= system_fpu_logic_io_port_0_completion_payload_written;
    if(io_port_0_rsp_rValidN) begin
      io_port_0_rsp_rData_value <= system_fpu_logic_io_port_0_rsp_payload_value;
      io_port_0_rsp_rData_NV <= system_fpu_logic_io_port_0_rsp_payload_NV;
      io_port_0_rsp_rData_NX <= system_fpu_logic_io_port_0_rsp_payload_NX;
    end
    if(system_cores_1_logic_cpu_FpuPlugin_port_commit_ready) begin
      FpuPlugin_port_commit_rData_opcode_1 <= system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_opcode;
      FpuPlugin_port_commit_rData_rd_1 <= system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_rd;
      FpuPlugin_port_commit_rData_write_1 <= system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_write;
      FpuPlugin_port_commit_rData_value_1 <= system_cores_1_logic_cpu_FpuPlugin_port_commit_payload_value;
    end
    io_port_1_completion_regNext_payload_flags_NX <= system_fpu_logic_io_port_1_completion_payload_flags_NX;
    io_port_1_completion_regNext_payload_flags_UF <= system_fpu_logic_io_port_1_completion_payload_flags_UF;
    io_port_1_completion_regNext_payload_flags_OF <= system_fpu_logic_io_port_1_completion_payload_flags_OF;
    io_port_1_completion_regNext_payload_flags_DZ <= system_fpu_logic_io_port_1_completion_payload_flags_DZ;
    io_port_1_completion_regNext_payload_flags_NV <= system_fpu_logic_io_port_1_completion_payload_flags_NV;
    io_port_1_completion_regNext_payload_written <= system_fpu_logic_io_port_1_completion_payload_written;
    if(io_port_1_rsp_rValidN) begin
      io_port_1_rsp_rData_value <= system_fpu_logic_io_port_1_rsp_payload_value;
      io_port_1_rsp_rData_NV <= system_fpu_logic_io_port_1_rsp_payload_NV;
      io_port_1_rsp_rData_NX <= system_fpu_logic_io_port_1_rsp_payload_NX;
    end
    if(_zz_system_fabric_invalidationMonitor_logic_input_inv_ready) begin
      _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all_1 <= _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_all;
      _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address_1 <= _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_address;
      _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length_1 <= _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_length;
      _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source_1 <= _zz_system_fabric_invalidationMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_inv_payload_source;
    end
    if(io_output_cmd_rValidN) begin
      io_output_cmd_rData_last <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_last;
      io_output_cmd_rData_fragment_source <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_source;
      io_output_cmd_rData_fragment_opcode <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_opcode;
      io_output_cmd_rData_fragment_address <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_address;
      io_output_cmd_rData_fragment_length <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_length;
      io_output_cmd_rData_fragment_data <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_data;
      io_output_cmd_rData_fragment_mask <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_mask;
      io_output_cmd_rData_fragment_context <= system_fabric_invalidationMonitor_logic_monitor_io_output_cmd_payload_fragment_context;
    end
    if(io_output_cmd_s2mPipe_ready) begin
      io_output_cmd_s2mPipe_rData_last <= io_output_cmd_s2mPipe_payload_last;
      io_output_cmd_s2mPipe_rData_fragment_source <= io_output_cmd_s2mPipe_payload_fragment_source;
      io_output_cmd_s2mPipe_rData_fragment_opcode <= io_output_cmd_s2mPipe_payload_fragment_opcode;
      io_output_cmd_s2mPipe_rData_fragment_address <= io_output_cmd_s2mPipe_payload_fragment_address;
      io_output_cmd_s2mPipe_rData_fragment_length <= io_output_cmd_s2mPipe_payload_fragment_length;
      io_output_cmd_s2mPipe_rData_fragment_data <= io_output_cmd_s2mPipe_payload_fragment_data;
      io_output_cmd_s2mPipe_rData_fragment_mask <= io_output_cmd_s2mPipe_payload_fragment_mask;
      io_output_cmd_s2mPipe_rData_fragment_context <= io_output_cmd_s2mPipe_payload_fragment_context;
    end
    if(_zz_system_fabric_invalidationMonitor_output_connector_decoder_rsp_ready) begin
      _zz_io_output_rsp_payload_last <= system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_last;
      _zz_io_output_rsp_payload_fragment_source <= system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_source;
      _zz_io_output_rsp_payload_fragment_opcode <= system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_opcode;
      _zz_io_output_rsp_payload_fragment_data <= system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_data;
      _zz_io_output_rsp_payload_fragment_context <= system_fabric_invalidationMonitor_output_connector_decoder_rsp_payload_fragment_context;
    end
    if(system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_exclusive <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_exclusive;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_exclusive <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_exclusive;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask;
      system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context <= system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context;
    end
    if(_zz_io_input_rsp_ready) begin
      _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last <= system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_last;
      _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source <= system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_source;
      _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode <= system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_opcode;
      _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_exclusive <= system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_exclusive;
      _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data <= system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_data;
      _zz_system_fabric_exclusiveMonitor_input_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context <= system_fabric_exclusiveMonitor_logic_io_input_rsp_payload_fragment_context;
    end
    if(system_fabric_iBus_bmb_cmd_ready) begin
      system_fabric_iBus_bmb_cmd_rData_last <= system_fabric_iBus_bmb_cmd_payload_last;
      system_fabric_iBus_bmb_cmd_rData_fragment_source <= system_fabric_iBus_bmb_cmd_payload_fragment_source;
      system_fabric_iBus_bmb_cmd_rData_fragment_opcode <= system_fabric_iBus_bmb_cmd_payload_fragment_opcode;
      system_fabric_iBus_bmb_cmd_rData_fragment_address <= system_fabric_iBus_bmb_cmd_payload_fragment_address;
      system_fabric_iBus_bmb_cmd_rData_fragment_length <= system_fabric_iBus_bmb_cmd_payload_fragment_length;
    end
    if(system_bridge_bmb_cmd_ready) begin
      system_bridge_bmb_cmd_rData_last <= system_bridge_bmb_cmd_payload_last;
      system_bridge_bmb_cmd_rData_fragment_source <= system_bridge_bmb_cmd_payload_fragment_source;
      system_bridge_bmb_cmd_rData_fragment_opcode <= system_bridge_bmb_cmd_payload_fragment_opcode;
      system_bridge_bmb_cmd_rData_fragment_address <= system_bridge_bmb_cmd_payload_fragment_address;
      system_bridge_bmb_cmd_rData_fragment_length <= system_bridge_bmb_cmd_payload_fragment_length;
      system_bridge_bmb_cmd_rData_fragment_data <= system_bridge_bmb_cmd_payload_fragment_data;
      system_bridge_bmb_cmd_rData_fragment_mask <= system_bridge_bmb_cmd_payload_fragment_mask;
      system_bridge_bmb_cmd_rData_fragment_context <= system_bridge_bmb_cmd_payload_fragment_context;
    end
    if(system_bridge_bmb_cmd_s2mPipe_ready) begin
      system_bridge_bmb_cmd_s2mPipe_rData_last <= system_bridge_bmb_cmd_s2mPipe_payload_last;
      system_bridge_bmb_cmd_s2mPipe_rData_fragment_source <= system_bridge_bmb_cmd_s2mPipe_payload_fragment_source;
      system_bridge_bmb_cmd_s2mPipe_rData_fragment_opcode <= system_bridge_bmb_cmd_s2mPipe_payload_fragment_opcode;
      system_bridge_bmb_cmd_s2mPipe_rData_fragment_address <= system_bridge_bmb_cmd_s2mPipe_payload_fragment_address;
      system_bridge_bmb_cmd_s2mPipe_rData_fragment_length <= system_bridge_bmb_cmd_s2mPipe_payload_fragment_length;
      system_bridge_bmb_cmd_s2mPipe_rData_fragment_data <= system_bridge_bmb_cmd_s2mPipe_payload_fragment_data;
      system_bridge_bmb_cmd_s2mPipe_rData_fragment_mask <= system_bridge_bmb_cmd_s2mPipe_payload_fragment_mask;
      system_bridge_bmb_cmd_s2mPipe_rData_fragment_context <= system_bridge_bmb_cmd_s2mPipe_payload_fragment_context;
    end
    if(system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_ready) begin
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_last <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_last;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_source <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_source;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_opcode <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_opcode;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_address <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_address;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_length <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_length;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_data <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_data;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_mask <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_mask;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_rData_fragment_context <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_payload_fragment_context;
    end
    if(system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_ready) begin
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_last <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_last;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_source <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_source;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_opcode <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_opcode;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_address <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_address;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_length <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_length;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_data <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_data;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_mask <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_mask;
      system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_rData_fragment_context <= system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_cmd_s2mPipe_payload_fragment_context;
    end
    if(_zz_io_input_rsp_ready_2) begin
      _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last <= system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_last;
      _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_source <= system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_source;
      _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode <= system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_opcode;
      _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data <= system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_data;
      _zz_system_ddr_bmb_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context <= system_ddr_ddrLogic_cc_fifo_io_input_rsp_payload_fragment_context;
    end
    if(_zz_io_bus_rsp_ready) begin
      _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_last <= system_ramA_logic_io_bus_rsp_payload_last;
      _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_opcode <= system_ramA_logic_io_bus_rsp_payload_fragment_opcode;
      _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_data <= system_ramA_logic_io_bus_rsp_payload_fragment_data;
      _zz_system_ramA_ctrl_slaveModel_arbiterGen_oneToOne_arbiter_rsp_payload_fragment_context <= system_ramA_logic_io_bus_rsp_payload_fragment_context;
    end
  end

  always @(posedge io_systemClk) begin
    if(debugCd_logic_outputReset) begin
      io_harts_0_dmToHart_regNext_valid <= 1'b0;
      io_harts_1_dmToHart_regNext_valid <= 1'b0;
      _zz_1 <= 1'b0;
    end else begin
      io_harts_0_dmToHart_regNext_valid <= system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_valid;
      io_harts_1_dmToHart_regNext_valid <= system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_valid;
      _zz_1 <= (&{system_cores_1_logic_cpu_stoptime,system_cores_0_logic_cpu_stoptime});
    end
  end

  always @(posedge io_systemClk) begin
    io_harts_0_dmToHart_regNext_payload_op <= system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_op;
    io_harts_0_dmToHart_regNext_payload_address <= system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_address;
    io_harts_0_dmToHart_regNext_payload_data <= system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_data;
    io_harts_0_dmToHart_regNext_payload_size <= system_riscvJtag_debug_logic_dm_io_harts_0_dmToHart_payload_size;
    io_harts_1_dmToHart_regNext_payload_op <= system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_op;
    io_harts_1_dmToHart_regNext_payload_address <= system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_address;
    io_harts_1_dmToHart_regNext_payload_data <= system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_data;
    io_harts_1_dmToHart_regNext_payload_size <= system_riscvJtag_debug_logic_dm_io_harts_1_dmToHart_payload_size;
  end

  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      io_output_cmd_rValid <= 1'b0;
      _zz_when_Stream_l375_3 <= 1'b0;
      io_output_arw_rValidN <= 1'b1;
      io_output_arw_s2mPipe_rValid <= 1'b0;
      io_output_arw_s2mPipe_m2sPipe_rValid <= 1'b0;
      io_output_w_rValidN <= 1'b1;
      io_output_w_s2mPipe_rValid <= 1'b0;
      io_output_w_s2mPipe_m2sPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_cpuAccess_b_rValidN <= 1'b1;
      system_ddr_ddrLogic_cpuAccess_b_s2mPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_cpuAccess_r_rValidN <= 1'b1;
      system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN <= 1'b1;
      system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN <= 1'b1;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN <= 1'b1;
      system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN <= 1'b1;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rValid <= 1'b0;
      io_output_aw_rValidN <= 1'b1;
      io_output_aw_s2mPipe_rValid <= 1'b0;
      io_output_ar_rValidN <= 1'b1;
      io_output_ar_s2mPipe_rValid <= 1'b0;
      io_output_w_rValid <= 1'b0;
      system_ddr_ddrLogic_ddrAAxi4_b_rValidN <= 1'b1;
      system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rValid <= 1'b0;
    end else begin
      if(system_ddr_ddrLogic_cc_fifo_io_output_cmd_ready) begin
        io_output_cmd_rValid <= system_ddr_ddrLogic_cc_fifo_io_output_cmd_valid;
      end
      if(_zz_io_input_rsp_ready_1) begin
        _zz_when_Stream_l375_3 <= system_ddr_ddrLogic_bmbToAxiBridge_io_input_rsp_valid;
      end
      if(system_ddr_ddrLogic_bmbToAxiBridge_io_output_arw_valid) begin
        io_output_arw_rValidN <= 1'b0;
      end
      if(io_output_arw_s2mPipe_ready) begin
        io_output_arw_rValidN <= 1'b1;
      end
      if(io_output_arw_s2mPipe_ready) begin
        io_output_arw_s2mPipe_rValid <= io_output_arw_s2mPipe_valid;
      end
      if(io_output_arw_s2mPipe_m2sPipe_ready) begin
        io_output_arw_s2mPipe_m2sPipe_rValid <= io_output_arw_s2mPipe_m2sPipe_valid;
      end
      if(system_ddr_ddrLogic_bmbToAxiBridge_io_output_w_valid) begin
        io_output_w_rValidN <= 1'b0;
      end
      if(io_output_w_s2mPipe_ready) begin
        io_output_w_rValidN <= 1'b1;
      end
      if(io_output_w_s2mPipe_ready) begin
        io_output_w_s2mPipe_rValid <= io_output_w_s2mPipe_valid;
      end
      if(io_output_w_s2mPipe_m2sPipe_ready) begin
        io_output_w_s2mPipe_m2sPipe_rValid <= io_output_w_s2mPipe_m2sPipe_valid;
      end
      if(system_ddr_ddrLogic_cpuAccess_b_valid) begin
        system_ddr_ddrLogic_cpuAccess_b_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_cpuAccess_b_s2mPipe_ready) begin
        system_ddr_ddrLogic_cpuAccess_b_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_cpuAccess_b_s2mPipe_ready) begin
        system_ddr_ddrLogic_cpuAccess_b_s2mPipe_rValid <= system_ddr_ddrLogic_cpuAccess_b_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_cpuAccess_r_valid) begin
        system_ddr_ddrLogic_cpuAccess_r_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_cpuAccess_r_s2mPipe_ready) begin
        system_ddr_ddrLogic_cpuAccess_r_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_cpuAccess_r_s2mPipe_ready) begin
        system_ddr_ddrLogic_cpuAccess_r_s2mPipe_rValid <= system_ddr_ddrLogic_cpuAccess_r_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_valid) begin
        system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rValid <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_halfPipe_fire) begin
        system_ddr_ddrLogic_userAdapters_0_userAxi4_ar_rValid <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_valid) begin
        system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rValid <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_halfPipe_fire) begin
        system_ddr_ddrLogic_userAdapters_0_userAxi4_aw_rValid <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_0_userAxi4_w_valid) begin
        system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_0_userAxi4_w_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_rValid <= system_ddr_ddrLogic_userAdapters_0_userAxi4_w_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_valid) begin
        system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_rValid <= system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_r_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_valid) begin
        system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rValid <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_halfPipe_fire) begin
        system_ddr_ddrLogic_userAdapters_0_pipelineAxi4_b_rValid <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_valid) begin
        system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rValid <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_halfPipe_fire) begin
        system_ddr_ddrLogic_userAdapters_1_userAxi4_ar_rValid <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_valid) begin
        system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rValid <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_halfPipe_fire) begin
        system_ddr_ddrLogic_userAdapters_1_userAxi4_aw_rValid <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_1_userAxi4_w_valid) begin
        system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_1_userAxi4_w_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_rValid <= system_ddr_ddrLogic_userAdapters_1_userAxi4_w_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_valid) begin
        system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_ready) begin
        system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_rValid <= system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_r_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_valid) begin
        system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rValid <= 1'b1;
      end
      if(system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_halfPipe_fire) begin
        system_ddr_ddrLogic_userAdapters_1_pipelineAxi4_b_rValid <= 1'b0;
      end
      if(system_ddr_ddrLogic_arbiterAxi4Write_io_output_aw_valid) begin
        io_output_aw_rValidN <= 1'b0;
      end
      if(io_output_aw_s2mPipe_ready) begin
        io_output_aw_rValidN <= 1'b1;
      end
      if(io_output_aw_s2mPipe_ready) begin
        io_output_aw_s2mPipe_rValid <= io_output_aw_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_arbiterAxi4Read_io_output_ar_valid) begin
        io_output_ar_rValidN <= 1'b0;
      end
      if(io_output_ar_s2mPipe_ready) begin
        io_output_ar_rValidN <= 1'b1;
      end
      if(io_output_ar_s2mPipe_ready) begin
        io_output_ar_s2mPipe_rValid <= io_output_ar_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_ready) begin
        io_output_w_rValid <= system_ddr_ddrLogic_arbiterAxi4Write_io_output_w_valid;
      end
      if(system_ddr_ddrLogic_ddrAAxi4_b_valid) begin
        system_ddr_ddrLogic_ddrAAxi4_b_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_ready) begin
        system_ddr_ddrLogic_ddrAAxi4_b_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_ready) begin
        system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_rValid <= system_ddr_ddrLogic_ddrAAxi4_b_s2mPipe_valid;
      end
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(io_ddrMasters_1_reset_read_buffer) begin
      io_ddrMasters_1_aw_rValidN <= 1'b1;
      io_ddrMasters_1_aw_s2mPipe_rValid <= 1'b0;
      io_ddrMasters_1_ar_rValid <= 1'b0;
      io_ddrMasters_1_w_rValidN <= 1'b1;
      io_ddrMasters_1_w_s2mPipe_rValid <= 1'b0;
      io_input_r_rValid <= 1'b0;
      io_input_b_rValidN <= 1'b1;
      io_input_b_s2mPipe_rValid <= 1'b0;
    end else begin
      if(io_ddrMasters_1_aw_valid) begin
        io_ddrMasters_1_aw_rValidN <= 1'b0;
      end
      if(io_ddrMasters_1_aw_s2mPipe_ready) begin
        io_ddrMasters_1_aw_rValidN <= 1'b1;
      end
      if(io_ddrMasters_1_aw_s2mPipe_ready) begin
        io_ddrMasters_1_aw_s2mPipe_rValid <= io_ddrMasters_1_aw_s2mPipe_valid;
      end
      if(io_ddrMasters_1_ar_valid) begin
        io_ddrMasters_1_ar_rValid <= 1'b1;
      end
      if(io_ddrMasters_1_ar_halfPipe_fire) begin
        io_ddrMasters_1_ar_rValid <= 1'b0;
      end
      if(io_ddrMasters_1_w_valid) begin
        io_ddrMasters_1_w_rValidN <= 1'b0;
      end
      if(io_ddrMasters_1_w_s2mPipe_ready) begin
        io_ddrMasters_1_w_rValidN <= 1'b1;
      end
      if(io_ddrMasters_1_w_s2mPipe_ready) begin
        io_ddrMasters_1_w_s2mPipe_rValid <= io_ddrMasters_1_w_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_ready) begin
        io_input_r_rValid <= system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_valid) begin
        io_input_b_rValidN <= 1'b0;
      end
      if(io_input_b_s2mPipe_ready) begin
        io_input_b_rValidN <= 1'b1;
      end
      if(io_input_b_s2mPipe_ready) begin
        io_input_b_s2mPipe_rValid <= io_input_b_s2mPipe_valid;
      end
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(io_ddrMasters_1_aw_ready) begin
      io_ddrMasters_1_aw_rData_addr <= io_ddrMasters_1_aw_payload_addr;
      io_ddrMasters_1_aw_rData_id <= io_ddrMasters_1_aw_payload_id;
      io_ddrMasters_1_aw_rData_region <= io_ddrMasters_1_aw_payload_region;
      io_ddrMasters_1_aw_rData_len <= io_ddrMasters_1_aw_payload_len;
      io_ddrMasters_1_aw_rData_size <= io_ddrMasters_1_aw_payload_size;
      io_ddrMasters_1_aw_rData_burst <= io_ddrMasters_1_aw_payload_burst;
      io_ddrMasters_1_aw_rData_lock <= io_ddrMasters_1_aw_payload_lock;
      io_ddrMasters_1_aw_rData_cache <= io_ddrMasters_1_aw_payload_cache;
      io_ddrMasters_1_aw_rData_qos <= io_ddrMasters_1_aw_payload_qos;
      io_ddrMasters_1_aw_rData_prot <= io_ddrMasters_1_aw_payload_prot;
    end
    if(io_ddrMasters_1_aw_s2mPipe_ready) begin
      io_ddrMasters_1_aw_s2mPipe_rData_addr <= io_ddrMasters_1_aw_s2mPipe_payload_addr;
      io_ddrMasters_1_aw_s2mPipe_rData_id <= io_ddrMasters_1_aw_s2mPipe_payload_id;
      io_ddrMasters_1_aw_s2mPipe_rData_region <= io_ddrMasters_1_aw_s2mPipe_payload_region;
      io_ddrMasters_1_aw_s2mPipe_rData_len <= io_ddrMasters_1_aw_s2mPipe_payload_len;
      io_ddrMasters_1_aw_s2mPipe_rData_size <= io_ddrMasters_1_aw_s2mPipe_payload_size;
      io_ddrMasters_1_aw_s2mPipe_rData_burst <= io_ddrMasters_1_aw_s2mPipe_payload_burst;
      io_ddrMasters_1_aw_s2mPipe_rData_lock <= io_ddrMasters_1_aw_s2mPipe_payload_lock;
      io_ddrMasters_1_aw_s2mPipe_rData_cache <= io_ddrMasters_1_aw_s2mPipe_payload_cache;
      io_ddrMasters_1_aw_s2mPipe_rData_qos <= io_ddrMasters_1_aw_s2mPipe_payload_qos;
      io_ddrMasters_1_aw_s2mPipe_rData_prot <= io_ddrMasters_1_aw_s2mPipe_payload_prot;
    end
    if(io_ddrMasters_1_ar_ready) begin
      io_ddrMasters_1_ar_rData_addr <= io_ddrMasters_1_ar_payload_addr;
      io_ddrMasters_1_ar_rData_id <= io_ddrMasters_1_ar_payload_id;
      io_ddrMasters_1_ar_rData_region <= io_ddrMasters_1_ar_payload_region;
      io_ddrMasters_1_ar_rData_len <= io_ddrMasters_1_ar_payload_len;
      io_ddrMasters_1_ar_rData_size <= io_ddrMasters_1_ar_payload_size;
      io_ddrMasters_1_ar_rData_burst <= io_ddrMasters_1_ar_payload_burst;
      io_ddrMasters_1_ar_rData_lock <= io_ddrMasters_1_ar_payload_lock;
      io_ddrMasters_1_ar_rData_cache <= io_ddrMasters_1_ar_payload_cache;
      io_ddrMasters_1_ar_rData_qos <= io_ddrMasters_1_ar_payload_qos;
      io_ddrMasters_1_ar_rData_prot <= io_ddrMasters_1_ar_payload_prot;
    end
    if(io_ddrMasters_1_w_ready) begin
      io_ddrMasters_1_w_rData_data <= io_ddrMasters_1_w_payload_data;
      io_ddrMasters_1_w_rData_strb <= io_ddrMasters_1_w_payload_strb;
      io_ddrMasters_1_w_rData_last <= io_ddrMasters_1_w_payload_last;
    end
    if(io_ddrMasters_1_w_s2mPipe_ready) begin
      io_ddrMasters_1_w_s2mPipe_rData_data <= io_ddrMasters_1_w_s2mPipe_payload_data;
      io_ddrMasters_1_w_s2mPipe_rData_strb <= io_ddrMasters_1_w_s2mPipe_payload_strb;
      io_ddrMasters_1_w_s2mPipe_rData_last <= io_ddrMasters_1_w_s2mPipe_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_ready) begin
      io_input_r_rData_data <= system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_data;
      io_input_r_rData_id <= system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_id;
      io_input_r_rData_resp <= system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_resp;
      io_input_r_rData_last <= system_ddr_ddrLogic_userAdapters_0_bridge_io_input_r_payload_last;
    end
    if(io_input_b_rValidN) begin
      io_input_b_rData_id <= system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_id;
      io_input_b_rData_resp <= system_ddr_ddrLogic_userAdapters_0_bridge_io_input_b_payload_resp;
    end
    if(io_input_b_s2mPipe_ready) begin
      io_input_b_s2mPipe_rData_id <= io_input_b_s2mPipe_payload_id;
      io_input_b_s2mPipe_rData_resp <= io_input_b_s2mPipe_payload_resp;
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(io_ddrMasters_0_reset_read_buffer) begin
      io_ddrMasters_0_aw_rValidN <= 1'b1;
      io_ddrMasters_0_aw_s2mPipe_rValid <= 1'b0;
      io_ddrMasters_0_ar_rValid <= 1'b0;
      io_ddrMasters_0_w_rValidN <= 1'b1;
      io_ddrMasters_0_w_s2mPipe_rValid <= 1'b0;
      io_input_r_rValid_1 <= 1'b0;
      io_input_b_rValidN_1 <= 1'b1;
      io_input_b_s2mPipe_rValid_1 <= 1'b0;
    end else begin
      if(io_ddrMasters_0_aw_valid) begin
        io_ddrMasters_0_aw_rValidN <= 1'b0;
      end
      if(io_ddrMasters_0_aw_s2mPipe_ready) begin
        io_ddrMasters_0_aw_rValidN <= 1'b1;
      end
      if(io_ddrMasters_0_aw_s2mPipe_ready) begin
        io_ddrMasters_0_aw_s2mPipe_rValid <= io_ddrMasters_0_aw_s2mPipe_valid;
      end
      if(io_ddrMasters_0_ar_valid) begin
        io_ddrMasters_0_ar_rValid <= 1'b1;
      end
      if(io_ddrMasters_0_ar_halfPipe_fire) begin
        io_ddrMasters_0_ar_rValid <= 1'b0;
      end
      if(io_ddrMasters_0_w_valid) begin
        io_ddrMasters_0_w_rValidN <= 1'b0;
      end
      if(io_ddrMasters_0_w_s2mPipe_ready) begin
        io_ddrMasters_0_w_rValidN <= 1'b1;
      end
      if(io_ddrMasters_0_w_s2mPipe_ready) begin
        io_ddrMasters_0_w_s2mPipe_rValid <= io_ddrMasters_0_w_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_ready) begin
        io_input_r_rValid_1 <= system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_valid;
      end
      if(system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_valid) begin
        io_input_b_rValidN_1 <= 1'b0;
      end
      if(io_input_b_s2mPipe_ready_1) begin
        io_input_b_rValidN_1 <= 1'b1;
      end
      if(io_input_b_s2mPipe_ready_1) begin
        io_input_b_s2mPipe_rValid_1 <= io_input_b_s2mPipe_valid_1;
      end
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(io_ddrMasters_0_aw_ready) begin
      io_ddrMasters_0_aw_rData_addr <= io_ddrMasters_0_aw_payload_addr;
      io_ddrMasters_0_aw_rData_id <= io_ddrMasters_0_aw_payload_id;
      io_ddrMasters_0_aw_rData_region <= io_ddrMasters_0_aw_payload_region;
      io_ddrMasters_0_aw_rData_len <= io_ddrMasters_0_aw_payload_len;
      io_ddrMasters_0_aw_rData_size <= io_ddrMasters_0_aw_payload_size;
      io_ddrMasters_0_aw_rData_burst <= io_ddrMasters_0_aw_payload_burst;
      io_ddrMasters_0_aw_rData_lock <= io_ddrMasters_0_aw_payload_lock;
      io_ddrMasters_0_aw_rData_cache <= io_ddrMasters_0_aw_payload_cache;
      io_ddrMasters_0_aw_rData_qos <= io_ddrMasters_0_aw_payload_qos;
      io_ddrMasters_0_aw_rData_prot <= io_ddrMasters_0_aw_payload_prot;
    end
    if(io_ddrMasters_0_aw_s2mPipe_ready) begin
      io_ddrMasters_0_aw_s2mPipe_rData_addr <= io_ddrMasters_0_aw_s2mPipe_payload_addr;
      io_ddrMasters_0_aw_s2mPipe_rData_id <= io_ddrMasters_0_aw_s2mPipe_payload_id;
      io_ddrMasters_0_aw_s2mPipe_rData_region <= io_ddrMasters_0_aw_s2mPipe_payload_region;
      io_ddrMasters_0_aw_s2mPipe_rData_len <= io_ddrMasters_0_aw_s2mPipe_payload_len;
      io_ddrMasters_0_aw_s2mPipe_rData_size <= io_ddrMasters_0_aw_s2mPipe_payload_size;
      io_ddrMasters_0_aw_s2mPipe_rData_burst <= io_ddrMasters_0_aw_s2mPipe_payload_burst;
      io_ddrMasters_0_aw_s2mPipe_rData_lock <= io_ddrMasters_0_aw_s2mPipe_payload_lock;
      io_ddrMasters_0_aw_s2mPipe_rData_cache <= io_ddrMasters_0_aw_s2mPipe_payload_cache;
      io_ddrMasters_0_aw_s2mPipe_rData_qos <= io_ddrMasters_0_aw_s2mPipe_payload_qos;
      io_ddrMasters_0_aw_s2mPipe_rData_prot <= io_ddrMasters_0_aw_s2mPipe_payload_prot;
    end
    if(io_ddrMasters_0_ar_ready) begin
      io_ddrMasters_0_ar_rData_addr <= io_ddrMasters_0_ar_payload_addr;
      io_ddrMasters_0_ar_rData_id <= io_ddrMasters_0_ar_payload_id;
      io_ddrMasters_0_ar_rData_region <= io_ddrMasters_0_ar_payload_region;
      io_ddrMasters_0_ar_rData_len <= io_ddrMasters_0_ar_payload_len;
      io_ddrMasters_0_ar_rData_size <= io_ddrMasters_0_ar_payload_size;
      io_ddrMasters_0_ar_rData_burst <= io_ddrMasters_0_ar_payload_burst;
      io_ddrMasters_0_ar_rData_lock <= io_ddrMasters_0_ar_payload_lock;
      io_ddrMasters_0_ar_rData_cache <= io_ddrMasters_0_ar_payload_cache;
      io_ddrMasters_0_ar_rData_qos <= io_ddrMasters_0_ar_payload_qos;
      io_ddrMasters_0_ar_rData_prot <= io_ddrMasters_0_ar_payload_prot;
    end
    if(io_ddrMasters_0_w_ready) begin
      io_ddrMasters_0_w_rData_data <= io_ddrMasters_0_w_payload_data;
      io_ddrMasters_0_w_rData_strb <= io_ddrMasters_0_w_payload_strb;
      io_ddrMasters_0_w_rData_last <= io_ddrMasters_0_w_payload_last;
    end
    if(io_ddrMasters_0_w_s2mPipe_ready) begin
      io_ddrMasters_0_w_s2mPipe_rData_data <= io_ddrMasters_0_w_s2mPipe_payload_data;
      io_ddrMasters_0_w_s2mPipe_rData_strb <= io_ddrMasters_0_w_s2mPipe_payload_strb;
      io_ddrMasters_0_w_s2mPipe_rData_last <= io_ddrMasters_0_w_s2mPipe_payload_last;
    end
    if(system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_ready) begin
      io_input_r_rData_data_1 <= system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_data;
      io_input_r_rData_id_1 <= system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_id;
      io_input_r_rData_resp_1 <= system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_resp;
      io_input_r_rData_last_1 <= system_ddr_ddrLogic_userAdapters_1_bridge_io_input_r_payload_last;
    end
    if(io_input_b_rValidN_1) begin
      io_input_b_rData_id_1 <= system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_id;
      io_input_b_rData_resp_1 <= system_ddr_ddrLogic_userAdapters_1_bridge_io_input_b_payload_resp;
    end
    if(io_input_b_s2mPipe_ready_1) begin
      io_input_b_s2mPipe_rData_id_1 <= io_input_b_s2mPipe_payload_id_1;
      io_input_b_s2mPipe_rData_resp_1 <= io_input_b_s2mPipe_payload_resp_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(when_TrionDdrGenerator_l257) begin
      if(ddrCd_logic_outputReset) begin
        system_ddr_ddrLogic_ddrAReset_counter <= (system_ddr_ddrLogic_ddrAReset_counter + 5'h01);
      end
    end
    system_ddr_ddrLogic_ddrAReset_reset <= system_ddr_ddrLogic_ddrAReset_resetUnbuffered;
  end

  always @(posedge io_memoryClk or posedge system_ddr_ddrLogic_ddrAReset_reset) begin
    if(system_ddr_ddrLogic_ddrAReset_reset) begin
      io_pop_rValidN_2 <= 1'b1;
      io_pop_s2mPipe_rValid_2 <= 1'b0;
      system_ddr_ddrLogic_ddrAToAxi4_ddrA_wCounter <= 8'h0;
      ddrCd_logic_outputReset_regNext <= 1'b0;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN <= 1'b1;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rValid <= 1'b0;
      system_ddr_ddrLogic_ddrAAxi4_ar_rValidN <= 1'b1;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rValid <= 1'b0;
      io_ddrA_r_rValid <= 1'b0;
      io_ddrA_b_rValidN <= 1'b1;
      io_ddrA_b_s2mPipe_rValid <= 1'b0;
      ddrCd_logic_outputReset_regNext_1 <= 1'b0;
    end else begin
      if(system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_valid) begin
        io_pop_rValidN_2 <= 1'b0;
      end
      if(io_pop_s2mPipe_ready_2) begin
        io_pop_rValidN_2 <= 1'b1;
      end
      if(io_pop_s2mPipe_ready_2) begin
        io_pop_s2mPipe_rValid_2 <= io_pop_s2mPipe_valid_2;
      end
      if(system_ddr_ddrLogic_ddrAAxi4_w_fire) begin
        system_ddr_ddrLogic_ddrAToAxi4_ddrA_wCounter <= (system_ddr_ddrLogic_ddrAToAxi4_ddrA_wCounter + 8'h01);
        if(system_ddr_ddrLogic_ddrAAxi4_w_payload_last) begin
          system_ddr_ddrLogic_ddrAToAxi4_ddrA_wCounter <= 8'h0;
        end
      end
      ddrCd_logic_outputReset_regNext <= ddrCd_logic_outputReset;
      if(system_ddr_ddrLogic_ddrAToAxi4_ioAw_valid) begin
        system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_ready) begin
        system_ddr_ddrLogic_ddrAToAxi4_ioAw_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_ready) begin
        system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rValid <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_valid;
      end
      if(system_ddr_ddrLogic_ddrAAxi4_ar_valid) begin
        system_ddr_ddrLogic_ddrAAxi4_ar_rValidN <= 1'b0;
      end
      if(system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_ready) begin
        system_ddr_ddrLogic_ddrAAxi4_ar_rValidN <= 1'b1;
      end
      if(system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_ready) begin
        system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rValid <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_valid;
      end
      if(io_ddrA_r_ready) begin
        io_ddrA_r_rValid <= io_ddrA_r_valid;
      end
      if(io_ddrA_b_valid) begin
        io_ddrA_b_rValidN <= 1'b0;
      end
      if(io_ddrA_b_s2mPipe_ready) begin
        io_ddrA_b_rValidN <= 1'b1;
      end
      if(io_ddrA_b_s2mPipe_ready) begin
        io_ddrA_b_s2mPipe_rValid <= io_ddrA_b_s2mPipe_valid;
      end
      ddrCd_logic_outputReset_regNext_1 <= ddrCd_logic_outputReset;
    end
  end

  always @(posedge io_memoryClk) begin
    if(io_pop_rValidN_2) begin
      io_pop_rData_len <= system_ddr_ddrLogic_ddrAToAxi4_patchAw_translated_fifo_io_pop_payload_len;
    end
    if(io_pop_s2mPipe_ready_2) begin
      io_pop_s2mPipe_rData_len <= io_pop_s2mPipe_payload_len;
    end
    if(system_ddr_ddrLogic_ddrAToAxi4_ioAw_ready) begin
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_addr <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_addr;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_id <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_id;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_region <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_region;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_len <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_len;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_size <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_size;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_burst <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_burst;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_lock <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_lock;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_cache <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_cache;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_qos <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_qos;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_rData_prot <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_payload_prot;
    end
    if(system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_ready) begin
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_addr <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_addr;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_id <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_id;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_region <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_region;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_len <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_len;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_size <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_size;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_burst <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_burst;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_lock <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_lock;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_cache <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_cache;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_qos <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_qos;
      system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_rData_prot <= system_ddr_ddrLogic_ddrAToAxi4_ioAw_s2mPipe_payload_prot;
    end
    if(system_ddr_ddrLogic_ddrAAxi4_ar_ready) begin
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_addr <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_addr;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_id <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_id;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_region <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_region;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_len <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_len;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_size <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_size;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_burst <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_burst;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_lock <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_lock;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_cache <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_cache;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_qos <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_qos;
      system_ddr_ddrLogic_ddrAAxi4_ar_rData_prot <= system_ddr_ddrLogic_ddrAAxi4_ar_payload_prot;
    end
    if(system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_ready) begin
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_addr <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_addr;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_id <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_id;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_region <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_region;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_len <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_len;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_size <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_size;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_burst <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_burst;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_lock <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_lock;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_cache <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_cache;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_qos <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_qos;
      system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_rData_prot <= system_ddr_ddrLogic_ddrAAxi4_ar_s2mPipe_payload_prot;
    end
    if(io_ddrA_r_ready) begin
      io_ddrA_r_rData_data <= io_ddrA_r_payload_data;
      io_ddrA_r_rData_id <= io_ddrA_r_payload_id;
      io_ddrA_r_rData_resp <= io_ddrA_r_payload_resp;
      io_ddrA_r_rData_last <= io_ddrA_r_payload_last;
    end
    if(io_ddrA_b_ready) begin
      io_ddrA_b_rData_id <= io_ddrA_b_payload_id;
      io_ddrA_b_rData_resp <= io_ddrA_b_payload_resp;
    end
    if(io_ddrA_b_s2mPipe_ready) begin
      io_ddrA_b_s2mPipe_rData_id <= io_ddrA_b_s2mPipe_payload_id;
      io_ddrA_b_s2mPipe_rData_resp <= io_ddrA_b_s2mPipe_payload_resp;
    end
  end


endmodule

//BufferCC_73 replaced by BufferCC

//BufferCC_72 replaced by BufferCC

//BufferCC_71 replaced by BufferCC

//BufferCC_70 replaced by BufferCC

//BufferCC_69 replaced by BufferCC

//BufferCC_68 replaced by BufferCC

//StreamCCByToggle_3 replaced by StreamCCByToggle_2

module StreamCCByToggle_2 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [63:0]   io_input_payload,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [63:0]   io_output_payload,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset,
  input  wire          io_systemClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1
);

  wire                outHitSignal_buffercc_io_dataOut;
  wire                pushArea_target_buffercc_io_dataOut;
  wire                outHitSignal;
  wire                pushArea_hit;
  wire                pushArea_accept;
  reg                 pushArea_target;
  reg        [63:0]   pushArea_data;
  wire                io_input_fire;
  wire                popArea_stream_valid;
  reg                 popArea_stream_ready;
  wire       [63:0]   popArea_stream_payload;
  wire                popArea_target;
  wire                popArea_stream_fire;
  reg                 popArea_hit;
  wire                popArea_stream_m2sPipe_valid;
  wire                popArea_stream_m2sPipe_ready;
  wire       [63:0]   popArea_stream_m2sPipe_payload;
  reg                 popArea_stream_rValid;
  (* async_reg = "true" *) reg        [63:0]   popArea_stream_rData;
  wire                when_Stream_l375;

  (* keep_hierarchy = "TRUE" *) BufferCC_45 outHitSignal_buffercc (
    .io_dataIn                      (outHitSignal                    ), //i
    .io_dataOut                     (outHitSignal_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset  )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_44 pushArea_target_buffercc (
    .io_dataIn                                                                           (pushArea_target                                                                    ), //i
    .io_dataOut                                                                          (pushArea_target_buffercc_io_dataOut                                                ), //o
    .io_systemClk                                                                        (io_systemClk                                                                       ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //i
  );
  assign pushArea_hit = outHitSignal_buffercc_io_dataOut;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign pushArea_accept = io_input_fire;
  assign io_input_ready = (pushArea_hit == pushArea_target);
  assign popArea_target = pushArea_target_buffercc_io_dataOut;
  assign popArea_stream_fire = (popArea_stream_valid && popArea_stream_ready);
  assign outHitSignal = popArea_hit;
  assign popArea_stream_valid = (popArea_target != popArea_hit);
  assign popArea_stream_payload = pushArea_data;
  always @(*) begin
    popArea_stream_ready = popArea_stream_m2sPipe_ready;
    if(when_Stream_l375) begin
      popArea_stream_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popArea_stream_m2sPipe_valid);
  assign popArea_stream_m2sPipe_valid = popArea_stream_rValid;
  assign popArea_stream_m2sPipe_payload = popArea_stream_rData;
  assign io_output_valid = popArea_stream_m2sPipe_valid;
  assign popArea_stream_m2sPipe_ready = io_output_ready;
  assign io_output_payload = popArea_stream_m2sPipe_payload;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      pushArea_target <= 1'b0;
    end else begin
      if(pushArea_accept) begin
        pushArea_target <= (! pushArea_target);
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(pushArea_accept) begin
      pushArea_data <= io_input_payload;
    end
  end

  always @(posedge io_systemClk) begin
    if(system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1) begin
      popArea_hit <= 1'b0;
      popArea_stream_rValid <= 1'b0;
    end else begin
      if(popArea_stream_fire) begin
        popArea_hit <= popArea_target;
      end
      if(popArea_stream_ready) begin
        popArea_stream_rValid <= popArea_stream_valid;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(popArea_stream_fire) begin
      popArea_stream_rData <= popArea_stream_payload;
    end
  end


endmodule

//BmbToApb3Bridge_4 replaced by BmbToApb3Bridge

//BmbToApb3Bridge_3 replaced by BmbToApb3Bridge

//BmbToApb3Bridge_2 replaced by BmbToApb3Bridge

//BmbToApb3Bridge_1 replaced by BmbToApb3Bridge

module BmbToApb3Bridge (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [15:0]   io_input_cmd_payload_fragment_address,
  input  wire [1:0]    io_input_cmd_payload_fragment_length,
  input  wire [31:0]   io_input_cmd_payload_fragment_data,
  input  wire [48:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [31:0]   io_input_rsp_payload_fragment_data,
  output wire [48:0]   io_input_rsp_payload_fragment_context,
  output wire [15:0]   io_output_PADDR,
  output wire [0:0]    io_output_PSEL,
  output wire          io_output_PENABLE,
  input  wire          io_output_PREADY,
  output wire          io_output_PWRITE,
  output wire [31:0]   io_output_PWDATA,
  input  wire [31:0]   io_output_PRDATA,
  input  wire          io_output_PSLVERROR,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire                bmbBuffer_cmd_valid;
  reg                 bmbBuffer_cmd_ready;
  wire                bmbBuffer_cmd_payload_last;
  wire       [0:0]    bmbBuffer_cmd_payload_fragment_opcode;
  wire       [15:0]   bmbBuffer_cmd_payload_fragment_address;
  wire       [1:0]    bmbBuffer_cmd_payload_fragment_length;
  wire       [31:0]   bmbBuffer_cmd_payload_fragment_data;
  wire       [48:0]   bmbBuffer_cmd_payload_fragment_context;
  reg                 bmbBuffer_rsp_valid;
  reg                 bmbBuffer_rsp_ready;
  wire                bmbBuffer_rsp_payload_last;
  reg        [0:0]    bmbBuffer_rsp_payload_fragment_opcode;
  wire       [31:0]   bmbBuffer_rsp_payload_fragment_data;
  wire       [48:0]   bmbBuffer_rsp_payload_fragment_context;
  wire                io_input_rsp_isStall;
  wire                _zz_io_input_cmd_ready;
  wire                bmbBuffer_rsp_m2sPipe_valid;
  wire                bmbBuffer_rsp_m2sPipe_ready;
  wire                bmbBuffer_rsp_m2sPipe_payload_last;
  wire       [0:0]    bmbBuffer_rsp_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   bmbBuffer_rsp_m2sPipe_payload_fragment_data;
  wire       [48:0]   bmbBuffer_rsp_m2sPipe_payload_fragment_context;
  reg                 bmbBuffer_rsp_rValid;
  reg                 bmbBuffer_rsp_rData_last;
  reg        [0:0]    bmbBuffer_rsp_rData_fragment_opcode;
  reg        [31:0]   bmbBuffer_rsp_rData_fragment_data;
  reg        [48:0]   bmbBuffer_rsp_rData_fragment_context;
  wire                when_Stream_l375;
  reg                 state;
  wire                when_BmbToApb3Bridge_l46;

  assign io_input_rsp_isStall = (io_input_rsp_valid && (! io_input_rsp_ready));
  assign _zz_io_input_cmd_ready = (! io_input_rsp_isStall);
  assign io_input_cmd_ready = (bmbBuffer_cmd_ready && _zz_io_input_cmd_ready);
  assign bmbBuffer_cmd_valid = (io_input_cmd_valid && _zz_io_input_cmd_ready);
  assign bmbBuffer_cmd_payload_last = io_input_cmd_payload_last;
  assign bmbBuffer_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign bmbBuffer_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign bmbBuffer_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign bmbBuffer_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign bmbBuffer_cmd_payload_fragment_context = io_input_cmd_payload_fragment_context;
  always @(*) begin
    bmbBuffer_rsp_ready = bmbBuffer_rsp_m2sPipe_ready;
    if(when_Stream_l375) begin
      bmbBuffer_rsp_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! bmbBuffer_rsp_m2sPipe_valid);
  assign bmbBuffer_rsp_m2sPipe_valid = bmbBuffer_rsp_rValid;
  assign bmbBuffer_rsp_m2sPipe_payload_last = bmbBuffer_rsp_rData_last;
  assign bmbBuffer_rsp_m2sPipe_payload_fragment_opcode = bmbBuffer_rsp_rData_fragment_opcode;
  assign bmbBuffer_rsp_m2sPipe_payload_fragment_data = bmbBuffer_rsp_rData_fragment_data;
  assign bmbBuffer_rsp_m2sPipe_payload_fragment_context = bmbBuffer_rsp_rData_fragment_context;
  assign io_input_rsp_valid = bmbBuffer_rsp_m2sPipe_valid;
  assign bmbBuffer_rsp_m2sPipe_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = bmbBuffer_rsp_m2sPipe_payload_last;
  assign io_input_rsp_payload_fragment_opcode = bmbBuffer_rsp_m2sPipe_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = bmbBuffer_rsp_m2sPipe_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = bmbBuffer_rsp_m2sPipe_payload_fragment_context;
  always @(*) begin
    bmbBuffer_cmd_ready = 1'b0;
    if(!when_BmbToApb3Bridge_l46) begin
      if(io_output_PREADY) begin
        bmbBuffer_cmd_ready = 1'b1;
      end
    end
  end

  assign io_output_PSEL[0] = bmbBuffer_cmd_valid;
  assign io_output_PENABLE = state;
  assign io_output_PWRITE = (bmbBuffer_cmd_payload_fragment_opcode == 1'b1);
  assign io_output_PADDR = bmbBuffer_cmd_payload_fragment_address;
  assign io_output_PWDATA = bmbBuffer_cmd_payload_fragment_data;
  always @(*) begin
    bmbBuffer_rsp_valid = 1'b0;
    if(!when_BmbToApb3Bridge_l46) begin
      if(io_output_PREADY) begin
        bmbBuffer_rsp_valid = 1'b1;
      end
    end
  end

  assign bmbBuffer_rsp_payload_fragment_data = io_output_PRDATA;
  assign when_BmbToApb3Bridge_l46 = (! state);
  assign bmbBuffer_rsp_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign bmbBuffer_rsp_payload_last = 1'b1;
  always @(*) begin
    bmbBuffer_rsp_payload_fragment_opcode = 1'b0;
    if(io_output_PSLVERROR) begin
      bmbBuffer_rsp_payload_fragment_opcode = 1'b1;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      bmbBuffer_rsp_rValid <= 1'b0;
      state <= 1'b0;
    end else begin
      if(bmbBuffer_rsp_ready) begin
        bmbBuffer_rsp_rValid <= bmbBuffer_rsp_valid;
      end
      if(when_BmbToApb3Bridge_l46) begin
        state <= bmbBuffer_cmd_valid;
      end else begin
        if(io_output_PREADY) begin
          state <= 1'b0;
        end
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(bmbBuffer_rsp_ready) begin
      bmbBuffer_rsp_rData_last <= bmbBuffer_rsp_payload_last;
      bmbBuffer_rsp_rData_fragment_opcode <= bmbBuffer_rsp_payload_fragment_opcode;
      bmbBuffer_rsp_rData_fragment_data <= bmbBuffer_rsp_payload_fragment_data;
      bmbBuffer_rsp_rData_fragment_context <= bmbBuffer_rsp_payload_fragment_context;
    end
  end


endmodule

module BmbWatchdog (
  input  wire          io_bus_cmd_valid,
  output wire          io_bus_cmd_ready,
  input  wire          io_bus_cmd_payload_last,
  input  wire [0:0]    io_bus_cmd_payload_fragment_opcode,
  input  wire [7:0]    io_bus_cmd_payload_fragment_address,
  input  wire [1:0]    io_bus_cmd_payload_fragment_length,
  input  wire [31:0]   io_bus_cmd_payload_fragment_data,
  input  wire [48:0]   io_bus_cmd_payload_fragment_context,
  output wire          io_bus_rsp_valid,
  input  wire          io_bus_rsp_ready,
  output wire          io_bus_rsp_payload_last,
  output wire [0:0]    io_bus_rsp_payload_fragment_opcode,
  output wire [31:0]   io_bus_rsp_payload_fragment_data,
  output wire [48:0]   io_bus_rsp_payload_fragment_context,
  output wire [1:0]    io_panics,
  input  wire          io_heartBeat,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire                wd_prescaler_io_clear;
  wire                wd_prescaler_io_overflow;
  wire                wd_counters_0_timer_io_full;
  wire       [15:0]   wd_counters_0_timer_io_value;
  wire                wd_counters_1_timer_io_full;
  wire       [15:0]   wd_counters_1_timer_io_value;
  reg        [1:0]    wd_api_enables;
  reg                 wd_api_heartbeat;
  reg        [1:0]    wd_api_panics;
  wire                wd_counters_0_clear;
  reg                 wd_counters_0_full;
  wire                wd_counters_1_clear;
  reg                 wd_counters_1_full;
  wire                busCtrl_readErrorFlag;
  wire                busCtrl_writeErrorFlag;
  wire                busCtrl_readHaltTrigger;
  wire                busCtrl_writeHaltTrigger;
  wire                busCtrl_rsp_valid;
  wire                busCtrl_rsp_ready;
  wire                busCtrl_rsp_payload_last;
  reg        [0:0]    busCtrl_rsp_payload_fragment_opcode;
  reg        [31:0]   busCtrl_rsp_payload_fragment_data;
  wire       [48:0]   busCtrl_rsp_payload_fragment_context;
  wire                _zz_busCtrl_rsp_ready;
  reg                 _zz_busCtrl_rsp_ready_1;
  wire                _zz_io_bus_rsp_valid;
  reg                 _zz_io_bus_rsp_valid_1;
  reg                 _zz_io_bus_rsp_payload_last;
  reg        [0:0]    _zz_io_bus_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_bus_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_bus_rsp_payload_fragment_context;
  wire                when_Stream_l375;
  wire                busCtrl_askWrite;
  wire                busCtrl_askRead;
  wire                io_bus_cmd_fire;
  wire                busCtrl_doWrite;
  wire                busCtrl_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  reg                 _zz_wd_api_heartbeat;
  wire       [1:0]    _zz_when_BusSlaveFactory_l379;
  reg                 when_BusSlaveFactory_l377;
  wire                when_BusSlaveFactory_l379;
  wire                when_BusSlaveFactory_l379_1;
  wire                when_Watchdog_l48;
  reg        [23:0]   _zz_io_limit;
  wire                when_Watchdog_l48_1;
  reg        [15:0]   _zz_io_limit_1;
  wire                when_Watchdog_l48_2;
  reg        [15:0]   _zz_io_limit_2;

  Prescaler_2 wd_prescaler (
    .io_clear                       (wd_prescaler_io_clear         ), //i
    .io_limit                       (_zz_io_limit[23:0]            ), //i
    .io_overflow                    (wd_prescaler_io_overflow      ), //o
    .io_peripheralClk               (io_peripheralClk              ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset)  //i
  );
  Timer_2 wd_counters_0_timer (
    .io_tick                        (wd_prescaler_io_overflow          ), //i
    .io_clear                       (wd_counters_0_clear               ), //i
    .io_limit                       (_zz_io_limit_1[15:0]              ), //i
    .io_full                        (wd_counters_0_timer_io_full       ), //o
    .io_value                       (wd_counters_0_timer_io_value[15:0]), //o
    .io_peripheralClk               (io_peripheralClk                  ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset    )  //i
  );
  Timer_2 wd_counters_1_timer (
    .io_tick                        (wd_prescaler_io_overflow          ), //i
    .io_clear                       (wd_counters_1_clear               ), //i
    .io_limit                       (_zz_io_limit_2[15:0]              ), //i
    .io_full                        (wd_counters_1_timer_io_full       ), //o
    .io_value                       (wd_counters_1_timer_io_value[15:0]), //o
    .io_peripheralClk               (io_peripheralClk                  ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset    )  //i
  );
  assign wd_prescaler_io_clear = (wd_api_heartbeat || (wd_api_enables == 2'b00));
  assign wd_counters_0_clear = ((! wd_api_enables[0]) || wd_api_heartbeat);
  always @(*) begin
    wd_api_panics[0] = wd_counters_0_full;
    wd_api_panics[1] = wd_counters_1_full;
  end

  assign wd_counters_1_clear = ((! wd_api_enables[1]) || wd_api_heartbeat);
  assign busCtrl_readErrorFlag = 1'b0;
  assign busCtrl_writeErrorFlag = 1'b0;
  assign busCtrl_readHaltTrigger = 1'b0;
  assign busCtrl_writeHaltTrigger = 1'b0;
  assign _zz_busCtrl_rsp_ready = (! (busCtrl_readHaltTrigger || busCtrl_writeHaltTrigger));
  assign busCtrl_rsp_ready = (_zz_busCtrl_rsp_ready_1 && _zz_busCtrl_rsp_ready);
  always @(*) begin
    _zz_busCtrl_rsp_ready_1 = io_bus_rsp_ready;
    if(when_Stream_l375) begin
      _zz_busCtrl_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375 = (! _zz_io_bus_rsp_valid);
  assign _zz_io_bus_rsp_valid = _zz_io_bus_rsp_valid_1;
  assign io_bus_rsp_valid = _zz_io_bus_rsp_valid;
  assign io_bus_rsp_payload_last = _zz_io_bus_rsp_payload_last;
  assign io_bus_rsp_payload_fragment_opcode = _zz_io_bus_rsp_payload_fragment_opcode;
  assign io_bus_rsp_payload_fragment_data = _zz_io_bus_rsp_payload_fragment_data;
  assign io_bus_rsp_payload_fragment_context = _zz_io_bus_rsp_payload_fragment_context;
  assign busCtrl_askWrite = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_askRead = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign io_bus_cmd_fire = (io_bus_cmd_valid && io_bus_cmd_ready);
  assign busCtrl_doWrite = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_doRead = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign busCtrl_rsp_valid = io_bus_cmd_valid;
  assign io_bus_cmd_ready = busCtrl_rsp_ready;
  assign busCtrl_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (busCtrl_doWrite && busCtrl_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      busCtrl_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        busCtrl_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        busCtrl_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (busCtrl_doRead && busCtrl_readErrorFlag);
  always @(*) begin
    busCtrl_rsp_payload_fragment_data = 32'h0;
    case(io_bus_cmd_payload_fragment_address)
      8'hc0 : begin
        busCtrl_rsp_payload_fragment_data[15 : 0] = wd_counters_0_timer_io_value;
      end
      8'hc4 : begin
        busCtrl_rsp_payload_fragment_data[15 : 0] = wd_counters_1_timer_io_value;
      end
      default : begin
      end
    endcase
  end

  assign busCtrl_rsp_payload_fragment_context = io_bus_cmd_payload_fragment_context;
  always @(*) begin
    _zz_wd_api_heartbeat = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      8'h0 : begin
        if(busCtrl_doWrite) begin
          _zz_wd_api_heartbeat = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    wd_api_heartbeat = (_zz_wd_api_heartbeat && (io_bus_cmd_payload_fragment_data[31 : 0] == 32'had68e70d));
    if(io_heartBeat) begin
      wd_api_heartbeat = 1'b1;
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377 = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      8'h04 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l377 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379 = _zz_when_BusSlaveFactory_l379[0];
  assign when_BusSlaveFactory_l379_1 = _zz_when_BusSlaveFactory_l379[1];
  assign when_Watchdog_l48 = (wd_api_enables == 2'b00);
  assign when_Watchdog_l48_1 = (! wd_api_enables[0]);
  assign when_Watchdog_l48_2 = (! wd_api_enables[1]);
  assign io_panics = wd_api_panics;
  assign _zz_when_BusSlaveFactory_l379 = io_bus_cmd_payload_fragment_data[1 : 0];
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      wd_counters_0_full <= 1'b0;
      wd_counters_1_full <= 1'b0;
      _zz_io_bus_rsp_valid_1 <= 1'b0;
      wd_api_enables <= 2'b00;
      _zz_io_limit <= 24'h0;
      _zz_io_limit_1 <= 16'h0;
      _zz_io_limit_2 <= 16'h0;
    end else begin
      if(wd_counters_0_timer_io_full) begin
        wd_counters_0_full <= 1'b1;
      end
      if(wd_counters_0_clear) begin
        wd_counters_0_full <= 1'b0;
      end
      if(wd_counters_1_timer_io_full) begin
        wd_counters_1_full <= 1'b1;
      end
      if(wd_counters_1_clear) begin
        wd_counters_1_full <= 1'b0;
      end
      if(_zz_busCtrl_rsp_ready_1) begin
        _zz_io_bus_rsp_valid_1 <= (busCtrl_rsp_valid && _zz_busCtrl_rsp_ready);
      end
      if(when_BusSlaveFactory_l377) begin
        if(when_BusSlaveFactory_l379) begin
          wd_api_enables[0 : 0] <= 1'b1;
        end
        if(when_BusSlaveFactory_l379_1) begin
          wd_api_enables[1 : 1] <= 1'b1;
        end
      end
      case(io_bus_cmd_payload_fragment_address)
        8'h40 : begin
          if(busCtrl_doWrite) begin
            if(when_Watchdog_l48) begin
              _zz_io_limit <= io_bus_cmd_payload_fragment_data[23 : 0];
            end
          end
        end
        8'h80 : begin
          if(busCtrl_doWrite) begin
            if(when_Watchdog_l48_1) begin
              _zz_io_limit_1 <= io_bus_cmd_payload_fragment_data[15 : 0];
            end
          end
        end
        8'h84 : begin
          if(busCtrl_doWrite) begin
            if(when_Watchdog_l48_2) begin
              _zz_io_limit_2 <= io_bus_cmd_payload_fragment_data[15 : 0];
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_peripheralClk) begin
    if(_zz_busCtrl_rsp_ready_1) begin
      _zz_io_bus_rsp_payload_last <= busCtrl_rsp_payload_last;
      _zz_io_bus_rsp_payload_fragment_opcode <= busCtrl_rsp_payload_fragment_opcode;
      _zz_io_bus_rsp_payload_fragment_data <= busCtrl_rsp_payload_fragment_data;
      _zz_io_bus_rsp_payload_fragment_context <= busCtrl_rsp_payload_fragment_context;
    end
  end


endmodule

module BmbGpio2 (
  input  wire [3:0]    io_gpio_read,
  output reg  [3:0]    io_gpio_write,
  output reg  [3:0]    io_gpio_writeEnable,
  input  wire          io_bus_cmd_valid,
  output wire          io_bus_cmd_ready,
  input  wire          io_bus_cmd_payload_last,
  input  wire [0:0]    io_bus_cmd_payload_fragment_opcode,
  input  wire [7:0]    io_bus_cmd_payload_fragment_address,
  input  wire [1:0]    io_bus_cmd_payload_fragment_length,
  input  wire [31:0]   io_bus_cmd_payload_fragment_data,
  input  wire [48:0]   io_bus_cmd_payload_fragment_context,
  output wire          io_bus_rsp_valid,
  input  wire          io_bus_rsp_ready,
  output wire          io_bus_rsp_payload_last,
  output wire [0:0]    io_bus_rsp_payload_fragment_opcode,
  output wire [31:0]   io_bus_rsp_payload_fragment_data,
  output wire [48:0]   io_bus_rsp_payload_fragment_context,
  output reg  [3:0]    io_interrupt,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire                mapper_readErrorFlag;
  wire                mapper_writeErrorFlag;
  wire                mapper_readHaltTrigger;
  wire                mapper_writeHaltTrigger;
  wire                mapper_rsp_valid;
  wire                mapper_rsp_ready;
  wire                mapper_rsp_payload_last;
  reg        [0:0]    mapper_rsp_payload_fragment_opcode;
  reg        [31:0]   mapper_rsp_payload_fragment_data;
  wire       [48:0]   mapper_rsp_payload_fragment_context;
  wire                _zz_mapper_rsp_ready;
  reg                 _zz_mapper_rsp_ready_1;
  wire                _zz_io_bus_rsp_valid;
  reg                 _zz_io_bus_rsp_valid_1;
  reg                 _zz_io_bus_rsp_payload_last;
  reg        [0:0]    _zz_io_bus_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_bus_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_bus_rsp_payload_fragment_context;
  wire                when_Stream_l375;
  wire                mapper_askWrite;
  wire                mapper_askRead;
  wire                io_bus_cmd_fire;
  wire                mapper_doWrite;
  wire                mapper_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  reg        [3:0]    io_gpio_read_delay_1;
  reg        [3:0]    syncronized;
  reg        [3:0]    last;
  reg                 _zz_io_gpio_write;
  reg                 _zz_io_gpio_writeEnable;
  reg                 _zz_io_gpio_write_1;
  reg                 _zz_io_gpio_writeEnable_1;
  reg                 _zz_io_gpio_write_2;
  reg                 _zz_io_gpio_writeEnable_2;
  reg                 _zz_io_gpio_write_3;
  reg                 _zz_io_gpio_writeEnable_3;
  reg        [3:0]    interrupt_enable_high;
  reg        [3:0]    interrupt_enable_low;
  reg        [3:0]    interrupt_enable_rise;
  reg        [3:0]    interrupt_enable_fall;
  wire       [3:0]    interrupt_valid;
  reg                 _zz_mapper_rsp_payload_fragment_data;
  reg                 _zz_mapper_rsp_payload_fragment_data_1;
  reg                 _zz_mapper_rsp_payload_fragment_data_2;
  reg                 _zz_mapper_rsp_payload_fragment_data_3;
  reg                 _zz_mapper_rsp_payload_fragment_data_4;
  reg                 _zz_mapper_rsp_payload_fragment_data_5;
  reg                 _zz_mapper_rsp_payload_fragment_data_6;
  reg                 _zz_mapper_rsp_payload_fragment_data_7;

  assign mapper_readErrorFlag = 1'b0;
  assign mapper_writeErrorFlag = 1'b0;
  assign mapper_readHaltTrigger = 1'b0;
  assign mapper_writeHaltTrigger = 1'b0;
  assign _zz_mapper_rsp_ready = (! (mapper_readHaltTrigger || mapper_writeHaltTrigger));
  assign mapper_rsp_ready = (_zz_mapper_rsp_ready_1 && _zz_mapper_rsp_ready);
  always @(*) begin
    _zz_mapper_rsp_ready_1 = io_bus_rsp_ready;
    if(when_Stream_l375) begin
      _zz_mapper_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375 = (! _zz_io_bus_rsp_valid);
  assign _zz_io_bus_rsp_valid = _zz_io_bus_rsp_valid_1;
  assign io_bus_rsp_valid = _zz_io_bus_rsp_valid;
  assign io_bus_rsp_payload_last = _zz_io_bus_rsp_payload_last;
  assign io_bus_rsp_payload_fragment_opcode = _zz_io_bus_rsp_payload_fragment_opcode;
  assign io_bus_rsp_payload_fragment_data = _zz_io_bus_rsp_payload_fragment_data;
  assign io_bus_rsp_payload_fragment_context = _zz_io_bus_rsp_payload_fragment_context;
  assign mapper_askWrite = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign mapper_askRead = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign io_bus_cmd_fire = (io_bus_cmd_valid && io_bus_cmd_ready);
  assign mapper_doWrite = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign mapper_doRead = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign mapper_rsp_valid = io_bus_cmd_valid;
  assign io_bus_cmd_ready = mapper_rsp_ready;
  assign mapper_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (mapper_doWrite && mapper_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      mapper_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        mapper_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        mapper_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (mapper_doRead && mapper_readErrorFlag);
  always @(*) begin
    mapper_rsp_payload_fragment_data = 32'h0;
    case(io_bus_cmd_payload_fragment_address)
      8'h0 : begin
        mapper_rsp_payload_fragment_data[0 : 0] = syncronized[0];
        mapper_rsp_payload_fragment_data[1 : 1] = syncronized[1];
        mapper_rsp_payload_fragment_data[2 : 2] = syncronized[2];
        mapper_rsp_payload_fragment_data[3 : 3] = syncronized[3];
      end
      8'h04 : begin
        mapper_rsp_payload_fragment_data[0 : 0] = _zz_io_gpio_write;
        mapper_rsp_payload_fragment_data[1 : 1] = _zz_io_gpio_write_1;
        mapper_rsp_payload_fragment_data[2 : 2] = _zz_io_gpio_write_2;
        mapper_rsp_payload_fragment_data[3 : 3] = _zz_io_gpio_write_3;
      end
      8'h08 : begin
        mapper_rsp_payload_fragment_data[0 : 0] = _zz_io_gpio_writeEnable;
        mapper_rsp_payload_fragment_data[1 : 1] = _zz_io_gpio_writeEnable_1;
        mapper_rsp_payload_fragment_data[2 : 2] = _zz_io_gpio_writeEnable_2;
        mapper_rsp_payload_fragment_data[3 : 3] = _zz_io_gpio_writeEnable_3;
      end
      8'h20 : begin
        mapper_rsp_payload_fragment_data[0 : 0] = _zz_mapper_rsp_payload_fragment_data;
        mapper_rsp_payload_fragment_data[1 : 1] = _zz_mapper_rsp_payload_fragment_data_4;
      end
      8'h24 : begin
        mapper_rsp_payload_fragment_data[0 : 0] = _zz_mapper_rsp_payload_fragment_data_1;
        mapper_rsp_payload_fragment_data[1 : 1] = _zz_mapper_rsp_payload_fragment_data_5;
      end
      8'h28 : begin
        mapper_rsp_payload_fragment_data[0 : 0] = _zz_mapper_rsp_payload_fragment_data_2;
        mapper_rsp_payload_fragment_data[1 : 1] = _zz_mapper_rsp_payload_fragment_data_6;
      end
      8'h2c : begin
        mapper_rsp_payload_fragment_data[0 : 0] = _zz_mapper_rsp_payload_fragment_data_3;
        mapper_rsp_payload_fragment_data[1 : 1] = _zz_mapper_rsp_payload_fragment_data_7;
      end
      default : begin
      end
    endcase
  end

  assign mapper_rsp_payload_fragment_context = io_bus_cmd_payload_fragment_context;
  always @(*) begin
    io_gpio_write[0] = _zz_io_gpio_write;
    io_gpio_write[1] = _zz_io_gpio_write_1;
    io_gpio_write[2] = _zz_io_gpio_write_2;
    io_gpio_write[3] = _zz_io_gpio_write_3;
  end

  always @(*) begin
    io_gpio_writeEnable[0] = _zz_io_gpio_writeEnable;
    io_gpio_writeEnable[1] = _zz_io_gpio_writeEnable_1;
    io_gpio_writeEnable[2] = _zz_io_gpio_writeEnable_2;
    io_gpio_writeEnable[3] = _zz_io_gpio_writeEnable_3;
  end

  assign interrupt_valid = ((((interrupt_enable_high & syncronized) | (interrupt_enable_low & (~ syncronized))) | (interrupt_enable_rise & (syncronized & (~ last)))) | (interrupt_enable_fall & ((~ syncronized) & last)));
  always @(*) begin
    io_interrupt[0] = interrupt_valid[0];
    io_interrupt[1] = interrupt_valid[1];
    io_interrupt[2] = 1'b0;
    io_interrupt[3] = 1'b0;
  end

  always @(*) begin
    interrupt_enable_rise[0] = _zz_mapper_rsp_payload_fragment_data;
    interrupt_enable_rise[1] = _zz_mapper_rsp_payload_fragment_data_4;
    interrupt_enable_rise[2] = 1'b0;
    interrupt_enable_rise[3] = 1'b0;
  end

  always @(*) begin
    interrupt_enable_fall[0] = _zz_mapper_rsp_payload_fragment_data_1;
    interrupt_enable_fall[1] = _zz_mapper_rsp_payload_fragment_data_5;
    interrupt_enable_fall[2] = 1'b0;
    interrupt_enable_fall[3] = 1'b0;
  end

  always @(*) begin
    interrupt_enable_high[0] = _zz_mapper_rsp_payload_fragment_data_2;
    interrupt_enable_high[1] = _zz_mapper_rsp_payload_fragment_data_6;
    interrupt_enable_high[2] = 1'b0;
    interrupt_enable_high[3] = 1'b0;
  end

  always @(*) begin
    interrupt_enable_low[0] = _zz_mapper_rsp_payload_fragment_data_3;
    interrupt_enable_low[1] = _zz_mapper_rsp_payload_fragment_data_7;
    interrupt_enable_low[2] = 1'b0;
    interrupt_enable_low[3] = 1'b0;
  end

  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      _zz_io_bus_rsp_valid_1 <= 1'b0;
      _zz_io_gpio_writeEnable <= 1'b0;
      _zz_io_gpio_writeEnable_1 <= 1'b0;
      _zz_io_gpio_writeEnable_2 <= 1'b0;
      _zz_io_gpio_writeEnable_3 <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data_1 <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data_2 <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data_3 <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data_4 <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data_5 <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data_6 <= 1'b0;
      _zz_mapper_rsp_payload_fragment_data_7 <= 1'b0;
    end else begin
      if(_zz_mapper_rsp_ready_1) begin
        _zz_io_bus_rsp_valid_1 <= (mapper_rsp_valid && _zz_mapper_rsp_ready);
      end
      case(io_bus_cmd_payload_fragment_address)
        8'h08 : begin
          if(mapper_doWrite) begin
            _zz_io_gpio_writeEnable <= io_bus_cmd_payload_fragment_data[0];
            _zz_io_gpio_writeEnable_1 <= io_bus_cmd_payload_fragment_data[1];
            _zz_io_gpio_writeEnable_2 <= io_bus_cmd_payload_fragment_data[2];
            _zz_io_gpio_writeEnable_3 <= io_bus_cmd_payload_fragment_data[3];
          end
        end
        8'h20 : begin
          if(mapper_doWrite) begin
            _zz_mapper_rsp_payload_fragment_data <= io_bus_cmd_payload_fragment_data[0];
            _zz_mapper_rsp_payload_fragment_data_4 <= io_bus_cmd_payload_fragment_data[1];
          end
        end
        8'h24 : begin
          if(mapper_doWrite) begin
            _zz_mapper_rsp_payload_fragment_data_1 <= io_bus_cmd_payload_fragment_data[0];
            _zz_mapper_rsp_payload_fragment_data_5 <= io_bus_cmd_payload_fragment_data[1];
          end
        end
        8'h28 : begin
          if(mapper_doWrite) begin
            _zz_mapper_rsp_payload_fragment_data_2 <= io_bus_cmd_payload_fragment_data[0];
            _zz_mapper_rsp_payload_fragment_data_6 <= io_bus_cmd_payload_fragment_data[1];
          end
        end
        8'h2c : begin
          if(mapper_doWrite) begin
            _zz_mapper_rsp_payload_fragment_data_3 <= io_bus_cmd_payload_fragment_data[0];
            _zz_mapper_rsp_payload_fragment_data_7 <= io_bus_cmd_payload_fragment_data[1];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_peripheralClk) begin
    if(_zz_mapper_rsp_ready_1) begin
      _zz_io_bus_rsp_payload_last <= mapper_rsp_payload_last;
      _zz_io_bus_rsp_payload_fragment_opcode <= mapper_rsp_payload_fragment_opcode;
      _zz_io_bus_rsp_payload_fragment_data <= mapper_rsp_payload_fragment_data;
      _zz_io_bus_rsp_payload_fragment_context <= mapper_rsp_payload_fragment_context;
    end
    io_gpio_read_delay_1 <= io_gpio_read;
    syncronized <= io_gpio_read_delay_1;
    last <= syncronized;
    case(io_bus_cmd_payload_fragment_address)
      8'h04 : begin
        if(mapper_doWrite) begin
          _zz_io_gpio_write <= io_bus_cmd_payload_fragment_data[0];
          _zz_io_gpio_write_1 <= io_bus_cmd_payload_fragment_data[1];
          _zz_io_gpio_write_2 <= io_bus_cmd_payload_fragment_data[2];
          _zz_io_gpio_write_3 <= io_bus_cmd_payload_fragment_data[3];
        end
      end
      default : begin
      end
    endcase
  end


endmodule

//EfxTimerCtrl_1 replaced by EfxTimerCtrl

module EfxTimerCtrl (
  input  wire          io_ctrl_cmd_valid,
  output wire          io_ctrl_cmd_ready,
  input  wire          io_ctrl_cmd_payload_last,
  input  wire [0:0]    io_ctrl_cmd_payload_fragment_opcode,
  input  wire [7:0]    io_ctrl_cmd_payload_fragment_address,
  input  wire [1:0]    io_ctrl_cmd_payload_fragment_length,
  input  wire [31:0]   io_ctrl_cmd_payload_fragment_data,
  input  wire [48:0]   io_ctrl_cmd_payload_fragment_context,
  output wire          io_ctrl_rsp_valid,
  input  wire          io_ctrl_rsp_ready,
  output wire          io_ctrl_rsp_payload_last,
  output wire [0:0]    io_ctrl_rsp_payload_fragment_opcode,
  output wire [31:0]   io_ctrl_rsp_payload_fragment_data,
  output wire [48:0]   io_ctrl_rsp_payload_fragment_context,
  output wire [0:0]    io_interrupts,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire                timer_4_io_tick;
  wire                timer_4_io_clear;
  wire                prescaler_3_io_overflow;
  wire                timer_4_io_full;
  wire       [11:0]   timer_4_io_value;
  wire                busCtrl_readErrorFlag;
  wire                busCtrl_writeErrorFlag;
  wire                busCtrl_readHaltTrigger;
  wire                busCtrl_writeHaltTrigger;
  wire                busCtrl_rsp_valid;
  wire                busCtrl_rsp_ready;
  wire                busCtrl_rsp_payload_last;
  reg        [0:0]    busCtrl_rsp_payload_fragment_opcode;
  reg        [31:0]   busCtrl_rsp_payload_fragment_data;
  wire       [48:0]   busCtrl_rsp_payload_fragment_context;
  wire                _zz_busCtrl_rsp_ready;
  reg                 _zz_busCtrl_rsp_ready_1;
  wire                _zz_io_ctrl_rsp_valid;
  reg                 _zz_io_ctrl_rsp_valid_1;
  reg                 _zz_io_ctrl_rsp_payload_last;
  reg        [0:0]    _zz_io_ctrl_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_ctrl_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_ctrl_rsp_payload_fragment_context;
  wire                when_Stream_l375;
  wire                busCtrl_askWrite;
  wire                busCtrl_askRead;
  wire                io_ctrl_cmd_fire;
  wire                busCtrl_doWrite;
  wire                busCtrl_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  reg        [7:0]    _zz_io_limit;
  reg                 _zz_io_clear;
  reg        [1:0]    _zz_busCtrl_rsp_payload_fragment_data;
  reg        [0:0]    _zz_busCtrl_rsp_payload_fragment_data_1;
  reg                 _zz_io_clear_1;
  reg        [11:0]   timer_4_io_limit_driver;
  reg                 when_Timer_l40;
  reg                 when_Timer_l44;

  Prescaler prescaler_3 (
    .io_clear                       (_zz_io_clear                  ), //i
    .io_limit                       (_zz_io_limit[7:0]             ), //i
    .io_overflow                    (prescaler_3_io_overflow       ), //o
    .io_peripheralClk               (io_peripheralClk              ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset)  //i
  );
  Timer timer_4 (
    .io_tick                        (timer_4_io_tick               ), //i
    .io_clear                       (timer_4_io_clear              ), //i
    .io_limit                       (timer_4_io_limit_driver[11:0] ), //i
    .io_full                        (timer_4_io_full               ), //o
    .io_value                       (timer_4_io_value[11:0]        ), //o
    .io_peripheralClk               (io_peripheralClk              ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset)  //i
  );
  assign busCtrl_readErrorFlag = 1'b0;
  assign busCtrl_writeErrorFlag = 1'b0;
  assign busCtrl_readHaltTrigger = 1'b0;
  assign busCtrl_writeHaltTrigger = 1'b0;
  assign _zz_busCtrl_rsp_ready = (! (busCtrl_readHaltTrigger || busCtrl_writeHaltTrigger));
  assign busCtrl_rsp_ready = (_zz_busCtrl_rsp_ready_1 && _zz_busCtrl_rsp_ready);
  always @(*) begin
    _zz_busCtrl_rsp_ready_1 = io_ctrl_rsp_ready;
    if(when_Stream_l375) begin
      _zz_busCtrl_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375 = (! _zz_io_ctrl_rsp_valid);
  assign _zz_io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid_1;
  assign io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid;
  assign io_ctrl_rsp_payload_last = _zz_io_ctrl_rsp_payload_last;
  assign io_ctrl_rsp_payload_fragment_opcode = _zz_io_ctrl_rsp_payload_fragment_opcode;
  assign io_ctrl_rsp_payload_fragment_data = _zz_io_ctrl_rsp_payload_fragment_data;
  assign io_ctrl_rsp_payload_fragment_context = _zz_io_ctrl_rsp_payload_fragment_context;
  assign busCtrl_askWrite = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_askRead = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign io_ctrl_cmd_fire = (io_ctrl_cmd_valid && io_ctrl_cmd_ready);
  assign busCtrl_doWrite = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_doRead = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign busCtrl_rsp_valid = io_ctrl_cmd_valid;
  assign io_ctrl_cmd_ready = busCtrl_rsp_ready;
  assign busCtrl_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (busCtrl_doWrite && busCtrl_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      busCtrl_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        busCtrl_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        busCtrl_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (busCtrl_doRead && busCtrl_readErrorFlag);
  always @(*) begin
    busCtrl_rsp_payload_fragment_data = 32'h0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h0 : begin
        busCtrl_rsp_payload_fragment_data[7 : 0] = _zz_io_limit;
      end
      8'h40 : begin
        busCtrl_rsp_payload_fragment_data[1 : 0] = _zz_busCtrl_rsp_payload_fragment_data;
        busCtrl_rsp_payload_fragment_data[16 : 16] = _zz_busCtrl_rsp_payload_fragment_data_1;
      end
      8'h44 : begin
        busCtrl_rsp_payload_fragment_data[11 : 0] = timer_4_io_limit_driver;
      end
      8'h48 : begin
        busCtrl_rsp_payload_fragment_data[11 : 0] = timer_4_io_value;
      end
      default : begin
      end
    endcase
  end

  assign busCtrl_rsp_payload_fragment_context = io_ctrl_cmd_payload_fragment_context;
  always @(*) begin
    _zz_io_clear = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h0 : begin
        if(busCtrl_doWrite) begin
          _zz_io_clear = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_clear_1 = 1'b0;
    if(when_Timer_l40) begin
      _zz_io_clear_1 = 1'b1;
    end
    if(when_Timer_l44) begin
      _zz_io_clear_1 = 1'b1;
    end
  end

  always @(*) begin
    when_Timer_l40 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h44 : begin
        if(busCtrl_doWrite) begin
          when_Timer_l40 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    when_Timer_l44 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h48 : begin
        if(busCtrl_doWrite) begin
          when_Timer_l44 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign timer_4_io_clear = ((|(_zz_busCtrl_rsp_payload_fragment_data_1 & timer_4_io_full)) || _zz_io_clear_1);
  assign timer_4_io_tick = (|(_zz_busCtrl_rsp_payload_fragment_data & {prescaler_3_io_overflow,1'b1}));
  assign io_interrupts[0] = timer_4_io_full;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      _zz_io_ctrl_rsp_valid_1 <= 1'b0;
      _zz_busCtrl_rsp_payload_fragment_data <= 2'b00;
      _zz_busCtrl_rsp_payload_fragment_data_1 <= 1'b0;
    end else begin
      if(_zz_busCtrl_rsp_ready_1) begin
        _zz_io_ctrl_rsp_valid_1 <= (busCtrl_rsp_valid && _zz_busCtrl_rsp_ready);
      end
      case(io_ctrl_cmd_payload_fragment_address)
        8'h40 : begin
          if(busCtrl_doWrite) begin
            _zz_busCtrl_rsp_payload_fragment_data <= io_ctrl_cmd_payload_fragment_data[1 : 0];
            _zz_busCtrl_rsp_payload_fragment_data_1 <= io_ctrl_cmd_payload_fragment_data[16 : 16];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_peripheralClk) begin
    if(_zz_busCtrl_rsp_ready_1) begin
      _zz_io_ctrl_rsp_payload_last <= busCtrl_rsp_payload_last;
      _zz_io_ctrl_rsp_payload_fragment_opcode <= busCtrl_rsp_payload_fragment_opcode;
      _zz_io_ctrl_rsp_payload_fragment_data <= busCtrl_rsp_payload_fragment_data;
      _zz_io_ctrl_rsp_payload_fragment_context <= busCtrl_rsp_payload_fragment_context;
    end
    case(io_ctrl_cmd_payload_fragment_address)
      8'h0 : begin
        if(busCtrl_doWrite) begin
          _zz_io_limit <= io_ctrl_cmd_payload_fragment_data[7 : 0];
        end
      end
      8'h44 : begin
        if(busCtrl_doWrite) begin
          timer_4_io_limit_driver <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      default : begin
      end
    endcase
  end


endmodule

//BmbI2cCtrl_2 replaced by BmbI2cCtrl

//BmbI2cCtrl_1 replaced by BmbI2cCtrl

module BmbI2cCtrl (
  input  wire          io_ctrl_cmd_valid,
  output wire          io_ctrl_cmd_ready,
  input  wire          io_ctrl_cmd_payload_last,
  input  wire [0:0]    io_ctrl_cmd_payload_fragment_opcode,
  input  wire [7:0]    io_ctrl_cmd_payload_fragment_address,
  input  wire [1:0]    io_ctrl_cmd_payload_fragment_length,
  input  wire [31:0]   io_ctrl_cmd_payload_fragment_data,
  input  wire [48:0]   io_ctrl_cmd_payload_fragment_context,
  output wire          io_ctrl_rsp_valid,
  input  wire          io_ctrl_rsp_ready,
  output wire          io_ctrl_rsp_payload_last,
  output wire [0:0]    io_ctrl_rsp_payload_fragment_opcode,
  output wire [31:0]   io_ctrl_rsp_payload_fragment_data,
  output wire [48:0]   io_ctrl_rsp_payload_fragment_context,
  output wire          io_i2c_sda_write,
  input  wire          io_i2c_sda_read,
  output wire          io_i2c_scl_write,
  input  wire          io_i2c_scl_read,
  output wire          io_interrupt,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);
  localparam bridge_masterLogic_fsm_enumDef_BOOT = 4'd0;
  localparam bridge_masterLogic_fsm_enumDef_IDLE = 4'd1;
  localparam bridge_masterLogic_fsm_enumDef_START1 = 4'd2;
  localparam bridge_masterLogic_fsm_enumDef_START2 = 4'd3;
  localparam bridge_masterLogic_fsm_enumDef_START3 = 4'd4;
  localparam bridge_masterLogic_fsm_enumDef_LOW = 4'd5;
  localparam bridge_masterLogic_fsm_enumDef_HIGH = 4'd6;
  localparam bridge_masterLogic_fsm_enumDef_RESTART = 4'd7;
  localparam bridge_masterLogic_fsm_enumDef_STOP1 = 4'd8;
  localparam bridge_masterLogic_fsm_enumDef_STOP2 = 4'd9;
  localparam bridge_masterLogic_fsm_enumDef_STOP3 = 4'd10;
  localparam bridge_masterLogic_fsm_enumDef_TBUF = 4'd11;
  localparam I2cSlaveCmdMode_NONE = 3'd0;
  localparam I2cSlaveCmdMode_START = 3'd1;
  localparam I2cSlaveCmdMode_RESTART = 3'd2;
  localparam I2cSlaveCmdMode_STOP = 3'd3;
  localparam I2cSlaveCmdMode_DROP = 3'd4;
  localparam I2cSlaveCmdMode_DRIVE = 3'd5;
  localparam I2cSlaveCmdMode_READ = 3'd6;

  reg                 i2cCtrl_io_config_timeoutClear;
  reg                 i2cCtrl_io_bus_rsp_valid;
  reg                 i2cCtrl_io_bus_rsp_enable;
  reg                 i2cCtrl_io_bus_rsp_data;
  wire                i2cCtrl_io_i2c_scl_write;
  wire                i2cCtrl_io_i2c_sda_write;
  wire       [2:0]    i2cCtrl_io_bus_cmd_kind;
  wire                i2cCtrl_io_bus_cmd_data;
  wire                i2cCtrl_io_timeout;
  wire                i2cCtrl_io_internals_inFrame;
  wire                i2cCtrl_io_internals_sdaRead;
  wire                i2cCtrl_io_internals_sclRead;
  wire       [6:0]    _zz_bridge_addressFilter_hits_0;
  wire       [6:0]    _zz_bridge_addressFilter_hits_1;
  wire       [0:0]    _zz_bridge_masterLogic_start;
  wire       [0:0]    _zz_bridge_masterLogic_stop;
  wire       [0:0]    _zz_bridge_masterLogic_drop;
  wire       [0:0]    _zz_bridge_masterLogic_recover;
  wire       [11:0]   _zz_bridge_masterLogic_timer_value;
  wire       [0:0]    _zz_bridge_masterLogic_timer_value_1;
  wire       [0:0]    _zz_bridge_masterLogic_fsm_dropped_start;
  wire       [0:0]    _zz_bridge_masterLogic_fsm_dropped_stop;
  wire       [0:0]    _zz_bridge_masterLogic_fsm_dropped_recover;
  wire       [2:0]    _zz_io_bus_rsp_data;
  wire       [2:0]    _zz_bridge_rxData_value;
  wire       [0:0]    _zz_bridge_interruptCtrl_start_flag;
  wire       [0:0]    _zz_bridge_interruptCtrl_restart_flag;
  wire       [0:0]    _zz_bridge_interruptCtrl_end_flag;
  wire       [0:0]    _zz_bridge_interruptCtrl_drop_flag;
  wire       [0:0]    _zz_bridge_interruptCtrl_filterGen_flag;
  wire       [0:0]    _zz_bridge_interruptCtrl_clockGenExit_flag;
  wire       [0:0]    _zz_bridge_interruptCtrl_clockGenEnter_flag;
  wire                busCtrl_readErrorFlag;
  wire                busCtrl_writeErrorFlag;
  wire                busCtrl_readHaltTrigger;
  wire                busCtrl_writeHaltTrigger;
  wire                busCtrl_rsp_valid;
  wire                busCtrl_rsp_ready;
  wire                busCtrl_rsp_payload_last;
  reg        [0:0]    busCtrl_rsp_payload_fragment_opcode;
  reg        [31:0]   busCtrl_rsp_payload_fragment_data;
  wire       [48:0]   busCtrl_rsp_payload_fragment_context;
  wire                _zz_busCtrl_rsp_ready;
  reg                 _zz_busCtrl_rsp_ready_1;
  wire                _zz_io_ctrl_rsp_valid;
  reg                 _zz_io_ctrl_rsp_valid_1;
  reg                 _zz_io_ctrl_rsp_payload_last;
  reg        [0:0]    _zz_io_ctrl_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_ctrl_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_ctrl_rsp_payload_fragment_context;
  wire                when_Stream_l375;
  wire                busCtrl_askWrite;
  wire                busCtrl_askRead;
  wire                io_ctrl_cmd_fire;
  wire                busCtrl_doWrite;
  wire                busCtrl_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  wire                bridge_busCtrlWithOffset_readErrorFlag;
  wire                bridge_busCtrlWithOffset_writeErrorFlag;
  reg                 bridge_frameReset;
  reg                 bridge_i2cBuffer_sda_write;
  wire                bridge_i2cBuffer_sda_read;
  reg                 bridge_i2cBuffer_scl_write;
  wire                bridge_i2cBuffer_scl_read;
  reg                 bridge_rxData_event;
  reg                 bridge_rxData_listen;
  reg                 bridge_rxData_valid;
  reg        [7:0]    bridge_rxData_value;
  reg                 when_I2cCtrl_l224;
  reg                 bridge_rxAck_listen;
  reg                 bridge_rxAck_valid;
  reg                 bridge_rxAck_value;
  reg                 when_I2cCtrl_l237;
  reg                 bridge_txData_valid;
  reg                 bridge_txData_repeat;
  reg                 bridge_txData_enable;
  reg        [7:0]    bridge_txData_value;
  reg                 bridge_txData_forceDisable;
  reg                 bridge_txData_disableOnDataConflict;
  reg                 bridge_txAck_valid;
  reg                 bridge_txAck_repeat;
  reg                 bridge_txAck_enable;
  reg                 bridge_txAck_value;
  reg                 bridge_txAck_forceAck;
  reg                 bridge_txAck_disableOnDataConflict;
  reg                 bridge_addressFilter_addresses_0_enable;
  reg        [9:0]    bridge_addressFilter_addresses_0_value;
  reg                 bridge_addressFilter_addresses_0_is10Bit;
  reg                 bridge_addressFilter_addresses_1_enable;
  reg        [9:0]    bridge_addressFilter_addresses_1_value;
  reg                 bridge_addressFilter_addresses_1_is10Bit;
  reg        [1:0]    bridge_addressFilter_state;
  reg        [7:0]    bridge_addressFilter_byte0;
  reg        [7:0]    bridge_addressFilter_byte1;
  wire                bridge_addressFilter_byte0Is10Bit;
  wire                bridge_addressFilter_hits_0;
  wire                bridge_addressFilter_hits_1;
  wire                when_I2cCtrl_l306;
  wire                _zz_when_I2cCtrl_l310;
  reg                 _zz_when_I2cCtrl_l310_1;
  wire                when_I2cCtrl_l310;
  reg                 bridge_masterLogic_start;
  reg                 when_BusSlaveFactory_l377;
  wire                when_BusSlaveFactory_l379;
  reg                 bridge_masterLogic_stop;
  reg                 when_BusSlaveFactory_l377_1;
  wire                when_BusSlaveFactory_l379_1;
  reg                 bridge_masterLogic_drop;
  reg                 when_BusSlaveFactory_l377_2;
  wire                when_BusSlaveFactory_l379_2;
  reg                 bridge_masterLogic_recover;
  reg                 when_BusSlaveFactory_l377_3;
  wire                when_BusSlaveFactory_l379_3;
  reg        [11:0]   bridge_masterLogic_timer_value;
  reg        [11:0]   bridge_masterLogic_timer_tLow;
  reg        [11:0]   bridge_masterLogic_timer_tHigh;
  reg        [11:0]   bridge_masterLogic_timer_tBuf;
  wire                bridge_masterLogic_timer_done;
  wire                bridge_masterLogic_txReady;
  wire                bridge_masterLogic_fsm_wantExit;
  reg                 bridge_masterLogic_fsm_wantStart;
  wire                bridge_masterLogic_fsm_wantKill;
  reg                 bridge_masterLogic_fsm_dropped_start;
  reg                 bridge_masterLogic_fsm_dropped_stop;
  reg                 bridge_masterLogic_fsm_dropped_recover;
  reg                 bridge_masterLogic_fsm_dropped_trigger;
  reg                 bridge_masterLogic_fsm_inFrameLate;
  wire                when_I2cCtrl_l363;
  wire                when_I2cCtrl_l363_1;
  wire                bridge_masterLogic_fsm_outOfSync;
  wire                bridge_masterLogic_fsm_isBusy;
  reg                 when_BusSlaveFactory_l341;
  wire                when_BusSlaveFactory_l347;
  reg                 when_BusSlaveFactory_l341_1;
  wire                when_BusSlaveFactory_l347_1;
  reg                 when_BusSlaveFactory_l341_2;
  wire                when_BusSlaveFactory_l347_2;
  reg        [2:0]    bridge_dataCounter;
  reg                 bridge_inAckState;
  reg                 bridge_wasntAck;
  wire                when_I2cCtrl_l523;
  wire                when_I2cCtrl_l546;
  wire                when_I2cCtrl_l566;
  wire                when_I2cCtrl_l570;
  wire                when_I2cCtrl_l574;
  wire                when_I2cCtrl_l578;
  wire                when_I2cCtrl_l588;
  wire                when_I2cCtrl_l601;
  reg                 bridge_interruptCtrl_rxDataEnable;
  reg                 bridge_interruptCtrl_rxAckEnable;
  reg                 bridge_interruptCtrl_txDataEnable;
  reg                 bridge_interruptCtrl_txAckEnable;
  reg                 bridge_interruptCtrl_interrupt;
  wire                when_I2cCtrl_l634;
  reg                 bridge_interruptCtrl_start_enable;
  reg                 bridge_interruptCtrl_start_flag;
  wire                when_I2cCtrl_l634_1;
  reg                 when_BusSlaveFactory_l341_3;
  wire                when_BusSlaveFactory_l347_3;
  wire                when_I2cCtrl_l634_2;
  reg                 bridge_interruptCtrl_restart_enable;
  reg                 bridge_interruptCtrl_restart_flag;
  wire                when_I2cCtrl_l634_3;
  reg                 when_BusSlaveFactory_l341_4;
  wire                when_BusSlaveFactory_l347_4;
  wire                when_I2cCtrl_l634_4;
  reg                 bridge_interruptCtrl_end_enable;
  reg                 bridge_interruptCtrl_end_flag;
  wire                when_I2cCtrl_l634_5;
  reg                 when_BusSlaveFactory_l341_5;
  wire                when_BusSlaveFactory_l347_5;
  wire                when_I2cCtrl_l634_6;
  reg                 bridge_interruptCtrl_drop_enable;
  reg                 bridge_interruptCtrl_drop_flag;
  wire                when_I2cCtrl_l634_7;
  reg                 when_BusSlaveFactory_l341_6;
  wire                when_BusSlaveFactory_l347_6;
  wire                _zz_when_I2cCtrl_l634;
  reg                 _zz_when_I2cCtrl_l634_1;
  wire                when_I2cCtrl_l634_8;
  reg                 bridge_interruptCtrl_filterGen_enable;
  reg                 bridge_interruptCtrl_filterGen_flag;
  wire                when_I2cCtrl_l634_9;
  reg                 when_BusSlaveFactory_l341_7;
  wire                when_BusSlaveFactory_l347_7;
  reg                 bridge_masterLogic_fsm_isBusy_regNext;
  wire                when_I2cCtrl_l634_10;
  reg                 bridge_interruptCtrl_clockGenExit_enable;
  reg                 bridge_interruptCtrl_clockGenExit_flag;
  wire                when_I2cCtrl_l634_11;
  reg                 when_BusSlaveFactory_l341_8;
  wire                when_BusSlaveFactory_l347_8;
  reg                 bridge_masterLogic_fsm_isBusy_regNext_1;
  wire                when_I2cCtrl_l634_12;
  reg                 bridge_interruptCtrl_clockGenEnter_enable;
  reg                 bridge_interruptCtrl_clockGenEnter_flag;
  wire                when_I2cCtrl_l634_13;
  reg                 when_BusSlaveFactory_l341_9;
  wire                when_BusSlaveFactory_l347_9;
  reg        [9:0]    _zz_io_config_samplingClockDivider;
  reg        [19:0]   _zz_io_config_timeout;
  reg        [5:0]    _zz_io_config_tsuData;
  reg                 bridge_timeoutClear;
  wire                when_I2cCtrl_l659;
  reg        [3:0]    bridge_masterLogic_fsm_stateReg;
  reg        [3:0]    bridge_masterLogic_fsm_stateNext;
  reg                 i2cCtrl_io_internals_inFrame_regNext;
  wire                when_I2cCtrl_l367;
  wire                when_I2cCtrl_l369;
  wire                when_I2cCtrl_l380;
  wire                when_I2cCtrl_l392;
  wire                when_I2cCtrl_l418;
  wire                when_I2cCtrl_l422;
  wire                when_I2cCtrl_l442;
  wire                when_I2cCtrl_l450;
  wire                when_I2cCtrl_l474;
  wire                when_StateMachine_l253;
  wire                when_StateMachine_l253_1;
  wire                when_StateMachine_l253_2;
  wire                when_StateMachine_l253_3;
  wire                when_StateMachine_l253_4;
  wire                when_StateMachine_l253_5;
  wire                when_I2cCtrl_l350;
  reg                 bridge_slaveOverride_sda;
  reg                 bridge_slaveOverride_scl;
  wire                when_I2cCtrl_l673;
  wire                when_I2cCtrl_l674;
  reg                 bridge_i2cBuffer_scl_write_regNext;
  reg                 bridge_i2cBuffer_sda_write_regNext;
  `ifndef SYNTHESIS
  reg [55:0] bridge_masterLogic_fsm_stateReg_string;
  reg [55:0] bridge_masterLogic_fsm_stateNext_string;
  `endif


  assign _zz_bridge_addressFilter_hits_0 = (bridge_addressFilter_byte0 >>> 1'd1);
  assign _zz_bridge_addressFilter_hits_1 = (bridge_addressFilter_byte0 >>> 1'd1);
  assign _zz_bridge_masterLogic_start = 1'b1;
  assign _zz_bridge_masterLogic_stop = 1'b1;
  assign _zz_bridge_masterLogic_drop = 1'b1;
  assign _zz_bridge_masterLogic_recover = 1'b1;
  assign _zz_bridge_masterLogic_timer_value_1 = (! bridge_masterLogic_timer_done);
  assign _zz_bridge_masterLogic_timer_value = {11'd0, _zz_bridge_masterLogic_timer_value_1};
  assign _zz_bridge_masterLogic_fsm_dropped_start = 1'b0;
  assign _zz_bridge_masterLogic_fsm_dropped_stop = 1'b0;
  assign _zz_bridge_masterLogic_fsm_dropped_recover = 1'b0;
  assign _zz_io_bus_rsp_data = (3'b111 - bridge_dataCounter);
  assign _zz_bridge_rxData_value = (3'b111 - bridge_dataCounter);
  assign _zz_bridge_interruptCtrl_start_flag = 1'b0;
  assign _zz_bridge_interruptCtrl_restart_flag = 1'b0;
  assign _zz_bridge_interruptCtrl_end_flag = 1'b0;
  assign _zz_bridge_interruptCtrl_drop_flag = 1'b0;
  assign _zz_bridge_interruptCtrl_filterGen_flag = 1'b0;
  assign _zz_bridge_interruptCtrl_clockGenExit_flag = 1'b0;
  assign _zz_bridge_interruptCtrl_clockGenEnter_flag = 1'b0;
  I2cSlave i2cCtrl (
    .io_i2c_sda_write               (i2cCtrl_io_i2c_sda_write               ), //o
    .io_i2c_sda_read                (bridge_i2cBuffer_sda_read              ), //i
    .io_i2c_scl_write               (i2cCtrl_io_i2c_scl_write               ), //o
    .io_i2c_scl_read                (bridge_i2cBuffer_scl_read              ), //i
    .io_config_samplingClockDivider (_zz_io_config_samplingClockDivider[9:0]), //i
    .io_config_timeout              (_zz_io_config_timeout[19:0]            ), //i
    .io_config_tsuData              (_zz_io_config_tsuData[5:0]             ), //i
    .io_config_timeoutClear         (i2cCtrl_io_config_timeoutClear         ), //i
    .io_bus_cmd_kind                (i2cCtrl_io_bus_cmd_kind[2:0]           ), //o
    .io_bus_cmd_data                (i2cCtrl_io_bus_cmd_data                ), //o
    .io_bus_rsp_valid               (i2cCtrl_io_bus_rsp_valid               ), //i
    .io_bus_rsp_enable              (i2cCtrl_io_bus_rsp_enable              ), //i
    .io_bus_rsp_data                (i2cCtrl_io_bus_rsp_data                ), //i
    .io_timeout                     (i2cCtrl_io_timeout                     ), //o
    .io_internals_inFrame           (i2cCtrl_io_internals_inFrame           ), //o
    .io_internals_sdaRead           (i2cCtrl_io_internals_sdaRead           ), //o
    .io_internals_sclRead           (i2cCtrl_io_internals_sclRead           ), //o
    .io_peripheralClk               (io_peripheralClk                       ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset         )  //i
  );
  initial begin
  `ifndef SYNTHESIS
    _zz_io_config_timeout = {$urandom};
    _zz_io_config_tsuData = {$urandom};
  `endif
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(bridge_masterLogic_fsm_stateReg)
      bridge_masterLogic_fsm_enumDef_BOOT : bridge_masterLogic_fsm_stateReg_string = "BOOT   ";
      bridge_masterLogic_fsm_enumDef_IDLE : bridge_masterLogic_fsm_stateReg_string = "IDLE   ";
      bridge_masterLogic_fsm_enumDef_START1 : bridge_masterLogic_fsm_stateReg_string = "START1 ";
      bridge_masterLogic_fsm_enumDef_START2 : bridge_masterLogic_fsm_stateReg_string = "START2 ";
      bridge_masterLogic_fsm_enumDef_START3 : bridge_masterLogic_fsm_stateReg_string = "START3 ";
      bridge_masterLogic_fsm_enumDef_LOW : bridge_masterLogic_fsm_stateReg_string = "LOW    ";
      bridge_masterLogic_fsm_enumDef_HIGH : bridge_masterLogic_fsm_stateReg_string = "HIGH   ";
      bridge_masterLogic_fsm_enumDef_RESTART : bridge_masterLogic_fsm_stateReg_string = "RESTART";
      bridge_masterLogic_fsm_enumDef_STOP1 : bridge_masterLogic_fsm_stateReg_string = "STOP1  ";
      bridge_masterLogic_fsm_enumDef_STOP2 : bridge_masterLogic_fsm_stateReg_string = "STOP2  ";
      bridge_masterLogic_fsm_enumDef_STOP3 : bridge_masterLogic_fsm_stateReg_string = "STOP3  ";
      bridge_masterLogic_fsm_enumDef_TBUF : bridge_masterLogic_fsm_stateReg_string = "TBUF   ";
      default : bridge_masterLogic_fsm_stateReg_string = "???????";
    endcase
  end
  always @(*) begin
    case(bridge_masterLogic_fsm_stateNext)
      bridge_masterLogic_fsm_enumDef_BOOT : bridge_masterLogic_fsm_stateNext_string = "BOOT   ";
      bridge_masterLogic_fsm_enumDef_IDLE : bridge_masterLogic_fsm_stateNext_string = "IDLE   ";
      bridge_masterLogic_fsm_enumDef_START1 : bridge_masterLogic_fsm_stateNext_string = "START1 ";
      bridge_masterLogic_fsm_enumDef_START2 : bridge_masterLogic_fsm_stateNext_string = "START2 ";
      bridge_masterLogic_fsm_enumDef_START3 : bridge_masterLogic_fsm_stateNext_string = "START3 ";
      bridge_masterLogic_fsm_enumDef_LOW : bridge_masterLogic_fsm_stateNext_string = "LOW    ";
      bridge_masterLogic_fsm_enumDef_HIGH : bridge_masterLogic_fsm_stateNext_string = "HIGH   ";
      bridge_masterLogic_fsm_enumDef_RESTART : bridge_masterLogic_fsm_stateNext_string = "RESTART";
      bridge_masterLogic_fsm_enumDef_STOP1 : bridge_masterLogic_fsm_stateNext_string = "STOP1  ";
      bridge_masterLogic_fsm_enumDef_STOP2 : bridge_masterLogic_fsm_stateNext_string = "STOP2  ";
      bridge_masterLogic_fsm_enumDef_STOP3 : bridge_masterLogic_fsm_stateNext_string = "STOP3  ";
      bridge_masterLogic_fsm_enumDef_TBUF : bridge_masterLogic_fsm_stateNext_string = "TBUF   ";
      default : bridge_masterLogic_fsm_stateNext_string = "???????";
    endcase
  end
  `endif

  assign busCtrl_readErrorFlag = 1'b0;
  assign busCtrl_writeErrorFlag = 1'b0;
  assign busCtrl_readHaltTrigger = 1'b0;
  assign busCtrl_writeHaltTrigger = 1'b0;
  assign _zz_busCtrl_rsp_ready = (! (busCtrl_readHaltTrigger || busCtrl_writeHaltTrigger));
  assign busCtrl_rsp_ready = (_zz_busCtrl_rsp_ready_1 && _zz_busCtrl_rsp_ready);
  always @(*) begin
    _zz_busCtrl_rsp_ready_1 = io_ctrl_rsp_ready;
    if(when_Stream_l375) begin
      _zz_busCtrl_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375 = (! _zz_io_ctrl_rsp_valid);
  assign _zz_io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid_1;
  assign io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid;
  assign io_ctrl_rsp_payload_last = _zz_io_ctrl_rsp_payload_last;
  assign io_ctrl_rsp_payload_fragment_opcode = _zz_io_ctrl_rsp_payload_fragment_opcode;
  assign io_ctrl_rsp_payload_fragment_data = _zz_io_ctrl_rsp_payload_fragment_data;
  assign io_ctrl_rsp_payload_fragment_context = _zz_io_ctrl_rsp_payload_fragment_context;
  assign busCtrl_askWrite = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_askRead = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign io_ctrl_cmd_fire = (io_ctrl_cmd_valid && io_ctrl_cmd_ready);
  assign busCtrl_doWrite = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_doRead = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign busCtrl_rsp_valid = io_ctrl_cmd_valid;
  assign io_ctrl_cmd_ready = busCtrl_rsp_ready;
  assign busCtrl_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (busCtrl_doWrite && busCtrl_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      busCtrl_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        busCtrl_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        busCtrl_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (busCtrl_doRead && busCtrl_readErrorFlag);
  always @(*) begin
    busCtrl_rsp_payload_fragment_data = 32'h0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h08 : begin
        busCtrl_rsp_payload_fragment_data[8 : 8] = bridge_rxData_valid;
        busCtrl_rsp_payload_fragment_data[7 : 0] = bridge_rxData_value;
      end
      8'h0c : begin
        busCtrl_rsp_payload_fragment_data[8 : 8] = bridge_rxAck_valid;
        busCtrl_rsp_payload_fragment_data[0 : 0] = bridge_rxAck_value;
      end
      8'h0 : begin
        busCtrl_rsp_payload_fragment_data[8 : 8] = bridge_txData_valid;
        busCtrl_rsp_payload_fragment_data[9 : 9] = bridge_txData_enable;
      end
      8'h04 : begin
        busCtrl_rsp_payload_fragment_data[8 : 8] = bridge_txAck_valid;
        busCtrl_rsp_payload_fragment_data[9 : 9] = bridge_txAck_enable;
      end
      8'h80 : begin
        busCtrl_rsp_payload_fragment_data[1 : 0] = {bridge_addressFilter_hits_1,bridge_addressFilter_hits_0};
      end
      8'h84 : begin
        busCtrl_rsp_payload_fragment_data[0 : 0] = bridge_addressFilter_byte0[0];
      end
      8'h40 : begin
        busCtrl_rsp_payload_fragment_data[4 : 4] = bridge_masterLogic_start;
        busCtrl_rsp_payload_fragment_data[5 : 5] = bridge_masterLogic_stop;
        busCtrl_rsp_payload_fragment_data[6 : 6] = bridge_masterLogic_drop;
        busCtrl_rsp_payload_fragment_data[7 : 7] = bridge_masterLogic_recover;
        busCtrl_rsp_payload_fragment_data[0 : 0] = bridge_masterLogic_fsm_isBusy;
        busCtrl_rsp_payload_fragment_data[9 : 9] = bridge_masterLogic_fsm_dropped_start;
        busCtrl_rsp_payload_fragment_data[10 : 10] = bridge_masterLogic_fsm_dropped_stop;
        busCtrl_rsp_payload_fragment_data[11 : 11] = bridge_masterLogic_fsm_dropped_recover;
      end
      8'h20 : begin
        busCtrl_rsp_payload_fragment_data[0 : 0] = bridge_interruptCtrl_rxDataEnable;
        busCtrl_rsp_payload_fragment_data[1 : 1] = bridge_interruptCtrl_rxAckEnable;
        busCtrl_rsp_payload_fragment_data[2 : 2] = bridge_interruptCtrl_txDataEnable;
        busCtrl_rsp_payload_fragment_data[3 : 3] = bridge_interruptCtrl_txAckEnable;
        busCtrl_rsp_payload_fragment_data[4 : 4] = bridge_interruptCtrl_start_enable;
        busCtrl_rsp_payload_fragment_data[5 : 5] = bridge_interruptCtrl_restart_enable;
        busCtrl_rsp_payload_fragment_data[6 : 6] = bridge_interruptCtrl_end_enable;
        busCtrl_rsp_payload_fragment_data[7 : 7] = bridge_interruptCtrl_drop_enable;
        busCtrl_rsp_payload_fragment_data[17 : 17] = bridge_interruptCtrl_filterGen_enable;
        busCtrl_rsp_payload_fragment_data[15 : 15] = bridge_interruptCtrl_clockGenExit_enable;
        busCtrl_rsp_payload_fragment_data[16 : 16] = bridge_interruptCtrl_clockGenEnter_enable;
      end
      8'h24 : begin
        busCtrl_rsp_payload_fragment_data[4 : 4] = bridge_interruptCtrl_start_flag;
        busCtrl_rsp_payload_fragment_data[5 : 5] = bridge_interruptCtrl_restart_flag;
        busCtrl_rsp_payload_fragment_data[6 : 6] = bridge_interruptCtrl_end_flag;
        busCtrl_rsp_payload_fragment_data[7 : 7] = bridge_interruptCtrl_drop_flag;
        busCtrl_rsp_payload_fragment_data[17 : 17] = bridge_interruptCtrl_filterGen_flag;
        busCtrl_rsp_payload_fragment_data[15 : 15] = bridge_interruptCtrl_clockGenExit_flag;
        busCtrl_rsp_payload_fragment_data[16 : 16] = bridge_interruptCtrl_clockGenEnter_flag;
      end
      8'h44 : begin
        busCtrl_rsp_payload_fragment_data[0 : 0] = i2cCtrl_io_internals_inFrame;
        busCtrl_rsp_payload_fragment_data[1 : 1] = i2cCtrl_io_internals_sdaRead;
        busCtrl_rsp_payload_fragment_data[2 : 2] = i2cCtrl_io_internals_sclRead;
      end
      8'h48 : begin
        busCtrl_rsp_payload_fragment_data[1 : 1] = bridge_slaveOverride_sda;
        busCtrl_rsp_payload_fragment_data[2 : 2] = bridge_slaveOverride_scl;
      end
      default : begin
      end
    endcase
  end

  assign busCtrl_rsp_payload_fragment_context = io_ctrl_cmd_payload_fragment_context;
  assign bridge_busCtrlWithOffset_readErrorFlag = 1'b0;
  assign bridge_busCtrlWithOffset_writeErrorFlag = 1'b0;
  always @(*) begin
    bridge_frameReset = 1'b0;
    case(i2cCtrl_io_bus_cmd_kind)
      I2cSlaveCmdMode_START : begin
        bridge_frameReset = 1'b1;
      end
      I2cSlaveCmdMode_RESTART : begin
        bridge_frameReset = 1'b1;
      end
      I2cSlaveCmdMode_STOP : begin
        bridge_frameReset = 1'b1;
      end
      I2cSlaveCmdMode_DROP : begin
        bridge_frameReset = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bridge_i2cBuffer_sda_write = i2cCtrl_io_i2c_sda_write;
    case(bridge_masterLogic_fsm_stateReg)
      bridge_masterLogic_fsm_enumDef_IDLE : begin
      end
      bridge_masterLogic_fsm_enumDef_START1 : begin
      end
      bridge_masterLogic_fsm_enumDef_START2 : begin
        bridge_i2cBuffer_sda_write = 1'b0;
      end
      bridge_masterLogic_fsm_enumDef_START3 : begin
        bridge_i2cBuffer_sda_write = 1'b0;
      end
      bridge_masterLogic_fsm_enumDef_LOW : begin
      end
      bridge_masterLogic_fsm_enumDef_HIGH : begin
      end
      bridge_masterLogic_fsm_enumDef_RESTART : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP1 : begin
        bridge_i2cBuffer_sda_write = 1'b0;
      end
      bridge_masterLogic_fsm_enumDef_STOP2 : begin
        bridge_i2cBuffer_sda_write = 1'b0;
      end
      bridge_masterLogic_fsm_enumDef_STOP3 : begin
      end
      bridge_masterLogic_fsm_enumDef_TBUF : begin
      end
      default : begin
      end
    endcase
    if(when_I2cCtrl_l673) begin
      bridge_i2cBuffer_sda_write = 1'b0;
    end
  end

  always @(*) begin
    bridge_i2cBuffer_scl_write = i2cCtrl_io_i2c_scl_write;
    case(bridge_masterLogic_fsm_stateReg)
      bridge_masterLogic_fsm_enumDef_IDLE : begin
      end
      bridge_masterLogic_fsm_enumDef_START1 : begin
      end
      bridge_masterLogic_fsm_enumDef_START2 : begin
      end
      bridge_masterLogic_fsm_enumDef_START3 : begin
        bridge_i2cBuffer_scl_write = 1'b0;
      end
      bridge_masterLogic_fsm_enumDef_LOW : begin
        if(bridge_masterLogic_timer_done) begin
          if(when_I2cCtrl_l418) begin
            bridge_i2cBuffer_scl_write = 1'b0;
          end else begin
            if(when_I2cCtrl_l422) begin
              bridge_i2cBuffer_scl_write = 1'b0;
            end
          end
        end else begin
          bridge_i2cBuffer_scl_write = 1'b0;
        end
      end
      bridge_masterLogic_fsm_enumDef_HIGH : begin
      end
      bridge_masterLogic_fsm_enumDef_RESTART : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP1 : begin
        bridge_i2cBuffer_scl_write = 1'b0;
      end
      bridge_masterLogic_fsm_enumDef_STOP2 : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP3 : begin
      end
      bridge_masterLogic_fsm_enumDef_TBUF : begin
      end
      default : begin
      end
    endcase
    if(when_I2cCtrl_l674) begin
      bridge_i2cBuffer_scl_write = 1'b0;
    end
  end

  always @(*) begin
    when_I2cCtrl_l224 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h08 : begin
        if(busCtrl_doRead) begin
          when_I2cCtrl_l224 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    when_I2cCtrl_l237 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h0c : begin
        if(busCtrl_doRead) begin
          when_I2cCtrl_l237 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bridge_txData_forceDisable = 1'b0;
    if(when_I2cCtrl_l601) begin
      bridge_txData_forceDisable = 1'b0;
    end
    case(bridge_masterLogic_fsm_stateReg)
      bridge_masterLogic_fsm_enumDef_IDLE : begin
      end
      bridge_masterLogic_fsm_enumDef_START1 : begin
      end
      bridge_masterLogic_fsm_enumDef_START2 : begin
      end
      bridge_masterLogic_fsm_enumDef_START3 : begin
      end
      bridge_masterLogic_fsm_enumDef_LOW : begin
        if(bridge_masterLogic_timer_done) begin
          if(when_I2cCtrl_l418) begin
            bridge_txData_forceDisable = 1'b1;
          end else begin
            if(when_I2cCtrl_l422) begin
              bridge_txData_forceDisable = 1'b1;
            end
          end
        end
      end
      bridge_masterLogic_fsm_enumDef_HIGH : begin
      end
      bridge_masterLogic_fsm_enumDef_RESTART : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP1 : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP2 : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP3 : begin
      end
      bridge_masterLogic_fsm_enumDef_TBUF : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bridge_txAck_forceAck = 1'b0;
    if(when_I2cCtrl_l306) begin
      bridge_txAck_forceAck = 1'b1;
    end
  end

  assign bridge_addressFilter_byte0Is10Bit = (bridge_addressFilter_byte0[7 : 3] == 5'h1e);
  assign bridge_addressFilter_hits_0 = (bridge_addressFilter_addresses_0_enable && ((! bridge_addressFilter_addresses_0_is10Bit) ? ((_zz_bridge_addressFilter_hits_0 == bridge_addressFilter_addresses_0_value[6 : 0]) && (bridge_addressFilter_state != 2'b00)) : (({bridge_addressFilter_byte0[2 : 1],bridge_addressFilter_byte1} == bridge_addressFilter_addresses_0_value) && (bridge_addressFilter_state == 2'b10))));
  assign bridge_addressFilter_hits_1 = (bridge_addressFilter_addresses_1_enable && ((! bridge_addressFilter_addresses_1_is10Bit) ? ((_zz_bridge_addressFilter_hits_1 == bridge_addressFilter_addresses_1_value[6 : 0]) && (bridge_addressFilter_state != 2'b00)) : (({bridge_addressFilter_byte0[2 : 1],bridge_addressFilter_byte1} == bridge_addressFilter_addresses_1_value) && (bridge_addressFilter_state == 2'b10))));
  assign when_I2cCtrl_l306 = ((bridge_addressFilter_byte0Is10Bit && (bridge_addressFilter_state == 2'b01)) && (|{((bridge_addressFilter_addresses_1_enable && bridge_addressFilter_addresses_1_is10Bit) && (bridge_addressFilter_byte0[2 : 1] == bridge_addressFilter_addresses_1_value[9 : 8])),((bridge_addressFilter_addresses_0_enable && bridge_addressFilter_addresses_0_is10Bit) && (bridge_addressFilter_byte0[2 : 1] == bridge_addressFilter_addresses_0_value[9 : 8]))}));
  assign _zz_when_I2cCtrl_l310 = (|{bridge_addressFilter_hits_1,bridge_addressFilter_hits_0});
  assign when_I2cCtrl_l310 = (_zz_when_I2cCtrl_l310 && (! _zz_when_I2cCtrl_l310_1));
  always @(*) begin
    when_BusSlaveFactory_l377 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h40 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l377 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379 = io_ctrl_cmd_payload_fragment_data[4];
  always @(*) begin
    when_BusSlaveFactory_l377_1 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h40 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l377_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_1 = io_ctrl_cmd_payload_fragment_data[5];
  always @(*) begin
    when_BusSlaveFactory_l377_2 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h40 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l377_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_2 = io_ctrl_cmd_payload_fragment_data[6];
  always @(*) begin
    when_BusSlaveFactory_l377_3 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h40 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l377_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_3 = io_ctrl_cmd_payload_fragment_data[7];
  assign bridge_masterLogic_timer_done = (bridge_masterLogic_timer_value == 12'h0);
  assign bridge_masterLogic_fsm_wantExit = 1'b0;
  always @(*) begin
    bridge_masterLogic_fsm_wantStart = 1'b0;
    case(bridge_masterLogic_fsm_stateReg)
      bridge_masterLogic_fsm_enumDef_IDLE : begin
      end
      bridge_masterLogic_fsm_enumDef_START1 : begin
      end
      bridge_masterLogic_fsm_enumDef_START2 : begin
      end
      bridge_masterLogic_fsm_enumDef_START3 : begin
      end
      bridge_masterLogic_fsm_enumDef_LOW : begin
      end
      bridge_masterLogic_fsm_enumDef_HIGH : begin
      end
      bridge_masterLogic_fsm_enumDef_RESTART : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP1 : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP2 : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP3 : begin
      end
      bridge_masterLogic_fsm_enumDef_TBUF : begin
      end
      default : begin
        bridge_masterLogic_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign bridge_masterLogic_fsm_wantKill = 1'b0;
  always @(*) begin
    bridge_masterLogic_fsm_dropped_trigger = 1'b0;
    if(when_I2cCtrl_l350) begin
      bridge_masterLogic_fsm_dropped_trigger = 1'b1;
    end
  end

  assign when_I2cCtrl_l363 = (! i2cCtrl_io_internals_sclRead);
  assign when_I2cCtrl_l363_1 = (! i2cCtrl_io_internals_inFrame);
  assign bridge_masterLogic_fsm_outOfSync = ((! i2cCtrl_io_internals_inFrame) && ((! i2cCtrl_io_internals_sdaRead) || (! i2cCtrl_io_internals_sclRead)));
  assign bridge_masterLogic_fsm_isBusy = ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_IDLE)) && (! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_TBUF)));
  always @(*) begin
    when_BusSlaveFactory_l341 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h40 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347 = io_ctrl_cmd_payload_fragment_data[9];
  always @(*) begin
    when_BusSlaveFactory_l341_1 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h40 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_1 = io_ctrl_cmd_payload_fragment_data[10];
  always @(*) begin
    when_BusSlaveFactory_l341_2 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h40 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_2 = io_ctrl_cmd_payload_fragment_data[11];
  assign bridge_masterLogic_txReady = (bridge_inAckState ? bridge_txAck_valid : bridge_txData_valid);
  assign when_I2cCtrl_l523 = (! bridge_inAckState);
  always @(*) begin
    if(when_I2cCtrl_l523) begin
      i2cCtrl_io_bus_rsp_valid = ((bridge_txData_valid && (! (bridge_rxData_valid && bridge_rxData_listen))) && (i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_DRIVE));
      if(bridge_txData_forceDisable) begin
        i2cCtrl_io_bus_rsp_valid = 1'b1;
      end
    end else begin
      i2cCtrl_io_bus_rsp_valid = ((bridge_txAck_valid && (! (bridge_rxAck_valid && bridge_rxAck_listen))) && (i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_DRIVE));
      if(bridge_txAck_forceAck) begin
        i2cCtrl_io_bus_rsp_valid = 1'b1;
      end
    end
    if(when_I2cCtrl_l546) begin
      i2cCtrl_io_bus_rsp_valid = (i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_DRIVE);
    end
  end

  always @(*) begin
    if(when_I2cCtrl_l523) begin
      i2cCtrl_io_bus_rsp_enable = bridge_txData_enable;
      if(bridge_txData_forceDisable) begin
        i2cCtrl_io_bus_rsp_enable = 1'b0;
      end
    end else begin
      i2cCtrl_io_bus_rsp_enable = bridge_txAck_enable;
      if(bridge_txAck_forceAck) begin
        i2cCtrl_io_bus_rsp_enable = 1'b1;
      end
    end
    if(when_I2cCtrl_l546) begin
      i2cCtrl_io_bus_rsp_enable = 1'b0;
    end
  end

  always @(*) begin
    if(when_I2cCtrl_l523) begin
      i2cCtrl_io_bus_rsp_data = bridge_txData_value[_zz_io_bus_rsp_data];
    end else begin
      i2cCtrl_io_bus_rsp_data = bridge_txAck_value;
      if(bridge_txAck_forceAck) begin
        i2cCtrl_io_bus_rsp_data = 1'b0;
      end
    end
  end

  assign when_I2cCtrl_l546 = (bridge_wasntAck && (! bridge_masterLogic_fsm_isBusy));
  assign when_I2cCtrl_l566 = (! bridge_inAckState);
  assign when_I2cCtrl_l570 = (i2cCtrl_io_bus_rsp_data != i2cCtrl_io_bus_cmd_data);
  assign when_I2cCtrl_l574 = (bridge_dataCounter == 3'b111);
  assign when_I2cCtrl_l578 = (bridge_txData_valid && (! bridge_txData_repeat));
  assign when_I2cCtrl_l588 = (bridge_txAck_valid && (! bridge_txAck_repeat));
  assign when_I2cCtrl_l601 = ((i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_STOP) || (i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_DROP));
  always @(*) begin
    bridge_interruptCtrl_interrupt = ((((bridge_interruptCtrl_rxDataEnable && bridge_rxData_valid) || (bridge_interruptCtrl_rxAckEnable && bridge_rxAck_valid)) || (bridge_interruptCtrl_txDataEnable && (! bridge_txData_valid))) || (bridge_interruptCtrl_txAckEnable && (! bridge_txAck_valid)));
    if(bridge_interruptCtrl_start_flag) begin
      bridge_interruptCtrl_interrupt = 1'b1;
    end
    if(bridge_interruptCtrl_restart_flag) begin
      bridge_interruptCtrl_interrupt = 1'b1;
    end
    if(bridge_interruptCtrl_end_flag) begin
      bridge_interruptCtrl_interrupt = 1'b1;
    end
    if(bridge_interruptCtrl_drop_flag) begin
      bridge_interruptCtrl_interrupt = 1'b1;
    end
    if(bridge_interruptCtrl_filterGen_flag) begin
      bridge_interruptCtrl_interrupt = 1'b1;
    end
    if(bridge_interruptCtrl_clockGenExit_flag) begin
      bridge_interruptCtrl_interrupt = 1'b1;
    end
    if(bridge_interruptCtrl_clockGenEnter_flag) begin
      bridge_interruptCtrl_interrupt = 1'b1;
    end
  end

  assign when_I2cCtrl_l634 = (i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_START);
  assign when_I2cCtrl_l634_1 = (! bridge_interruptCtrl_start_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_3 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h24 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_3 = io_ctrl_cmd_payload_fragment_data[4];
  assign when_I2cCtrl_l634_2 = (i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_RESTART);
  assign when_I2cCtrl_l634_3 = (! bridge_interruptCtrl_restart_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_4 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h24 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_4 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_4 = io_ctrl_cmd_payload_fragment_data[5];
  assign when_I2cCtrl_l634_4 = (i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_STOP);
  assign when_I2cCtrl_l634_5 = (! bridge_interruptCtrl_end_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_5 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h24 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_5 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_5 = io_ctrl_cmd_payload_fragment_data[6];
  assign when_I2cCtrl_l634_6 = ((i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_DROP) || bridge_masterLogic_fsm_dropped_trigger);
  assign when_I2cCtrl_l634_7 = (! bridge_interruptCtrl_drop_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_6 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h24 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_6 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_6 = io_ctrl_cmd_payload_fragment_data[7];
  assign _zz_when_I2cCtrl_l634 = (|{bridge_addressFilter_hits_1,bridge_addressFilter_hits_0});
  assign when_I2cCtrl_l634_8 = (_zz_when_I2cCtrl_l634 && (! _zz_when_I2cCtrl_l634_1));
  assign when_I2cCtrl_l634_9 = (! bridge_interruptCtrl_filterGen_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_7 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h24 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_7 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_7 = io_ctrl_cmd_payload_fragment_data[17];
  assign when_I2cCtrl_l634_10 = ((! bridge_masterLogic_fsm_isBusy) && bridge_masterLogic_fsm_isBusy_regNext);
  assign when_I2cCtrl_l634_11 = (! bridge_interruptCtrl_clockGenExit_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_8 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h24 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_8 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_8 = io_ctrl_cmd_payload_fragment_data[15];
  assign when_I2cCtrl_l634_12 = (bridge_masterLogic_fsm_isBusy && (! bridge_masterLogic_fsm_isBusy_regNext_1));
  assign when_I2cCtrl_l634_13 = (! bridge_interruptCtrl_clockGenEnter_enable);
  always @(*) begin
    when_BusSlaveFactory_l341_9 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      8'h24 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_9 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_9 = io_ctrl_cmd_payload_fragment_data[16];
  always @(*) begin
    i2cCtrl_io_config_timeoutClear = bridge_timeoutClear;
    if(when_I2cCtrl_l659) begin
      i2cCtrl_io_config_timeoutClear = 1'b1;
    end
  end

  assign when_I2cCtrl_l659 = ((! i2cCtrl_io_internals_inFrame) && (! bridge_masterLogic_fsm_isBusy));
  always @(*) begin
    bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_stateReg;
    case(bridge_masterLogic_fsm_stateReg)
      bridge_masterLogic_fsm_enumDef_IDLE : begin
        if(when_I2cCtrl_l367) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_TBUF;
        end else begin
          if(when_I2cCtrl_l369) begin
            bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_START1;
          end else begin
            if(bridge_masterLogic_recover) begin
              bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_LOW;
            end
          end
        end
      end
      bridge_masterLogic_fsm_enumDef_START1 : begin
        if(when_I2cCtrl_l380) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_START2;
        end
      end
      bridge_masterLogic_fsm_enumDef_START2 : begin
        if(when_I2cCtrl_l392) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_START3;
        end
      end
      bridge_masterLogic_fsm_enumDef_START3 : begin
        if(bridge_masterLogic_timer_done) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_LOW;
        end
      end
      bridge_masterLogic_fsm_enumDef_LOW : begin
        if(bridge_masterLogic_timer_done) begin
          if(when_I2cCtrl_l418) begin
            bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_STOP1;
          end else begin
            if(when_I2cCtrl_l422) begin
              bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_RESTART;
            end else begin
              if(i2cCtrl_io_internals_sclRead) begin
                bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_HIGH;
              end
            end
          end
        end
      end
      bridge_masterLogic_fsm_enumDef_HIGH : begin
        if(when_I2cCtrl_l442) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_LOW;
        end
      end
      bridge_masterLogic_fsm_enumDef_RESTART : begin
        if(!when_I2cCtrl_l450) begin
          if(bridge_masterLogic_timer_done) begin
            bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_START1;
          end
        end
      end
      bridge_masterLogic_fsm_enumDef_STOP1 : begin
        if(bridge_masterLogic_timer_done) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_STOP2;
        end
      end
      bridge_masterLogic_fsm_enumDef_STOP2 : begin
        if(!when_I2cCtrl_l474) begin
          if(bridge_masterLogic_timer_done) begin
            bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_STOP3;
          end
        end
      end
      bridge_masterLogic_fsm_enumDef_STOP3 : begin
        if(i2cCtrl_io_internals_sdaRead) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_TBUF;
        end
      end
      bridge_masterLogic_fsm_enumDef_TBUF : begin
        if(bridge_masterLogic_timer_done) begin
          bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(when_I2cCtrl_l350) begin
      bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_TBUF;
    end
    if(bridge_masterLogic_fsm_wantStart) begin
      bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_IDLE;
    end
    if(bridge_masterLogic_fsm_wantKill) begin
      bridge_masterLogic_fsm_stateNext = bridge_masterLogic_fsm_enumDef_BOOT;
    end
  end

  assign when_I2cCtrl_l367 = ((! i2cCtrl_io_internals_inFrame) && i2cCtrl_io_internals_inFrame_regNext);
  assign when_I2cCtrl_l369 = (bridge_masterLogic_start && (! bridge_masterLogic_fsm_inFrameLate));
  assign when_I2cCtrl_l380 = (! bridge_masterLogic_fsm_outOfSync);
  assign when_I2cCtrl_l392 = (bridge_masterLogic_timer_done || (! i2cCtrl_io_internals_sclRead));
  assign when_I2cCtrl_l418 = ((bridge_masterLogic_stop && (! bridge_inAckState)) || (bridge_masterLogic_recover && i2cCtrl_io_internals_sdaRead));
  assign when_I2cCtrl_l422 = (bridge_masterLogic_start && (! bridge_inAckState));
  assign when_I2cCtrl_l442 = (bridge_masterLogic_timer_done || (! i2cCtrl_io_internals_sclRead));
  assign when_I2cCtrl_l450 = (! i2cCtrl_io_internals_sclRead);
  assign when_I2cCtrl_l474 = (! i2cCtrl_io_internals_sclRead);
  assign when_StateMachine_l253 = ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_START2)) && (bridge_masterLogic_fsm_stateNext == bridge_masterLogic_fsm_enumDef_START2));
  assign when_StateMachine_l253_1 = ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_START3)) && (bridge_masterLogic_fsm_stateNext == bridge_masterLogic_fsm_enumDef_START3));
  assign when_StateMachine_l253_2 = ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_LOW)) && (bridge_masterLogic_fsm_stateNext == bridge_masterLogic_fsm_enumDef_LOW));
  assign when_StateMachine_l253_3 = ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_HIGH)) && (bridge_masterLogic_fsm_stateNext == bridge_masterLogic_fsm_enumDef_HIGH));
  assign when_StateMachine_l253_4 = ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_STOP1)) && (bridge_masterLogic_fsm_stateNext == bridge_masterLogic_fsm_enumDef_STOP1));
  assign when_StateMachine_l253_5 = ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_TBUF)) && (bridge_masterLogic_fsm_stateNext == bridge_masterLogic_fsm_enumDef_TBUF));
  assign when_I2cCtrl_l350 = (bridge_masterLogic_drop || ((! (bridge_masterLogic_fsm_stateReg == bridge_masterLogic_fsm_enumDef_IDLE)) && ((i2cCtrl_io_bus_cmd_kind == I2cSlaveCmdMode_DROP) || i2cCtrl_io_timeout)));
  assign when_I2cCtrl_l673 = (! bridge_slaveOverride_sda);
  assign when_I2cCtrl_l674 = (! bridge_slaveOverride_scl);
  assign io_i2c_scl_write = bridge_i2cBuffer_scl_write_regNext;
  assign io_i2c_sda_write = bridge_i2cBuffer_sda_write_regNext;
  assign bridge_i2cBuffer_scl_read = io_i2c_scl_read;
  assign bridge_i2cBuffer_sda_read = io_i2c_sda_read;
  assign io_interrupt = bridge_interruptCtrl_interrupt;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      _zz_io_ctrl_rsp_valid_1 <= 1'b0;
      bridge_rxData_event <= 1'b0;
      bridge_rxData_listen <= 1'b0;
      bridge_rxData_valid <= 1'b0;
      bridge_rxAck_listen <= 1'b0;
      bridge_rxAck_valid <= 1'b0;
      bridge_txData_valid <= 1'b1;
      bridge_txData_repeat <= 1'b1;
      bridge_txData_enable <= 1'b0;
      bridge_txAck_valid <= 1'b1;
      bridge_txAck_repeat <= 1'b1;
      bridge_txAck_enable <= 1'b0;
      bridge_addressFilter_addresses_0_enable <= 1'b0;
      bridge_addressFilter_addresses_1_enable <= 1'b0;
      bridge_addressFilter_state <= 2'b00;
      bridge_masterLogic_start <= 1'b0;
      bridge_masterLogic_stop <= 1'b0;
      bridge_masterLogic_drop <= 1'b0;
      bridge_masterLogic_recover <= 1'b0;
      bridge_masterLogic_fsm_dropped_start <= 1'b0;
      bridge_masterLogic_fsm_dropped_stop <= 1'b0;
      bridge_masterLogic_fsm_dropped_recover <= 1'b0;
      bridge_dataCounter <= 3'b000;
      bridge_inAckState <= 1'b0;
      bridge_wasntAck <= 1'b0;
      bridge_interruptCtrl_rxDataEnable <= 1'b0;
      bridge_interruptCtrl_rxAckEnable <= 1'b0;
      bridge_interruptCtrl_txDataEnable <= 1'b0;
      bridge_interruptCtrl_txAckEnable <= 1'b0;
      bridge_interruptCtrl_start_enable <= 1'b0;
      bridge_interruptCtrl_start_flag <= 1'b0;
      bridge_interruptCtrl_restart_enable <= 1'b0;
      bridge_interruptCtrl_restart_flag <= 1'b0;
      bridge_interruptCtrl_end_enable <= 1'b0;
      bridge_interruptCtrl_end_flag <= 1'b0;
      bridge_interruptCtrl_drop_enable <= 1'b0;
      bridge_interruptCtrl_drop_flag <= 1'b0;
      bridge_interruptCtrl_filterGen_enable <= 1'b0;
      bridge_interruptCtrl_filterGen_flag <= 1'b0;
      bridge_interruptCtrl_clockGenExit_enable <= 1'b0;
      bridge_interruptCtrl_clockGenExit_flag <= 1'b0;
      bridge_interruptCtrl_clockGenEnter_enable <= 1'b0;
      bridge_interruptCtrl_clockGenEnter_flag <= 1'b0;
      _zz_io_config_samplingClockDivider <= 10'h0;
      bridge_masterLogic_fsm_stateReg <= bridge_masterLogic_fsm_enumDef_BOOT;
      bridge_slaveOverride_sda <= 1'b1;
      bridge_slaveOverride_scl <= 1'b1;
      bridge_i2cBuffer_scl_write_regNext <= 1'b1;
      bridge_i2cBuffer_sda_write_regNext <= 1'b1;
    end else begin
      if(_zz_busCtrl_rsp_ready_1) begin
        _zz_io_ctrl_rsp_valid_1 <= (busCtrl_rsp_valid && _zz_busCtrl_rsp_ready);
      end
      bridge_rxData_event <= 1'b0;
      if(when_I2cCtrl_l224) begin
        bridge_rxData_valid <= 1'b0;
      end
      if(when_I2cCtrl_l237) begin
        bridge_rxAck_valid <= 1'b0;
      end
      if(bridge_rxData_event) begin
        case(bridge_addressFilter_state)
          2'b00 : begin
            bridge_addressFilter_state <= 2'b01;
          end
          2'b01 : begin
            bridge_addressFilter_state <= 2'b10;
          end
          default : begin
          end
        endcase
      end
      if(bridge_frameReset) begin
        bridge_addressFilter_state <= 2'b00;
      end
      if(when_I2cCtrl_l310) begin
        bridge_txAck_valid <= 1'b0;
      end
      if(when_BusSlaveFactory_l377) begin
        if(when_BusSlaveFactory_l379) begin
          bridge_masterLogic_start <= _zz_bridge_masterLogic_start[0];
        end
      end
      if(when_BusSlaveFactory_l377_1) begin
        if(when_BusSlaveFactory_l379_1) begin
          bridge_masterLogic_stop <= _zz_bridge_masterLogic_stop[0];
        end
      end
      if(when_BusSlaveFactory_l377_2) begin
        if(when_BusSlaveFactory_l379_2) begin
          bridge_masterLogic_drop <= _zz_bridge_masterLogic_drop[0];
        end
      end
      if(when_BusSlaveFactory_l377_3) begin
        if(when_BusSlaveFactory_l379_3) begin
          bridge_masterLogic_recover <= _zz_bridge_masterLogic_recover[0];
        end
      end
      if(when_BusSlaveFactory_l341) begin
        if(when_BusSlaveFactory_l347) begin
          bridge_masterLogic_fsm_dropped_start <= _zz_bridge_masterLogic_fsm_dropped_start[0];
        end
      end
      if(when_BusSlaveFactory_l341_1) begin
        if(when_BusSlaveFactory_l347_1) begin
          bridge_masterLogic_fsm_dropped_stop <= _zz_bridge_masterLogic_fsm_dropped_stop[0];
        end
      end
      if(when_BusSlaveFactory_l341_2) begin
        if(when_BusSlaveFactory_l347_2) begin
          bridge_masterLogic_fsm_dropped_recover <= _zz_bridge_masterLogic_fsm_dropped_recover[0];
        end
      end
      case(i2cCtrl_io_bus_cmd_kind)
        I2cSlaveCmdMode_READ : begin
          if(when_I2cCtrl_l566) begin
            bridge_dataCounter <= (bridge_dataCounter + 3'b001);
            if(when_I2cCtrl_l570) begin
              if(bridge_txData_disableOnDataConflict) begin
                bridge_txData_enable <= 1'b0;
              end
              if(bridge_txAck_disableOnDataConflict) begin
                bridge_txAck_enable <= 1'b0;
              end
            end
            if(when_I2cCtrl_l574) begin
              if(bridge_rxData_listen) begin
                bridge_rxData_valid <= 1'b1;
              end
              bridge_rxData_event <= 1'b1;
              bridge_inAckState <= 1'b1;
              if(when_I2cCtrl_l578) begin
                bridge_txData_valid <= 1'b0;
              end
            end
          end else begin
            if(bridge_rxAck_listen) begin
              bridge_rxAck_valid <= 1'b1;
            end
            bridge_inAckState <= 1'b0;
            bridge_wasntAck <= i2cCtrl_io_bus_cmd_data;
            if(when_I2cCtrl_l588) begin
              bridge_txAck_valid <= 1'b0;
            end
          end
        end
        default : begin
        end
      endcase
      if(bridge_frameReset) begin
        bridge_inAckState <= 1'b0;
        bridge_dataCounter <= 3'b000;
        bridge_wasntAck <= 1'b0;
      end
      if(when_I2cCtrl_l601) begin
        bridge_txData_valid <= 1'b1;
        bridge_txData_enable <= 1'b0;
        bridge_txData_repeat <= 1'b1;
        bridge_txAck_valid <= 1'b1;
        bridge_txAck_enable <= 1'b0;
        bridge_txAck_repeat <= 1'b1;
        bridge_rxData_listen <= 1'b0;
        bridge_rxAck_listen <= 1'b0;
      end
      if(when_I2cCtrl_l634) begin
        bridge_interruptCtrl_start_flag <= 1'b1;
      end
      if(when_I2cCtrl_l634_1) begin
        bridge_interruptCtrl_start_flag <= 1'b0;
      end
      if(when_BusSlaveFactory_l341_3) begin
        if(when_BusSlaveFactory_l347_3) begin
          bridge_interruptCtrl_start_flag <= _zz_bridge_interruptCtrl_start_flag[0];
        end
      end
      if(when_I2cCtrl_l634_2) begin
        bridge_interruptCtrl_restart_flag <= 1'b1;
      end
      if(when_I2cCtrl_l634_3) begin
        bridge_interruptCtrl_restart_flag <= 1'b0;
      end
      if(when_BusSlaveFactory_l341_4) begin
        if(when_BusSlaveFactory_l347_4) begin
          bridge_interruptCtrl_restart_flag <= _zz_bridge_interruptCtrl_restart_flag[0];
        end
      end
      if(when_I2cCtrl_l634_4) begin
        bridge_interruptCtrl_end_flag <= 1'b1;
      end
      if(when_I2cCtrl_l634_5) begin
        bridge_interruptCtrl_end_flag <= 1'b0;
      end
      if(when_BusSlaveFactory_l341_5) begin
        if(when_BusSlaveFactory_l347_5) begin
          bridge_interruptCtrl_end_flag <= _zz_bridge_interruptCtrl_end_flag[0];
        end
      end
      if(when_I2cCtrl_l634_6) begin
        bridge_interruptCtrl_drop_flag <= 1'b1;
      end
      if(when_I2cCtrl_l634_7) begin
        bridge_interruptCtrl_drop_flag <= 1'b0;
      end
      if(when_BusSlaveFactory_l341_6) begin
        if(when_BusSlaveFactory_l347_6) begin
          bridge_interruptCtrl_drop_flag <= _zz_bridge_interruptCtrl_drop_flag[0];
        end
      end
      if(when_I2cCtrl_l634_8) begin
        bridge_interruptCtrl_filterGen_flag <= 1'b1;
      end
      if(when_I2cCtrl_l634_9) begin
        bridge_interruptCtrl_filterGen_flag <= 1'b0;
      end
      if(when_BusSlaveFactory_l341_7) begin
        if(when_BusSlaveFactory_l347_7) begin
          bridge_interruptCtrl_filterGen_flag <= _zz_bridge_interruptCtrl_filterGen_flag[0];
        end
      end
      if(when_I2cCtrl_l634_10) begin
        bridge_interruptCtrl_clockGenExit_flag <= 1'b1;
      end
      if(when_I2cCtrl_l634_11) begin
        bridge_interruptCtrl_clockGenExit_flag <= 1'b0;
      end
      if(when_BusSlaveFactory_l341_8) begin
        if(when_BusSlaveFactory_l347_8) begin
          bridge_interruptCtrl_clockGenExit_flag <= _zz_bridge_interruptCtrl_clockGenExit_flag[0];
        end
      end
      if(when_I2cCtrl_l634_12) begin
        bridge_interruptCtrl_clockGenEnter_flag <= 1'b1;
      end
      if(when_I2cCtrl_l634_13) begin
        bridge_interruptCtrl_clockGenEnter_flag <= 1'b0;
      end
      if(when_BusSlaveFactory_l341_9) begin
        if(when_BusSlaveFactory_l347_9) begin
          bridge_interruptCtrl_clockGenEnter_flag <= _zz_bridge_interruptCtrl_clockGenEnter_flag[0];
        end
      end
      bridge_masterLogic_fsm_stateReg <= bridge_masterLogic_fsm_stateNext;
      case(bridge_masterLogic_fsm_stateReg)
        bridge_masterLogic_fsm_enumDef_IDLE : begin
          if(!when_I2cCtrl_l367) begin
            if(when_I2cCtrl_l369) begin
              bridge_txData_valid <= 1'b0;
            end
          end
        end
        bridge_masterLogic_fsm_enumDef_START1 : begin
        end
        bridge_masterLogic_fsm_enumDef_START2 : begin
        end
        bridge_masterLogic_fsm_enumDef_START3 : begin
          if(bridge_masterLogic_timer_done) begin
            bridge_masterLogic_start <= 1'b0;
          end
        end
        bridge_masterLogic_fsm_enumDef_LOW : begin
        end
        bridge_masterLogic_fsm_enumDef_HIGH : begin
        end
        bridge_masterLogic_fsm_enumDef_RESTART : begin
        end
        bridge_masterLogic_fsm_enumDef_STOP1 : begin
        end
        bridge_masterLogic_fsm_enumDef_STOP2 : begin
        end
        bridge_masterLogic_fsm_enumDef_STOP3 : begin
          if(i2cCtrl_io_internals_sdaRead) begin
            bridge_masterLogic_stop <= 1'b0;
            bridge_masterLogic_recover <= 1'b0;
          end
        end
        bridge_masterLogic_fsm_enumDef_TBUF : begin
        end
        default : begin
        end
      endcase
      if(when_I2cCtrl_l350) begin
        bridge_masterLogic_start <= 1'b0;
        bridge_masterLogic_stop <= 1'b0;
        bridge_masterLogic_drop <= 1'b0;
        bridge_masterLogic_recover <= 1'b0;
        if(bridge_masterLogic_start) begin
          bridge_masterLogic_fsm_dropped_start <= 1'b1;
        end
        if(bridge_masterLogic_stop) begin
          bridge_masterLogic_fsm_dropped_stop <= 1'b1;
        end
      end
      bridge_i2cBuffer_scl_write_regNext <= bridge_i2cBuffer_scl_write;
      bridge_i2cBuffer_sda_write_regNext <= bridge_i2cBuffer_sda_write;
      case(io_ctrl_cmd_payload_fragment_address)
        8'h08 : begin
          if(busCtrl_doWrite) begin
            bridge_rxData_listen <= io_ctrl_cmd_payload_fragment_data[9];
          end
        end
        8'h0c : begin
          if(busCtrl_doWrite) begin
            bridge_rxAck_listen <= io_ctrl_cmd_payload_fragment_data[9];
          end
        end
        8'h0 : begin
          if(busCtrl_doWrite) begin
            bridge_txData_repeat <= io_ctrl_cmd_payload_fragment_data[10];
            bridge_txData_valid <= io_ctrl_cmd_payload_fragment_data[8];
            bridge_txData_enable <= io_ctrl_cmd_payload_fragment_data[9];
          end
        end
        8'h04 : begin
          if(busCtrl_doWrite) begin
            bridge_txAck_repeat <= io_ctrl_cmd_payload_fragment_data[10];
            bridge_txAck_valid <= io_ctrl_cmd_payload_fragment_data[8];
            bridge_txAck_enable <= io_ctrl_cmd_payload_fragment_data[9];
          end
        end
        8'h88 : begin
          if(busCtrl_doWrite) begin
            bridge_addressFilter_addresses_0_enable <= io_ctrl_cmd_payload_fragment_data[15];
          end
        end
        8'h8c : begin
          if(busCtrl_doWrite) begin
            bridge_addressFilter_addresses_1_enable <= io_ctrl_cmd_payload_fragment_data[15];
          end
        end
        8'h20 : begin
          if(busCtrl_doWrite) begin
            bridge_interruptCtrl_rxDataEnable <= io_ctrl_cmd_payload_fragment_data[0];
            bridge_interruptCtrl_rxAckEnable <= io_ctrl_cmd_payload_fragment_data[1];
            bridge_interruptCtrl_txDataEnable <= io_ctrl_cmd_payload_fragment_data[2];
            bridge_interruptCtrl_txAckEnable <= io_ctrl_cmd_payload_fragment_data[3];
            bridge_interruptCtrl_start_enable <= io_ctrl_cmd_payload_fragment_data[4];
            bridge_interruptCtrl_restart_enable <= io_ctrl_cmd_payload_fragment_data[5];
            bridge_interruptCtrl_end_enable <= io_ctrl_cmd_payload_fragment_data[6];
            bridge_interruptCtrl_drop_enable <= io_ctrl_cmd_payload_fragment_data[7];
            bridge_interruptCtrl_filterGen_enable <= io_ctrl_cmd_payload_fragment_data[17];
            bridge_interruptCtrl_clockGenExit_enable <= io_ctrl_cmd_payload_fragment_data[15];
            bridge_interruptCtrl_clockGenEnter_enable <= io_ctrl_cmd_payload_fragment_data[16];
          end
        end
        8'h28 : begin
          if(busCtrl_doWrite) begin
            _zz_io_config_samplingClockDivider <= io_ctrl_cmd_payload_fragment_data[9 : 0];
          end
        end
        8'h48 : begin
          if(busCtrl_doWrite) begin
            bridge_slaveOverride_sda <= io_ctrl_cmd_payload_fragment_data[1];
            bridge_slaveOverride_scl <= io_ctrl_cmd_payload_fragment_data[2];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_peripheralClk) begin
    if(_zz_busCtrl_rsp_ready_1) begin
      _zz_io_ctrl_rsp_payload_last <= busCtrl_rsp_payload_last;
      _zz_io_ctrl_rsp_payload_fragment_opcode <= busCtrl_rsp_payload_fragment_opcode;
      _zz_io_ctrl_rsp_payload_fragment_data <= busCtrl_rsp_payload_fragment_data;
      _zz_io_ctrl_rsp_payload_fragment_context <= busCtrl_rsp_payload_fragment_context;
    end
    if(bridge_rxData_event) begin
      case(bridge_addressFilter_state)
        2'b00 : begin
          bridge_addressFilter_byte0 <= bridge_rxData_value;
        end
        2'b01 : begin
          bridge_addressFilter_byte1 <= bridge_rxData_value;
        end
        default : begin
        end
      endcase
    end
    _zz_when_I2cCtrl_l310_1 <= _zz_when_I2cCtrl_l310;
    bridge_masterLogic_timer_value <= (bridge_masterLogic_timer_value - _zz_bridge_masterLogic_timer_value);
    if(when_I2cCtrl_l363) begin
      bridge_masterLogic_fsm_inFrameLate <= 1'b1;
    end
    if(when_I2cCtrl_l363_1) begin
      bridge_masterLogic_fsm_inFrameLate <= 1'b0;
    end
    case(i2cCtrl_io_bus_cmd_kind)
      I2cSlaveCmdMode_READ : begin
        if(when_I2cCtrl_l566) begin
          bridge_rxData_value[_zz_bridge_rxData_value] <= i2cCtrl_io_bus_cmd_data;
        end else begin
          bridge_rxAck_value <= i2cCtrl_io_bus_cmd_data;
        end
      end
      default : begin
      end
    endcase
    if(when_I2cCtrl_l601) begin
      bridge_txData_disableOnDataConflict <= 1'b0;
      bridge_txAck_disableOnDataConflict <= 1'b0;
    end
    _zz_when_I2cCtrl_l634_1 <= _zz_when_I2cCtrl_l634;
    bridge_masterLogic_fsm_isBusy_regNext <= bridge_masterLogic_fsm_isBusy;
    bridge_masterLogic_fsm_isBusy_regNext_1 <= bridge_masterLogic_fsm_isBusy;
    bridge_timeoutClear <= 1'b0;
    case(bridge_masterLogic_fsm_stateReg)
      bridge_masterLogic_fsm_enumDef_IDLE : begin
      end
      bridge_masterLogic_fsm_enumDef_START1 : begin
      end
      bridge_masterLogic_fsm_enumDef_START2 : begin
      end
      bridge_masterLogic_fsm_enumDef_START3 : begin
      end
      bridge_masterLogic_fsm_enumDef_LOW : begin
      end
      bridge_masterLogic_fsm_enumDef_HIGH : begin
      end
      bridge_masterLogic_fsm_enumDef_RESTART : begin
        if(when_I2cCtrl_l450) begin
          bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tHigh;
        end
      end
      bridge_masterLogic_fsm_enumDef_STOP1 : begin
      end
      bridge_masterLogic_fsm_enumDef_STOP2 : begin
        if(when_I2cCtrl_l474) begin
          bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tHigh;
        end
      end
      bridge_masterLogic_fsm_enumDef_STOP3 : begin
      end
      bridge_masterLogic_fsm_enumDef_TBUF : begin
      end
      default : begin
      end
    endcase
    if(when_StateMachine_l253) begin
      bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tHigh;
    end
    if(when_StateMachine_l253_1) begin
      bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tLow;
    end
    if(when_StateMachine_l253_2) begin
      bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tLow;
    end
    if(when_StateMachine_l253_3) begin
      bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tHigh;
    end
    if(when_StateMachine_l253_4) begin
      bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tHigh;
    end
    if(when_StateMachine_l253_5) begin
      bridge_masterLogic_timer_value <= bridge_masterLogic_timer_tBuf;
    end
    case(io_ctrl_cmd_payload_fragment_address)
      8'h0 : begin
        if(busCtrl_doWrite) begin
          bridge_txData_value <= io_ctrl_cmd_payload_fragment_data[7 : 0];
          bridge_txData_disableOnDataConflict <= io_ctrl_cmd_payload_fragment_data[11];
        end
      end
      8'h04 : begin
        if(busCtrl_doWrite) begin
          bridge_txAck_value <= io_ctrl_cmd_payload_fragment_data[0];
          bridge_txAck_disableOnDataConflict <= io_ctrl_cmd_payload_fragment_data[11];
        end
      end
      8'h88 : begin
        if(busCtrl_doWrite) begin
          bridge_addressFilter_addresses_0_value <= io_ctrl_cmd_payload_fragment_data[9 : 0];
          bridge_addressFilter_addresses_0_is10Bit <= io_ctrl_cmd_payload_fragment_data[14];
        end
      end
      8'h8c : begin
        if(busCtrl_doWrite) begin
          bridge_addressFilter_addresses_1_value <= io_ctrl_cmd_payload_fragment_data[9 : 0];
          bridge_addressFilter_addresses_1_is10Bit <= io_ctrl_cmd_payload_fragment_data[14];
        end
      end
      8'h50 : begin
        if(busCtrl_doWrite) begin
          bridge_masterLogic_timer_tLow <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      8'h54 : begin
        if(busCtrl_doWrite) begin
          bridge_masterLogic_timer_tHigh <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      8'h58 : begin
        if(busCtrl_doWrite) begin
          bridge_masterLogic_timer_tBuf <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      8'h2c : begin
        if(busCtrl_doWrite) begin
          _zz_io_config_timeout <= io_ctrl_cmd_payload_fragment_data[19 : 0];
          bridge_timeoutClear <= 1'b1;
        end
      end
      8'h30 : begin
        if(busCtrl_doWrite) begin
          _zz_io_config_tsuData <= io_ctrl_cmd_payload_fragment_data[5 : 0];
        end
      end
      default : begin
      end
    endcase
  end

  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      i2cCtrl_io_internals_inFrame_regNext <= 1'b0;
    end else begin
      i2cCtrl_io_internals_inFrame_regNext <= i2cCtrl_io_internals_inFrame;
    end
  end


endmodule

//BmbSpiXdrMasterCtrl_1 replaced by BmbSpiXdrMasterCtrl

module BmbSpiXdrMasterCtrl (
  input  wire          io_ctrl_cmd_valid,
  output wire          io_ctrl_cmd_ready,
  input  wire          io_ctrl_cmd_payload_last,
  input  wire [0:0]    io_ctrl_cmd_payload_fragment_opcode,
  input  wire [11:0]   io_ctrl_cmd_payload_fragment_address,
  input  wire [1:0]    io_ctrl_cmd_payload_fragment_length,
  input  wire [31:0]   io_ctrl_cmd_payload_fragment_data,
  input  wire [48:0]   io_ctrl_cmd_payload_fragment_context,
  output wire          io_ctrl_rsp_valid,
  input  wire          io_ctrl_rsp_ready,
  output wire          io_ctrl_rsp_payload_last,
  output wire [0:0]    io_ctrl_rsp_payload_fragment_opcode,
  output wire [31:0]   io_ctrl_rsp_payload_fragment_data,
  output wire [48:0]   io_ctrl_rsp_payload_fragment_context,
  output wire [0:0]    io_spi_sclk_write,
  output wire          io_spi_data_0_writeEnable,
  input  wire [0:0]    io_spi_data_0_read,
  output wire [0:0]    io_spi_data_0_write,
  output wire          io_spi_data_1_writeEnable,
  input  wire [0:0]    io_spi_data_1_read,
  output wire [0:0]    io_spi_data_1_write,
  output wire          io_spi_data_2_writeEnable,
  input  wire [0:0]    io_spi_data_2_read,
  output wire [0:0]    io_spi_data_2_write,
  output wire          io_spi_data_3_writeEnable,
  input  wire [0:0]    io_spi_data_3_read,
  output wire [0:0]    io_spi_data_3_write,
  output wire [0:0]    io_spi_ss,
  output wire          io_interrupt,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire                ctrl_io_rsp_queueWithOccupancy_io_pop_ready;
  wire                ctrl_io_cmd_ready;
  wire                ctrl_io_rsp_valid;
  wire       [7:0]    ctrl_io_rsp_payload_data;
  wire       [0:0]    ctrl_io_spi_sclk_write;
  wire       [0:0]    ctrl_io_spi_ss;
  wire       [0:0]    ctrl_io_spi_data_0_write;
  wire                ctrl_io_spi_data_0_writeEnable;
  wire       [0:0]    ctrl_io_spi_data_1_write;
  wire                ctrl_io_spi_data_1_writeEnable;
  wire       [0:0]    ctrl_io_spi_data_2_write;
  wire                ctrl_io_spi_data_2_writeEnable;
  wire       [0:0]    ctrl_io_spi_data_3_write;
  wire                ctrl_io_spi_data_3_writeEnable;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_push_ready;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_valid;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_kind;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_read;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_write;
  wire       [7:0]    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_data;
  wire       [8:0]    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_occupancy;
  wire       [8:0]    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_availability;
  wire                ctrl_io_rsp_queueWithOccupancy_io_push_ready;
  wire                ctrl_io_rsp_queueWithOccupancy_io_pop_valid;
  wire       [7:0]    ctrl_io_rsp_queueWithOccupancy_io_pop_payload_data;
  wire       [8:0]    ctrl_io_rsp_queueWithOccupancy_io_occupancy;
  wire       [8:0]    ctrl_io_rsp_queueWithOccupancy_io_availability;
  wire                factory_readErrorFlag;
  wire                factory_writeErrorFlag;
  wire                factory_readHaltTrigger;
  wire                factory_writeHaltTrigger;
  wire                factory_rsp_valid;
  wire                factory_rsp_ready;
  wire                factory_rsp_payload_last;
  reg        [0:0]    factory_rsp_payload_fragment_opcode;
  reg        [31:0]   factory_rsp_payload_fragment_data;
  wire       [48:0]   factory_rsp_payload_fragment_context;
  wire                _zz_factory_rsp_ready;
  reg                 _zz_factory_rsp_ready_1;
  wire                _zz_io_ctrl_rsp_valid;
  reg                 _zz_io_ctrl_rsp_valid_1;
  reg                 _zz_io_ctrl_rsp_payload_last;
  reg        [0:0]    _zz_io_ctrl_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_ctrl_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_ctrl_rsp_payload_fragment_context;
  wire                when_Stream_l375;
  wire                factory_askWrite;
  wire                factory_askRead;
  wire                io_ctrl_cmd_fire;
  wire                factory_doWrite;
  wire                factory_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  wire       [31:0]   mapping_cmdLogic_writeData;
  reg                 mapping_cmdLogic_doRegular;
  reg                 mapping_cmdLogic_doWriteLarge;
  reg                 mapping_cmdLogic_doReadWriteLarge;
  wire                mapping_cmdLogic_streamUnbuffered_valid;
  wire                mapping_cmdLogic_streamUnbuffered_ready;
  wire                mapping_cmdLogic_streamUnbuffered_payload_kind;
  wire                mapping_cmdLogic_streamUnbuffered_payload_read;
  wire                mapping_cmdLogic_streamUnbuffered_payload_write;
  wire       [7:0]    mapping_cmdLogic_streamUnbuffered_payload_data;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_valid;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_ready;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_kind;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_read;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_write;
  wire       [7:0]    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_data;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_kind;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_read;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_write;
  reg        [7:0]    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_data;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_valid;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_ready;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_kind;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_read;
  wire                mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_write;
  wire       [7:0]    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_data;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rValid;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_kind;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_read;
  reg                 mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_write;
  reg        [7:0]    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_data;
  wire                when_Stream_l375_1;
  wire                ctrl_io_rsp_toStream_valid;
  wire                ctrl_io_rsp_toStream_ready;
  wire       [7:0]    ctrl_io_rsp_toStream_payload_data;
  reg                 _zz_io_pop_ready;
  reg                 _zz_io_pop_ready_1;
  reg                 mapping_interruptCtrl_cmdIntEnable;
  reg                 mapping_interruptCtrl_rspIntEnable;
  wire                mapping_interruptCtrl_cmdInt;
  wire                mapping_interruptCtrl_rspInt;
  wire                mapping_interruptCtrl_interrupt;
  reg                 _zz_io_config_kind_cpol;
  reg                 _zz_io_config_kind_cpha;
  reg        [1:0]    _zz_io_config_mod;
  reg        [11:0]   _zz_io_config_sclkToggle;
  reg        [11:0]   _zz_io_config_ss_setup;
  reg        [11:0]   _zz_io_config_ss_hold;
  reg        [11:0]   _zz_io_config_ss_disable;
  reg        [0:0]    _zz_io_config_ss_activeHigh;
  wire       [1:0]    _zz_io_config_kind_cpol_1;

  TopLevel ctrl (
    .io_config_kind_cpol            (_zz_io_config_kind_cpol                                                                         ), //i
    .io_config_kind_cpha            (_zz_io_config_kind_cpha                                                                         ), //i
    .io_config_sclkToggle           (_zz_io_config_sclkToggle[11:0]                                                                  ), //i
    .io_config_mod                  (_zz_io_config_mod[1:0]                                                                          ), //i
    .io_config_ss_activeHigh        (_zz_io_config_ss_activeHigh                                                                     ), //i
    .io_config_ss_setup             (_zz_io_config_ss_setup[11:0]                                                                    ), //i
    .io_config_ss_hold              (_zz_io_config_ss_hold[11:0]                                                                     ), //i
    .io_config_ss_disable           (_zz_io_config_ss_disable[11:0]                                                                  ), //i
    .io_cmd_valid                   (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_valid            ), //i
    .io_cmd_ready                   (ctrl_io_cmd_ready                                                                               ), //o
    .io_cmd_payload_kind            (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_kind     ), //i
    .io_cmd_payload_read            (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_read     ), //i
    .io_cmd_payload_write           (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_write    ), //i
    .io_cmd_payload_data            (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_data[7:0]), //i
    .io_rsp_valid                   (ctrl_io_rsp_valid                                                                               ), //o
    .io_rsp_payload_data            (ctrl_io_rsp_payload_data[7:0]                                                                   ), //o
    .io_spi_sclk_write              (ctrl_io_spi_sclk_write                                                                          ), //o
    .io_spi_data_0_writeEnable      (ctrl_io_spi_data_0_writeEnable                                                                  ), //o
    .io_spi_data_0_read             (io_spi_data_0_read                                                                              ), //i
    .io_spi_data_0_write            (ctrl_io_spi_data_0_write                                                                        ), //o
    .io_spi_data_1_writeEnable      (ctrl_io_spi_data_1_writeEnable                                                                  ), //o
    .io_spi_data_1_read             (io_spi_data_1_read                                                                              ), //i
    .io_spi_data_1_write            (ctrl_io_spi_data_1_write                                                                        ), //o
    .io_spi_data_2_writeEnable      (ctrl_io_spi_data_2_writeEnable                                                                  ), //o
    .io_spi_data_2_read             (io_spi_data_2_read                                                                              ), //i
    .io_spi_data_2_write            (ctrl_io_spi_data_2_write                                                                        ), //o
    .io_spi_data_3_writeEnable      (ctrl_io_spi_data_3_writeEnable                                                                  ), //o
    .io_spi_data_3_read             (io_spi_data_3_read                                                                              ), //i
    .io_spi_data_3_write            (ctrl_io_spi_data_3_write                                                                        ), //o
    .io_spi_ss                      (ctrl_io_spi_ss                                                                                  ), //o
    .io_peripheralClk               (io_peripheralClk                                                                                ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                                                                  )  //i
  );
  StreamFifo_11 mapping_cmdLogic_streamUnbuffered_queueWithAvailability (
    .io_push_valid                  (mapping_cmdLogic_streamUnbuffered_valid                                         ), //i
    .io_push_ready                  (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_push_ready           ), //o
    .io_push_payload_kind           (mapping_cmdLogic_streamUnbuffered_payload_kind                                  ), //i
    .io_push_payload_read           (mapping_cmdLogic_streamUnbuffered_payload_read                                  ), //i
    .io_push_payload_write          (mapping_cmdLogic_streamUnbuffered_payload_write                                 ), //i
    .io_push_payload_data           (mapping_cmdLogic_streamUnbuffered_payload_data[7:0]                             ), //i
    .io_pop_valid                   (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_valid            ), //o
    .io_pop_ready                   (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN          ), //i
    .io_pop_payload_kind            (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_kind     ), //o
    .io_pop_payload_read            (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_read     ), //o
    .io_pop_payload_write           (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_write    ), //o
    .io_pop_payload_data            (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_data[7:0]), //o
    .io_flush                       (1'b0                                                                            ), //i
    .io_occupancy                   (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_occupancy[8:0]       ), //o
    .io_availability                (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_availability[8:0]    ), //o
    .io_peripheralClk               (io_peripheralClk                                                                ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                                                  )  //i
  );
  StreamFifo_12 ctrl_io_rsp_queueWithOccupancy (
    .io_push_valid                  (ctrl_io_rsp_toStream_valid                             ), //i
    .io_push_ready                  (ctrl_io_rsp_queueWithOccupancy_io_push_ready           ), //o
    .io_push_payload_data           (ctrl_io_rsp_toStream_payload_data[7:0]                 ), //i
    .io_pop_valid                   (ctrl_io_rsp_queueWithOccupancy_io_pop_valid            ), //o
    .io_pop_ready                   (ctrl_io_rsp_queueWithOccupancy_io_pop_ready            ), //i
    .io_pop_payload_data            (ctrl_io_rsp_queueWithOccupancy_io_pop_payload_data[7:0]), //o
    .io_flush                       (1'b0                                                   ), //i
    .io_occupancy                   (ctrl_io_rsp_queueWithOccupancy_io_occupancy[8:0]       ), //o
    .io_availability                (ctrl_io_rsp_queueWithOccupancy_io_availability[8:0]    ), //o
    .io_peripheralClk               (io_peripheralClk                                       ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                         )  //i
  );
  assign factory_readErrorFlag = 1'b0;
  assign factory_writeErrorFlag = 1'b0;
  assign factory_readHaltTrigger = 1'b0;
  assign factory_writeHaltTrigger = 1'b0;
  assign _zz_factory_rsp_ready = (! (factory_readHaltTrigger || factory_writeHaltTrigger));
  assign factory_rsp_ready = (_zz_factory_rsp_ready_1 && _zz_factory_rsp_ready);
  always @(*) begin
    _zz_factory_rsp_ready_1 = io_ctrl_rsp_ready;
    if(when_Stream_l375) begin
      _zz_factory_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375 = (! _zz_io_ctrl_rsp_valid);
  assign _zz_io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid_1;
  assign io_ctrl_rsp_valid = _zz_io_ctrl_rsp_valid;
  assign io_ctrl_rsp_payload_last = _zz_io_ctrl_rsp_payload_last;
  assign io_ctrl_rsp_payload_fragment_opcode = _zz_io_ctrl_rsp_payload_fragment_opcode;
  assign io_ctrl_rsp_payload_fragment_data = _zz_io_ctrl_rsp_payload_fragment_data;
  assign io_ctrl_rsp_payload_fragment_context = _zz_io_ctrl_rsp_payload_fragment_context;
  assign factory_askWrite = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign factory_askRead = (io_ctrl_cmd_valid && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign io_ctrl_cmd_fire = (io_ctrl_cmd_valid && io_ctrl_cmd_ready);
  assign factory_doWrite = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b1));
  assign factory_doRead = (io_ctrl_cmd_fire && (io_ctrl_cmd_payload_fragment_opcode == 1'b0));
  assign factory_rsp_valid = io_ctrl_cmd_valid;
  assign io_ctrl_cmd_ready = factory_rsp_ready;
  assign factory_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (factory_doWrite && factory_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      factory_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        factory_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        factory_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (factory_doRead && factory_readErrorFlag);
  always @(*) begin
    factory_rsp_payload_fragment_data = 32'h0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h0 : begin
        factory_rsp_payload_fragment_data[31 : 31] = (! ctrl_io_rsp_queueWithOccupancy_io_pop_valid);
        factory_rsp_payload_fragment_data[7 : 0] = ctrl_io_rsp_queueWithOccupancy_io_pop_payload_data;
      end
      12'h004 : begin
        factory_rsp_payload_fragment_data[8 : 0] = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_availability;
        factory_rsp_payload_fragment_data[24 : 16] = ctrl_io_rsp_queueWithOccupancy_io_occupancy;
      end
      12'h00c : begin
        factory_rsp_payload_fragment_data[16 : 16] = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_valid;
        factory_rsp_payload_fragment_data[0 : 0] = mapping_interruptCtrl_cmdIntEnable;
        factory_rsp_payload_fragment_data[1 : 1] = mapping_interruptCtrl_rspIntEnable;
        factory_rsp_payload_fragment_data[8 : 8] = mapping_interruptCtrl_cmdInt;
        factory_rsp_payload_fragment_data[9 : 9] = mapping_interruptCtrl_rspInt;
      end
      12'h058 : begin
        factory_rsp_payload_fragment_data[7 : 0] = ctrl_io_rsp_queueWithOccupancy_io_pop_payload_data;
      end
      default : begin
      end
    endcase
  end

  assign factory_rsp_payload_fragment_context = io_ctrl_cmd_payload_fragment_context;
  always @(*) begin
    mapping_cmdLogic_doRegular = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h0 : begin
        if(factory_doWrite) begin
          mapping_cmdLogic_doRegular = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mapping_cmdLogic_doWriteLarge = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h050 : begin
        if(factory_doWrite) begin
          mapping_cmdLogic_doWriteLarge = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    mapping_cmdLogic_doReadWriteLarge = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h054 : begin
        if(factory_doWrite) begin
          mapping_cmdLogic_doReadWriteLarge = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign mapping_cmdLogic_streamUnbuffered_valid = ((mapping_cmdLogic_doRegular || mapping_cmdLogic_doWriteLarge) || mapping_cmdLogic_doReadWriteLarge);
  assign mapping_cmdLogic_streamUnbuffered_payload_write = (((mapping_cmdLogic_doRegular && mapping_cmdLogic_writeData[8]) || mapping_cmdLogic_doWriteLarge) || mapping_cmdLogic_doReadWriteLarge);
  assign mapping_cmdLogic_streamUnbuffered_payload_read = ((mapping_cmdLogic_doRegular && mapping_cmdLogic_writeData[9]) || mapping_cmdLogic_doReadWriteLarge);
  assign mapping_cmdLogic_streamUnbuffered_payload_kind = (mapping_cmdLogic_doRegular && mapping_cmdLogic_writeData[11]);
  assign mapping_cmdLogic_streamUnbuffered_payload_data = mapping_cmdLogic_writeData[7:0];
  assign mapping_cmdLogic_streamUnbuffered_ready = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_push_ready;
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_valid = (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_valid || (! mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN));
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_kind = (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN ? mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_kind : mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_kind);
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_read = (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN ? mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_read : mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_read);
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_write = (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN ? mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_write : mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_write);
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_data = (mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN ? mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_data : mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_data);
  always @(*) begin
    mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_ready = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_1) begin
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_valid);
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_valid = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rValid;
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_kind = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_kind;
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_read = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_read;
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_write = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_write;
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_payload_data = mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_data;
  assign mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_m2sPipe_ready = ctrl_io_cmd_ready;
  assign ctrl_io_rsp_toStream_valid = ctrl_io_rsp_valid;
  assign ctrl_io_rsp_toStream_payload_data = ctrl_io_rsp_payload_data;
  assign ctrl_io_rsp_toStream_ready = ctrl_io_rsp_queueWithOccupancy_io_push_ready;
  always @(*) begin
    _zz_io_pop_ready = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h0 : begin
        if(factory_doRead) begin
          _zz_io_pop_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_pop_ready_1 = 1'b0;
    case(io_ctrl_cmd_payload_fragment_address)
      12'h058 : begin
        if(factory_doRead) begin
          _zz_io_pop_ready_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign ctrl_io_rsp_queueWithOccupancy_io_pop_ready = (_zz_io_pop_ready || _zz_io_pop_ready_1);
  assign mapping_interruptCtrl_cmdInt = (mapping_interruptCtrl_cmdIntEnable && (! mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_valid));
  assign mapping_interruptCtrl_rspInt = (mapping_interruptCtrl_rspIntEnable && ctrl_io_rsp_queueWithOccupancy_io_pop_valid);
  assign mapping_interruptCtrl_interrupt = (mapping_interruptCtrl_rspInt || mapping_interruptCtrl_cmdInt);
  assign io_spi_sclk_write = ctrl_io_spi_sclk_write;
  assign io_spi_data_0_writeEnable = ctrl_io_spi_data_0_writeEnable;
  assign io_spi_data_0_write = ctrl_io_spi_data_0_write;
  assign io_spi_data_1_writeEnable = ctrl_io_spi_data_1_writeEnable;
  assign io_spi_data_1_write = ctrl_io_spi_data_1_write;
  assign io_spi_data_2_writeEnable = ctrl_io_spi_data_2_writeEnable;
  assign io_spi_data_2_write = ctrl_io_spi_data_2_write;
  assign io_spi_data_3_writeEnable = ctrl_io_spi_data_3_writeEnable;
  assign io_spi_data_3_write = ctrl_io_spi_data_3_write;
  assign io_spi_ss = ctrl_io_spi_ss;
  assign io_interrupt = mapping_interruptCtrl_interrupt;
  assign mapping_cmdLogic_writeData = io_ctrl_cmd_payload_fragment_data[31 : 0];
  assign _zz_io_config_kind_cpol_1 = io_ctrl_cmd_payload_fragment_data[1 : 0];
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      _zz_io_ctrl_rsp_valid_1 <= 1'b0;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN <= 1'b1;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rValid <= 1'b0;
      mapping_interruptCtrl_cmdIntEnable <= 1'b0;
      mapping_interruptCtrl_rspIntEnable <= 1'b0;
      _zz_io_config_ss_activeHigh <= 1'b0;
    end else begin
      if(_zz_factory_rsp_ready_1) begin
        _zz_io_ctrl_rsp_valid_1 <= (factory_rsp_valid && _zz_factory_rsp_ready);
      end
      if(mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_valid) begin
        mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN <= 1'b0;
      end
      if(mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_ready) begin
        mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN <= 1'b1;
      end
      if(mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_ready) begin
        mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rValid <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_valid;
      end
      case(io_ctrl_cmd_payload_fragment_address)
        12'h00c : begin
          if(factory_doWrite) begin
            mapping_interruptCtrl_cmdIntEnable <= io_ctrl_cmd_payload_fragment_data[0];
            mapping_interruptCtrl_rspIntEnable <= io_ctrl_cmd_payload_fragment_data[1];
          end
        end
        12'h030 : begin
          if(factory_doWrite) begin
            _zz_io_config_ss_activeHigh <= io_ctrl_cmd_payload_fragment_data[0 : 0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_peripheralClk) begin
    if(_zz_factory_rsp_ready_1) begin
      _zz_io_ctrl_rsp_payload_last <= factory_rsp_payload_last;
      _zz_io_ctrl_rsp_payload_fragment_opcode <= factory_rsp_payload_fragment_opcode;
      _zz_io_ctrl_rsp_payload_fragment_data <= factory_rsp_payload_fragment_data;
      _zz_io_ctrl_rsp_payload_fragment_context <= factory_rsp_payload_fragment_context;
    end
    if(mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rValidN) begin
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_kind <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_kind;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_read <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_read;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_write <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_write;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_rData_data <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_payload_data;
    end
    if(mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_ready) begin
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_kind <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_kind;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_read <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_read;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_write <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_write;
      mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_rData_data <= mapping_cmdLogic_streamUnbuffered_queueWithAvailability_io_pop_s2mPipe_payload_data;
    end
    case(io_ctrl_cmd_payload_fragment_address)
      12'h008 : begin
        if(factory_doWrite) begin
          _zz_io_config_kind_cpol <= _zz_io_config_kind_cpol_1[0];
          _zz_io_config_kind_cpha <= _zz_io_config_kind_cpol_1[1];
          _zz_io_config_mod <= io_ctrl_cmd_payload_fragment_data[5 : 4];
        end
      end
      12'h020 : begin
        if(factory_doWrite) begin
          _zz_io_config_sclkToggle <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      12'h024 : begin
        if(factory_doWrite) begin
          _zz_io_config_ss_setup <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      12'h028 : begin
        if(factory_doWrite) begin
          _zz_io_config_ss_hold <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      12'h02c : begin
        if(factory_doWrite) begin
          _zz_io_config_ss_disable <= io_ctrl_cmd_payload_fragment_data[11 : 0];
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module BmbUartCtrl (
  input  wire          io_bus_cmd_valid,
  output wire          io_bus_cmd_ready,
  input  wire          io_bus_cmd_payload_last,
  input  wire [0:0]    io_bus_cmd_payload_fragment_opcode,
  input  wire [5:0]    io_bus_cmd_payload_fragment_address,
  input  wire [1:0]    io_bus_cmd_payload_fragment_length,
  input  wire [31:0]   io_bus_cmd_payload_fragment_data,
  input  wire [48:0]   io_bus_cmd_payload_fragment_context,
  output wire          io_bus_rsp_valid,
  input  wire          io_bus_rsp_ready,
  output wire          io_bus_rsp_payload_last,
  output wire [0:0]    io_bus_rsp_payload_fragment_opcode,
  output wire [31:0]   io_bus_rsp_payload_fragment_data,
  output wire [48:0]   io_bus_rsp_payload_fragment_context,
  output wire          io_uart_txd,
  input  wire          io_uart_rxd,
  output wire          io_interrupt,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;

  reg                 uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready;
  wire                uartCtrl_1_io_write_ready;
  wire                uartCtrl_1_io_read_valid;
  wire       [7:0]    uartCtrl_1_io_read_payload;
  wire                uartCtrl_1_io_uart_txd;
  wire                uartCtrl_1_io_readError;
  wire                uartCtrl_1_io_readBreak;
  wire                bridge_write_streamUnbuffered_queueWithOccupancy_io_push_ready;
  wire                bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid;
  wire       [7:0]    bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_payload;
  wire       [7:0]    bridge_write_streamUnbuffered_queueWithOccupancy_io_occupancy;
  wire       [7:0]    bridge_write_streamUnbuffered_queueWithOccupancy_io_availability;
  wire                uartCtrl_1_io_read_queueWithOccupancy_io_push_ready;
  wire                uartCtrl_1_io_read_queueWithOccupancy_io_pop_valid;
  wire       [7:0]    uartCtrl_1_io_read_queueWithOccupancy_io_pop_payload;
  wire       [7:0]    uartCtrl_1_io_read_queueWithOccupancy_io_occupancy;
  wire       [7:0]    uartCtrl_1_io_read_queueWithOccupancy_io_availability;
  wire       [0:0]    _zz_bridge_misc_readError;
  wire       [0:0]    _zz_bridge_misc_readOverflowError;
  wire       [0:0]    _zz_bridge_misc_breakDetected;
  wire       [0:0]    _zz_bridge_misc_doBreak;
  wire       [0:0]    _zz_bridge_misc_doBreak_1;
  wire       [7:0]    _zz_busCtrl_rsp_payload_fragment_data;
  wire                busCtrl_readErrorFlag;
  wire                busCtrl_writeErrorFlag;
  wire                busCtrl_readHaltTrigger;
  wire                busCtrl_writeHaltTrigger;
  wire                busCtrl_rsp_valid;
  wire                busCtrl_rsp_ready;
  wire                busCtrl_rsp_payload_last;
  reg        [0:0]    busCtrl_rsp_payload_fragment_opcode;
  reg        [31:0]   busCtrl_rsp_payload_fragment_data;
  wire       [48:0]   busCtrl_rsp_payload_fragment_context;
  wire                _zz_busCtrl_rsp_ready;
  reg                 _zz_busCtrl_rsp_ready_1;
  wire                _zz_io_bus_rsp_valid;
  reg                 _zz_io_bus_rsp_valid_1;
  reg                 _zz_io_bus_rsp_payload_last;
  reg        [0:0]    _zz_io_bus_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_bus_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_bus_rsp_payload_fragment_context;
  wire                when_Stream_l375;
  wire                busCtrl_askWrite;
  wire                busCtrl_askRead;
  wire                io_bus_cmd_fire;
  wire                busCtrl_doWrite;
  wire                busCtrl_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  wire                bridge_busCtrlWrapped_readErrorFlag;
  wire                bridge_busCtrlWrapped_writeErrorFlag;
  reg        [2:0]    bridge_uartConfigReg_frame_dataLength;
  reg        [0:0]    bridge_uartConfigReg_frame_stop;
  reg        [1:0]    bridge_uartConfigReg_frame_parity;
  reg        [19:0]   bridge_uartConfigReg_clockDivider;
  reg                 _zz_bridge_write_streamUnbuffered_valid;
  wire                bridge_write_streamUnbuffered_valid;
  wire                bridge_write_streamUnbuffered_ready;
  wire       [7:0]    bridge_write_streamUnbuffered_payload;
  reg                 bridge_read_streamBreaked_valid;
  reg                 bridge_read_streamBreaked_ready;
  wire       [7:0]    bridge_read_streamBreaked_payload;
  reg                 bridge_interruptCtrl_writeIntEnable;
  reg                 bridge_interruptCtrl_readIntEnable;
  wire                bridge_interruptCtrl_readInt;
  wire                bridge_interruptCtrl_writeInt;
  wire                bridge_interruptCtrl_interrupt;
  reg                 bridge_misc_readError;
  reg                 when_BusSlaveFactory_l341;
  wire                when_BusSlaveFactory_l347;
  reg                 bridge_misc_readOverflowError;
  reg                 when_BusSlaveFactory_l341_1;
  wire                when_BusSlaveFactory_l347_1;
  wire                uartCtrl_1_io_read_isStall;
  reg                 bridge_misc_breakDetected;
  reg                 uartCtrl_1_io_readBreak_regNext;
  wire                when_UartCtrl_l155;
  reg                 when_BusSlaveFactory_l341_2;
  wire                when_BusSlaveFactory_l347_2;
  reg                 bridge_misc_doBreak;
  reg                 when_BusSlaveFactory_l377;
  wire                when_BusSlaveFactory_l379;
  reg                 when_BusSlaveFactory_l341_3;
  wire                when_BusSlaveFactory_l347_3;
  wire       [1:0]    _zz_bridge_uartConfigReg_frame_parity;
  wire       [0:0]    _zz_bridge_uartConfigReg_frame_stop;
  wire                when_BmbSlaveFactory_l77;
  `ifndef SYNTHESIS
  reg [23:0] bridge_uartConfigReg_frame_stop_string;
  reg [31:0] bridge_uartConfigReg_frame_parity_string;
  reg [31:0] _zz_bridge_uartConfigReg_frame_parity_string;
  reg [23:0] _zz_bridge_uartConfigReg_frame_stop_string;
  `endif


  assign _zz_bridge_misc_readError = 1'b0;
  assign _zz_bridge_misc_readOverflowError = 1'b0;
  assign _zz_bridge_misc_breakDetected = 1'b0;
  assign _zz_bridge_misc_doBreak = 1'b1;
  assign _zz_bridge_misc_doBreak_1 = 1'b0;
  assign _zz_busCtrl_rsp_payload_fragment_data = (8'h80 - bridge_write_streamUnbuffered_queueWithOccupancy_io_occupancy);
  UartCtrl uartCtrl_1 (
    .io_config_frame_dataLength     (bridge_uartConfigReg_frame_dataLength[2:0]                          ), //i
    .io_config_frame_stop           (bridge_uartConfigReg_frame_stop                                     ), //i
    .io_config_frame_parity         (bridge_uartConfigReg_frame_parity[1:0]                              ), //i
    .io_config_clockDivider         (bridge_uartConfigReg_clockDivider[19:0]                             ), //i
    .io_write_valid                 (bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid       ), //i
    .io_write_ready                 (uartCtrl_1_io_write_ready                                           ), //o
    .io_write_payload               (bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_payload[7:0]), //i
    .io_read_valid                  (uartCtrl_1_io_read_valid                                            ), //o
    .io_read_ready                  (uartCtrl_1_io_read_queueWithOccupancy_io_push_ready                 ), //i
    .io_read_payload                (uartCtrl_1_io_read_payload[7:0]                                     ), //o
    .io_uart_txd                    (uartCtrl_1_io_uart_txd                                              ), //o
    .io_uart_rxd                    (io_uart_rxd                                                         ), //i
    .io_readError                   (uartCtrl_1_io_readError                                             ), //o
    .io_writeBreak                  (bridge_misc_doBreak                                                 ), //i
    .io_readBreak                   (uartCtrl_1_io_readBreak                                             ), //o
    .io_peripheralClk               (io_peripheralClk                                                    ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                                      )  //i
  );
  StreamFifo_9 bridge_write_streamUnbuffered_queueWithOccupancy (
    .io_push_valid                  (bridge_write_streamUnbuffered_valid                                  ), //i
    .io_push_ready                  (bridge_write_streamUnbuffered_queueWithOccupancy_io_push_ready       ), //o
    .io_push_payload                (bridge_write_streamUnbuffered_payload[7:0]                           ), //i
    .io_pop_valid                   (bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid        ), //o
    .io_pop_ready                   (uartCtrl_1_io_write_ready                                            ), //i
    .io_pop_payload                 (bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_payload[7:0] ), //o
    .io_flush                       (1'b0                                                                 ), //i
    .io_occupancy                   (bridge_write_streamUnbuffered_queueWithOccupancy_io_occupancy[7:0]   ), //o
    .io_availability                (bridge_write_streamUnbuffered_queueWithOccupancy_io_availability[7:0]), //o
    .io_peripheralClk               (io_peripheralClk                                                     ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                                       )  //i
  );
  StreamFifo_9 uartCtrl_1_io_read_queueWithOccupancy (
    .io_push_valid                  (uartCtrl_1_io_read_valid                                  ), //i
    .io_push_ready                  (uartCtrl_1_io_read_queueWithOccupancy_io_push_ready       ), //o
    .io_push_payload                (uartCtrl_1_io_read_payload[7:0]                           ), //i
    .io_pop_valid                   (uartCtrl_1_io_read_queueWithOccupancy_io_pop_valid        ), //o
    .io_pop_ready                   (uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready        ), //i
    .io_pop_payload                 (uartCtrl_1_io_read_queueWithOccupancy_io_pop_payload[7:0] ), //o
    .io_flush                       (1'b0                                                      ), //i
    .io_occupancy                   (uartCtrl_1_io_read_queueWithOccupancy_io_occupancy[7:0]   ), //o
    .io_availability                (uartCtrl_1_io_read_queueWithOccupancy_io_availability[7:0]), //o
    .io_peripheralClk               (io_peripheralClk                                          ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                            )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(bridge_uartConfigReg_frame_stop)
      UartStopType_ONE : bridge_uartConfigReg_frame_stop_string = "ONE";
      UartStopType_TWO : bridge_uartConfigReg_frame_stop_string = "TWO";
      default : bridge_uartConfigReg_frame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(bridge_uartConfigReg_frame_parity)
      UartParityType_NONE : bridge_uartConfigReg_frame_parity_string = "NONE";
      UartParityType_EVEN : bridge_uartConfigReg_frame_parity_string = "EVEN";
      UartParityType_ODD : bridge_uartConfigReg_frame_parity_string = "ODD ";
      default : bridge_uartConfigReg_frame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_bridge_uartConfigReg_frame_parity)
      UartParityType_NONE : _zz_bridge_uartConfigReg_frame_parity_string = "NONE";
      UartParityType_EVEN : _zz_bridge_uartConfigReg_frame_parity_string = "EVEN";
      UartParityType_ODD : _zz_bridge_uartConfigReg_frame_parity_string = "ODD ";
      default : _zz_bridge_uartConfigReg_frame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_bridge_uartConfigReg_frame_stop)
      UartStopType_ONE : _zz_bridge_uartConfigReg_frame_stop_string = "ONE";
      UartStopType_TWO : _zz_bridge_uartConfigReg_frame_stop_string = "TWO";
      default : _zz_bridge_uartConfigReg_frame_stop_string = "???";
    endcase
  end
  `endif

  assign io_uart_txd = uartCtrl_1_io_uart_txd;
  assign busCtrl_readErrorFlag = 1'b0;
  assign busCtrl_writeErrorFlag = 1'b0;
  assign busCtrl_readHaltTrigger = 1'b0;
  assign busCtrl_writeHaltTrigger = 1'b0;
  assign _zz_busCtrl_rsp_ready = (! (busCtrl_readHaltTrigger || busCtrl_writeHaltTrigger));
  assign busCtrl_rsp_ready = (_zz_busCtrl_rsp_ready_1 && _zz_busCtrl_rsp_ready);
  always @(*) begin
    _zz_busCtrl_rsp_ready_1 = io_bus_rsp_ready;
    if(when_Stream_l375) begin
      _zz_busCtrl_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375 = (! _zz_io_bus_rsp_valid);
  assign _zz_io_bus_rsp_valid = _zz_io_bus_rsp_valid_1;
  assign io_bus_rsp_valid = _zz_io_bus_rsp_valid;
  assign io_bus_rsp_payload_last = _zz_io_bus_rsp_payload_last;
  assign io_bus_rsp_payload_fragment_opcode = _zz_io_bus_rsp_payload_fragment_opcode;
  assign io_bus_rsp_payload_fragment_data = _zz_io_bus_rsp_payload_fragment_data;
  assign io_bus_rsp_payload_fragment_context = _zz_io_bus_rsp_payload_fragment_context;
  assign busCtrl_askWrite = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_askRead = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign io_bus_cmd_fire = (io_bus_cmd_valid && io_bus_cmd_ready);
  assign busCtrl_doWrite = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign busCtrl_doRead = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign busCtrl_rsp_valid = io_bus_cmd_valid;
  assign io_bus_cmd_ready = busCtrl_rsp_ready;
  assign busCtrl_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (busCtrl_doWrite && busCtrl_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      busCtrl_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        busCtrl_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        busCtrl_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (busCtrl_doRead && busCtrl_readErrorFlag);
  always @(*) begin
    busCtrl_rsp_payload_fragment_data = 32'h0;
    case(io_bus_cmd_payload_fragment_address)
      6'h0 : begin
        busCtrl_rsp_payload_fragment_data[16 : 16] = (bridge_read_streamBreaked_valid ^ 1'b0);
        busCtrl_rsp_payload_fragment_data[7 : 0] = bridge_read_streamBreaked_payload;
      end
      6'h04 : begin
        busCtrl_rsp_payload_fragment_data[23 : 16] = _zz_busCtrl_rsp_payload_fragment_data;
        busCtrl_rsp_payload_fragment_data[15 : 15] = bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid;
        busCtrl_rsp_payload_fragment_data[31 : 24] = uartCtrl_1_io_read_queueWithOccupancy_io_occupancy;
        busCtrl_rsp_payload_fragment_data[0 : 0] = bridge_interruptCtrl_writeIntEnable;
        busCtrl_rsp_payload_fragment_data[1 : 1] = bridge_interruptCtrl_readIntEnable;
        busCtrl_rsp_payload_fragment_data[8 : 8] = bridge_interruptCtrl_writeInt;
        busCtrl_rsp_payload_fragment_data[9 : 9] = bridge_interruptCtrl_readInt;
      end
      6'h10 : begin
        busCtrl_rsp_payload_fragment_data[0 : 0] = bridge_misc_readError;
        busCtrl_rsp_payload_fragment_data[1 : 1] = bridge_misc_readOverflowError;
        busCtrl_rsp_payload_fragment_data[8 : 8] = uartCtrl_1_io_readBreak;
        busCtrl_rsp_payload_fragment_data[9 : 9] = bridge_misc_breakDetected;
      end
      default : begin
      end
    endcase
  end

  assign busCtrl_rsp_payload_fragment_context = io_bus_cmd_payload_fragment_context;
  assign bridge_busCtrlWrapped_readErrorFlag = 1'b0;
  assign bridge_busCtrlWrapped_writeErrorFlag = 1'b0;
  always @(*) begin
    _zz_bridge_write_streamUnbuffered_valid = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      6'h0 : begin
        if(busCtrl_doWrite) begin
          _zz_bridge_write_streamUnbuffered_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign bridge_write_streamUnbuffered_valid = _zz_bridge_write_streamUnbuffered_valid;
  assign bridge_write_streamUnbuffered_payload = io_bus_cmd_payload_fragment_data[7 : 0];
  assign bridge_write_streamUnbuffered_ready = bridge_write_streamUnbuffered_queueWithOccupancy_io_push_ready;
  always @(*) begin
    bridge_read_streamBreaked_valid = uartCtrl_1_io_read_queueWithOccupancy_io_pop_valid;
    if(uartCtrl_1_io_readBreak) begin
      bridge_read_streamBreaked_valid = 1'b0;
    end
  end

  always @(*) begin
    uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready = bridge_read_streamBreaked_ready;
    if(uartCtrl_1_io_readBreak) begin
      uartCtrl_1_io_read_queueWithOccupancy_io_pop_ready = 1'b1;
    end
  end

  assign bridge_read_streamBreaked_payload = uartCtrl_1_io_read_queueWithOccupancy_io_pop_payload;
  always @(*) begin
    bridge_read_streamBreaked_ready = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      6'h0 : begin
        if(busCtrl_doRead) begin
          bridge_read_streamBreaked_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign bridge_interruptCtrl_readInt = (bridge_interruptCtrl_readIntEnable && bridge_read_streamBreaked_valid);
  assign bridge_interruptCtrl_writeInt = (bridge_interruptCtrl_writeIntEnable && (! bridge_write_streamUnbuffered_queueWithOccupancy_io_pop_valid));
  assign bridge_interruptCtrl_interrupt = (bridge_interruptCtrl_readInt || bridge_interruptCtrl_writeInt);
  always @(*) begin
    when_BusSlaveFactory_l341 = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      6'h10 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347 = io_bus_cmd_payload_fragment_data[0];
  always @(*) begin
    when_BusSlaveFactory_l341_1 = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      6'h10 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_1 = io_bus_cmd_payload_fragment_data[1];
  assign uartCtrl_1_io_read_isStall = (uartCtrl_1_io_read_valid && (! uartCtrl_1_io_read_queueWithOccupancy_io_push_ready));
  assign when_UartCtrl_l155 = (uartCtrl_1_io_readBreak && (! uartCtrl_1_io_readBreak_regNext));
  always @(*) begin
    when_BusSlaveFactory_l341_2 = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      6'h10 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_2 = io_bus_cmd_payload_fragment_data[9];
  always @(*) begin
    when_BusSlaveFactory_l377 = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      6'h10 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l377 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379 = io_bus_cmd_payload_fragment_data[10];
  always @(*) begin
    when_BusSlaveFactory_l341_3 = 1'b0;
    case(io_bus_cmd_payload_fragment_address)
      6'h10 : begin
        if(busCtrl_doWrite) begin
          when_BusSlaveFactory_l341_3 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l347_3 = io_bus_cmd_payload_fragment_data[11];
  assign io_interrupt = bridge_interruptCtrl_interrupt;
  assign _zz_bridge_uartConfigReg_frame_parity = io_bus_cmd_payload_fragment_data[9 : 8];
  assign _zz_bridge_uartConfigReg_frame_stop = io_bus_cmd_payload_fragment_data[16 : 16];
  assign when_BmbSlaveFactory_l77 = ((io_bus_cmd_payload_fragment_address & (~ 6'h03)) == 6'h08);
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      _zz_io_bus_rsp_valid_1 <= 1'b0;
      bridge_uartConfigReg_clockDivider <= 20'h0;
      bridge_uartConfigReg_clockDivider <= 20'h00035;
      bridge_uartConfigReg_frame_dataLength <= 3'b111;
      bridge_uartConfigReg_frame_parity <= UartParityType_NONE;
      bridge_uartConfigReg_frame_stop <= UartStopType_ONE;
      bridge_interruptCtrl_writeIntEnable <= 1'b0;
      bridge_interruptCtrl_readIntEnable <= 1'b0;
      bridge_misc_readError <= 1'b0;
      bridge_misc_readOverflowError <= 1'b0;
      bridge_misc_breakDetected <= 1'b0;
      bridge_misc_doBreak <= 1'b0;
    end else begin
      if(_zz_busCtrl_rsp_ready_1) begin
        _zz_io_bus_rsp_valid_1 <= (busCtrl_rsp_valid && _zz_busCtrl_rsp_ready);
      end
      if(when_BusSlaveFactory_l341) begin
        if(when_BusSlaveFactory_l347) begin
          bridge_misc_readError <= _zz_bridge_misc_readError[0];
        end
      end
      if(uartCtrl_1_io_readError) begin
        bridge_misc_readError <= 1'b1;
      end
      if(when_BusSlaveFactory_l341_1) begin
        if(when_BusSlaveFactory_l347_1) begin
          bridge_misc_readOverflowError <= _zz_bridge_misc_readOverflowError[0];
        end
      end
      if(uartCtrl_1_io_read_isStall) begin
        bridge_misc_readOverflowError <= 1'b1;
      end
      if(when_UartCtrl_l155) begin
        bridge_misc_breakDetected <= 1'b1;
      end
      if(when_BusSlaveFactory_l341_2) begin
        if(when_BusSlaveFactory_l347_2) begin
          bridge_misc_breakDetected <= _zz_bridge_misc_breakDetected[0];
        end
      end
      if(when_BusSlaveFactory_l377) begin
        if(when_BusSlaveFactory_l379) begin
          bridge_misc_doBreak <= _zz_bridge_misc_doBreak[0];
        end
      end
      if(when_BusSlaveFactory_l341_3) begin
        if(when_BusSlaveFactory_l347_3) begin
          bridge_misc_doBreak <= _zz_bridge_misc_doBreak_1[0];
        end
      end
      case(io_bus_cmd_payload_fragment_address)
        6'h0c : begin
          if(busCtrl_doWrite) begin
            bridge_uartConfigReg_frame_dataLength <= io_bus_cmd_payload_fragment_data[2 : 0];
            bridge_uartConfigReg_frame_parity <= _zz_bridge_uartConfigReg_frame_parity;
            bridge_uartConfigReg_frame_stop <= _zz_bridge_uartConfigReg_frame_stop;
          end
        end
        6'h04 : begin
          if(busCtrl_doWrite) begin
            bridge_interruptCtrl_writeIntEnable <= io_bus_cmd_payload_fragment_data[0];
            bridge_interruptCtrl_readIntEnable <= io_bus_cmd_payload_fragment_data[1];
          end
        end
        default : begin
        end
      endcase
      if(when_BmbSlaveFactory_l77) begin
        if(busCtrl_doWrite) begin
          bridge_uartConfigReg_clockDivider[19 : 0] <= io_bus_cmd_payload_fragment_data[19 : 0];
        end
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(_zz_busCtrl_rsp_ready_1) begin
      _zz_io_bus_rsp_payload_last <= busCtrl_rsp_payload_last;
      _zz_io_bus_rsp_payload_fragment_opcode <= busCtrl_rsp_payload_fragment_opcode;
      _zz_io_bus_rsp_payload_fragment_data <= busCtrl_rsp_payload_fragment_data;
      _zz_io_bus_rsp_payload_fragment_context <= busCtrl_rsp_payload_fragment_context;
    end
    uartCtrl_1_io_readBreak_regNext <= uartCtrl_1_io_readBreak;
  end


endmodule

module BmbClint (
  input  wire          io_bus_cmd_valid,
  output wire          io_bus_cmd_ready,
  input  wire          io_bus_cmd_payload_last,
  input  wire [0:0]    io_bus_cmd_payload_fragment_opcode,
  input  wire [15:0]   io_bus_cmd_payload_fragment_address,
  input  wire [1:0]    io_bus_cmd_payload_fragment_length,
  input  wire [31:0]   io_bus_cmd_payload_fragment_data,
  input  wire [48:0]   io_bus_cmd_payload_fragment_context,
  output wire          io_bus_rsp_valid,
  input  wire          io_bus_rsp_ready,
  output wire          io_bus_rsp_payload_last,
  output wire [0:0]    io_bus_rsp_payload_fragment_opcode,
  output wire [31:0]   io_bus_rsp_payload_fragment_data,
  output wire [48:0]   io_bus_rsp_payload_fragment_context,
  output reg  [1:0]    io_timerInterrupt,
  output reg  [1:0]    io_softwareInterrupt,
  output wire [63:0]   io_time,
  input  wire          io_stop,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire                factory_readErrorFlag;
  wire                factory_writeErrorFlag;
  wire                factory_readHaltTrigger;
  wire                factory_writeHaltTrigger;
  wire                factory_rsp_valid;
  wire                factory_rsp_ready;
  wire                factory_rsp_payload_last;
  reg        [0:0]    factory_rsp_payload_fragment_opcode;
  reg        [31:0]   factory_rsp_payload_fragment_data;
  wire       [48:0]   factory_rsp_payload_fragment_context;
  wire                _zz_factory_rsp_ready;
  reg                 _zz_factory_rsp_ready_1;
  wire                _zz_io_bus_rsp_valid;
  reg                 _zz_io_bus_rsp_valid_1;
  reg                 _zz_io_bus_rsp_payload_last;
  reg        [0:0]    _zz_io_bus_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_bus_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_bus_rsp_payload_fragment_context;
  wire                when_Stream_l375;
  wire                factory_askWrite;
  wire                factory_askRead;
  wire                io_bus_cmd_fire;
  wire                factory_doWrite;
  wire                factory_doRead;
  wire                when_BmbSlaveFactory_l33;
  wire                when_BmbSlaveFactory_l35;
  reg                 logic_stop;
  reg        [63:0]   logic_time;
  wire                when_Clint_l39;
  reg        [63:0]   logic_harts_0_cmp;
  reg                 logic_harts_0_timerInterrupt;
  reg                 logic_harts_0_softwareInterrupt;
  reg        [63:0]   logic_harts_1_cmp;
  reg                 logic_harts_1_timerInterrupt;
  reg                 logic_harts_1_softwareInterrupt;
  wire       [63:0]   _zz_factory_rsp_payload_fragment_data;
  wire                when_BmbSlaveFactory_l77;
  wire                when_BmbSlaveFactory_l77_1;
  wire                when_BmbSlaveFactory_l77_2;
  wire                when_BmbSlaveFactory_l77_3;
  wire                when_BmbSlaveFactory_l77_4;
  wire                when_BmbSlaveFactory_l77_5;

  assign factory_readErrorFlag = 1'b0;
  assign factory_writeErrorFlag = 1'b0;
  assign factory_readHaltTrigger = 1'b0;
  assign factory_writeHaltTrigger = 1'b0;
  assign _zz_factory_rsp_ready = (! (factory_readHaltTrigger || factory_writeHaltTrigger));
  assign factory_rsp_ready = (_zz_factory_rsp_ready_1 && _zz_factory_rsp_ready);
  always @(*) begin
    _zz_factory_rsp_ready_1 = io_bus_rsp_ready;
    if(when_Stream_l375) begin
      _zz_factory_rsp_ready_1 = 1'b1;
    end
  end

  assign when_Stream_l375 = (! _zz_io_bus_rsp_valid);
  assign _zz_io_bus_rsp_valid = _zz_io_bus_rsp_valid_1;
  assign io_bus_rsp_valid = _zz_io_bus_rsp_valid;
  assign io_bus_rsp_payload_last = _zz_io_bus_rsp_payload_last;
  assign io_bus_rsp_payload_fragment_opcode = _zz_io_bus_rsp_payload_fragment_opcode;
  assign io_bus_rsp_payload_fragment_data = _zz_io_bus_rsp_payload_fragment_data;
  assign io_bus_rsp_payload_fragment_context = _zz_io_bus_rsp_payload_fragment_context;
  assign factory_askWrite = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign factory_askRead = (io_bus_cmd_valid && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign io_bus_cmd_fire = (io_bus_cmd_valid && io_bus_cmd_ready);
  assign factory_doWrite = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b1));
  assign factory_doRead = (io_bus_cmd_fire && (io_bus_cmd_payload_fragment_opcode == 1'b0));
  assign factory_rsp_valid = io_bus_cmd_valid;
  assign io_bus_cmd_ready = factory_rsp_ready;
  assign factory_rsp_payload_last = 1'b1;
  assign when_BmbSlaveFactory_l33 = (factory_doWrite && factory_writeErrorFlag);
  always @(*) begin
    if(when_BmbSlaveFactory_l33) begin
      factory_rsp_payload_fragment_opcode = 1'b1;
    end else begin
      if(when_BmbSlaveFactory_l35) begin
        factory_rsp_payload_fragment_opcode = 1'b1;
      end else begin
        factory_rsp_payload_fragment_opcode = 1'b0;
      end
    end
  end

  assign when_BmbSlaveFactory_l35 = (factory_doRead && factory_readErrorFlag);
  always @(*) begin
    factory_rsp_payload_fragment_data = 32'h0;
    case(io_bus_cmd_payload_fragment_address)
      16'h0 : begin
        factory_rsp_payload_fragment_data[0 : 0] = logic_harts_0_softwareInterrupt;
      end
      16'h0004 : begin
        factory_rsp_payload_fragment_data[0 : 0] = logic_harts_1_softwareInterrupt;
      end
      default : begin
      end
    endcase
    if(when_BmbSlaveFactory_l77) begin
      factory_rsp_payload_fragment_data[31 : 0] = _zz_factory_rsp_payload_fragment_data[31 : 0];
    end
    if(when_BmbSlaveFactory_l77_1) begin
      factory_rsp_payload_fragment_data[31 : 0] = _zz_factory_rsp_payload_fragment_data[63 : 32];
    end
  end

  assign factory_rsp_payload_fragment_context = io_bus_cmd_payload_fragment_context;
  always @(*) begin
    logic_stop = 1'b0;
    if(io_stop) begin
      logic_stop = 1'b1;
    end
  end

  assign when_Clint_l39 = (! logic_stop);
  assign _zz_factory_rsp_payload_fragment_data = logic_time;
  always @(*) begin
    io_timerInterrupt[0] = logic_harts_0_timerInterrupt;
    io_timerInterrupt[1] = logic_harts_1_timerInterrupt;
  end

  always @(*) begin
    io_softwareInterrupt[0] = logic_harts_0_softwareInterrupt;
    io_softwareInterrupt[1] = logic_harts_1_softwareInterrupt;
  end

  assign io_time = logic_time;
  assign when_BmbSlaveFactory_l77 = ((io_bus_cmd_payload_fragment_address & (~ 16'h0003)) == 16'hbff8);
  assign when_BmbSlaveFactory_l77_1 = ((io_bus_cmd_payload_fragment_address & (~ 16'h0003)) == 16'hbffc);
  assign when_BmbSlaveFactory_l77_2 = ((io_bus_cmd_payload_fragment_address & (~ 16'h0003)) == 16'h4000);
  assign when_BmbSlaveFactory_l77_3 = ((io_bus_cmd_payload_fragment_address & (~ 16'h0003)) == 16'h4004);
  assign when_BmbSlaveFactory_l77_4 = ((io_bus_cmd_payload_fragment_address & (~ 16'h0003)) == 16'h4008);
  assign when_BmbSlaveFactory_l77_5 = ((io_bus_cmd_payload_fragment_address & (~ 16'h0003)) == 16'h400c);
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      _zz_io_bus_rsp_valid_1 <= 1'b0;
      logic_time <= 64'h0;
      logic_harts_0_softwareInterrupt <= 1'b0;
      logic_harts_1_softwareInterrupt <= 1'b0;
    end else begin
      if(_zz_factory_rsp_ready_1) begin
        _zz_io_bus_rsp_valid_1 <= (factory_rsp_valid && _zz_factory_rsp_ready);
      end
      if(when_Clint_l39) begin
        logic_time <= (logic_time + 64'h0000000000000001);
      end
      case(io_bus_cmd_payload_fragment_address)
        16'h0 : begin
          if(factory_doWrite) begin
            logic_harts_0_softwareInterrupt <= io_bus_cmd_payload_fragment_data[0];
          end
        end
        16'h0004 : begin
          if(factory_doWrite) begin
            logic_harts_1_softwareInterrupt <= io_bus_cmd_payload_fragment_data[0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_peripheralClk) begin
    if(_zz_factory_rsp_ready_1) begin
      _zz_io_bus_rsp_payload_last <= factory_rsp_payload_last;
      _zz_io_bus_rsp_payload_fragment_opcode <= factory_rsp_payload_fragment_opcode;
      _zz_io_bus_rsp_payload_fragment_data <= factory_rsp_payload_fragment_data;
      _zz_io_bus_rsp_payload_fragment_context <= factory_rsp_payload_fragment_context;
    end
    logic_harts_0_timerInterrupt <= (logic_harts_0_cmp <= logic_time);
    logic_harts_1_timerInterrupt <= (logic_harts_1_cmp <= logic_time);
    if(when_BmbSlaveFactory_l77_2) begin
      if(factory_doWrite) begin
        logic_harts_0_cmp[31 : 0] <= io_bus_cmd_payload_fragment_data[31 : 0];
      end
    end
    if(when_BmbSlaveFactory_l77_3) begin
      if(factory_doWrite) begin
        logic_harts_0_cmp[63 : 32] <= io_bus_cmd_payload_fragment_data[31 : 0];
      end
    end
    if(when_BmbSlaveFactory_l77_4) begin
      if(factory_doWrite) begin
        logic_harts_1_cmp[31 : 0] <= io_bus_cmd_payload_fragment_data[31 : 0];
      end
    end
    if(when_BmbSlaveFactory_l77_5) begin
      if(factory_doWrite) begin
        logic_harts_1_cmp[63 : 32] <= io_bus_cmd_payload_fragment_data[31 : 0];
      end
    end
  end


endmodule

module BmbDecoder_1 (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [23:0]   io_input_cmd_payload_fragment_address,
  input  wire [1:0]    io_input_cmd_payload_fragment_length,
  input  wire [31:0]   io_input_cmd_payload_fragment_data,
  input  wire [3:0]    io_input_cmd_payload_fragment_mask,
  input  wire [48:0]   io_input_cmd_payload_fragment_context,
  output reg           io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output reg           io_input_rsp_payload_last,
  output reg  [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [31:0]   io_input_rsp_payload_fragment_data,
  output reg  [48:0]   io_input_rsp_payload_fragment_context,
  output reg           io_outputs_0_cmd_valid,
  input  wire          io_outputs_0_cmd_ready,
  output wire          io_outputs_0_cmd_payload_last,
  output wire [0:0]    io_outputs_0_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_0_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_0_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_0_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_0_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_0_cmd_payload_fragment_context,
  input  wire          io_outputs_0_rsp_valid,
  output wire          io_outputs_0_rsp_ready,
  input  wire          io_outputs_0_rsp_payload_last,
  input  wire [0:0]    io_outputs_0_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_0_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_0_rsp_payload_fragment_context,
  output reg           io_outputs_1_cmd_valid,
  input  wire          io_outputs_1_cmd_ready,
  output wire          io_outputs_1_cmd_payload_last,
  output wire [0:0]    io_outputs_1_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_1_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_1_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_1_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_1_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_1_cmd_payload_fragment_context,
  input  wire          io_outputs_1_rsp_valid,
  output wire          io_outputs_1_rsp_ready,
  input  wire          io_outputs_1_rsp_payload_last,
  input  wire [0:0]    io_outputs_1_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_1_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_1_rsp_payload_fragment_context,
  output reg           io_outputs_2_cmd_valid,
  input  wire          io_outputs_2_cmd_ready,
  output wire          io_outputs_2_cmd_payload_last,
  output wire [0:0]    io_outputs_2_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_2_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_2_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_2_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_2_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_2_cmd_payload_fragment_context,
  input  wire          io_outputs_2_rsp_valid,
  output wire          io_outputs_2_rsp_ready,
  input  wire          io_outputs_2_rsp_payload_last,
  input  wire [0:0]    io_outputs_2_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_2_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_2_rsp_payload_fragment_context,
  output reg           io_outputs_3_cmd_valid,
  input  wire          io_outputs_3_cmd_ready,
  output wire          io_outputs_3_cmd_payload_last,
  output wire [0:0]    io_outputs_3_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_3_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_3_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_3_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_3_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_3_cmd_payload_fragment_context,
  input  wire          io_outputs_3_rsp_valid,
  output wire          io_outputs_3_rsp_ready,
  input  wire          io_outputs_3_rsp_payload_last,
  input  wire [0:0]    io_outputs_3_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_3_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_3_rsp_payload_fragment_context,
  output reg           io_outputs_4_cmd_valid,
  input  wire          io_outputs_4_cmd_ready,
  output wire          io_outputs_4_cmd_payload_last,
  output wire [0:0]    io_outputs_4_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_4_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_4_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_4_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_4_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_4_cmd_payload_fragment_context,
  input  wire          io_outputs_4_rsp_valid,
  output wire          io_outputs_4_rsp_ready,
  input  wire          io_outputs_4_rsp_payload_last,
  input  wire [0:0]    io_outputs_4_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_4_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_4_rsp_payload_fragment_context,
  output reg           io_outputs_5_cmd_valid,
  input  wire          io_outputs_5_cmd_ready,
  output wire          io_outputs_5_cmd_payload_last,
  output wire [0:0]    io_outputs_5_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_5_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_5_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_5_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_5_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_5_cmd_payload_fragment_context,
  input  wire          io_outputs_5_rsp_valid,
  output wire          io_outputs_5_rsp_ready,
  input  wire          io_outputs_5_rsp_payload_last,
  input  wire [0:0]    io_outputs_5_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_5_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_5_rsp_payload_fragment_context,
  output reg           io_outputs_6_cmd_valid,
  input  wire          io_outputs_6_cmd_ready,
  output wire          io_outputs_6_cmd_payload_last,
  output wire [0:0]    io_outputs_6_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_6_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_6_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_6_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_6_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_6_cmd_payload_fragment_context,
  input  wire          io_outputs_6_rsp_valid,
  output wire          io_outputs_6_rsp_ready,
  input  wire          io_outputs_6_rsp_payload_last,
  input  wire [0:0]    io_outputs_6_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_6_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_6_rsp_payload_fragment_context,
  output reg           io_outputs_7_cmd_valid,
  input  wire          io_outputs_7_cmd_ready,
  output wire          io_outputs_7_cmd_payload_last,
  output wire [0:0]    io_outputs_7_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_7_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_7_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_7_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_7_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_7_cmd_payload_fragment_context,
  input  wire          io_outputs_7_rsp_valid,
  output wire          io_outputs_7_rsp_ready,
  input  wire          io_outputs_7_rsp_payload_last,
  input  wire [0:0]    io_outputs_7_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_7_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_7_rsp_payload_fragment_context,
  output reg           io_outputs_8_cmd_valid,
  input  wire          io_outputs_8_cmd_ready,
  output wire          io_outputs_8_cmd_payload_last,
  output wire [0:0]    io_outputs_8_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_8_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_8_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_8_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_8_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_8_cmd_payload_fragment_context,
  input  wire          io_outputs_8_rsp_valid,
  output wire          io_outputs_8_rsp_ready,
  input  wire          io_outputs_8_rsp_payload_last,
  input  wire [0:0]    io_outputs_8_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_8_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_8_rsp_payload_fragment_context,
  output reg           io_outputs_9_cmd_valid,
  input  wire          io_outputs_9_cmd_ready,
  output wire          io_outputs_9_cmd_payload_last,
  output wire [0:0]    io_outputs_9_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_9_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_9_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_9_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_9_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_9_cmd_payload_fragment_context,
  input  wire          io_outputs_9_rsp_valid,
  output wire          io_outputs_9_rsp_ready,
  input  wire          io_outputs_9_rsp_payload_last,
  input  wire [0:0]    io_outputs_9_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_9_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_9_rsp_payload_fragment_context,
  output reg           io_outputs_10_cmd_valid,
  input  wire          io_outputs_10_cmd_ready,
  output wire          io_outputs_10_cmd_payload_last,
  output wire [0:0]    io_outputs_10_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_10_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_10_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_10_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_10_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_10_cmd_payload_fragment_context,
  input  wire          io_outputs_10_rsp_valid,
  output wire          io_outputs_10_rsp_ready,
  input  wire          io_outputs_10_rsp_payload_last,
  input  wire [0:0]    io_outputs_10_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_10_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_10_rsp_payload_fragment_context,
  output reg           io_outputs_11_cmd_valid,
  input  wire          io_outputs_11_cmd_ready,
  output wire          io_outputs_11_cmd_payload_last,
  output wire [0:0]    io_outputs_11_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_11_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_11_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_11_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_11_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_11_cmd_payload_fragment_context,
  input  wire          io_outputs_11_rsp_valid,
  output wire          io_outputs_11_rsp_ready,
  input  wire          io_outputs_11_rsp_payload_last,
  input  wire [0:0]    io_outputs_11_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_11_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_11_rsp_payload_fragment_context,
  output reg           io_outputs_12_cmd_valid,
  input  wire          io_outputs_12_cmd_ready,
  output wire          io_outputs_12_cmd_payload_last,
  output wire [0:0]    io_outputs_12_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_12_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_12_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_12_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_12_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_12_cmd_payload_fragment_context,
  input  wire          io_outputs_12_rsp_valid,
  output wire          io_outputs_12_rsp_ready,
  input  wire          io_outputs_12_rsp_payload_last,
  input  wire [0:0]    io_outputs_12_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_12_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_12_rsp_payload_fragment_context,
  output reg           io_outputs_13_cmd_valid,
  input  wire          io_outputs_13_cmd_ready,
  output wire          io_outputs_13_cmd_payload_last,
  output wire [0:0]    io_outputs_13_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_13_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_13_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_13_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_13_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_13_cmd_payload_fragment_context,
  input  wire          io_outputs_13_rsp_valid,
  output wire          io_outputs_13_rsp_ready,
  input  wire          io_outputs_13_rsp_payload_last,
  input  wire [0:0]    io_outputs_13_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_13_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_13_rsp_payload_fragment_context,
  output reg           io_outputs_14_cmd_valid,
  input  wire          io_outputs_14_cmd_ready,
  output wire          io_outputs_14_cmd_payload_last,
  output wire [0:0]    io_outputs_14_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_14_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_14_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_14_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_14_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_14_cmd_payload_fragment_context,
  input  wire          io_outputs_14_rsp_valid,
  output wire          io_outputs_14_rsp_ready,
  input  wire          io_outputs_14_rsp_payload_last,
  input  wire [0:0]    io_outputs_14_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_14_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_14_rsp_payload_fragment_context,
  output reg           io_outputs_15_cmd_valid,
  input  wire          io_outputs_15_cmd_ready,
  output wire          io_outputs_15_cmd_payload_last,
  output wire [0:0]    io_outputs_15_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_15_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_15_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_15_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_15_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_15_cmd_payload_fragment_context,
  input  wire          io_outputs_15_rsp_valid,
  output wire          io_outputs_15_rsp_ready,
  input  wire          io_outputs_15_rsp_payload_last,
  input  wire [0:0]    io_outputs_15_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_15_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_15_rsp_payload_fragment_context,
  output reg           io_outputs_16_cmd_valid,
  input  wire          io_outputs_16_cmd_ready,
  output wire          io_outputs_16_cmd_payload_last,
  output wire [0:0]    io_outputs_16_cmd_payload_fragment_opcode,
  output wire [23:0]   io_outputs_16_cmd_payload_fragment_address,
  output wire [1:0]    io_outputs_16_cmd_payload_fragment_length,
  output wire [31:0]   io_outputs_16_cmd_payload_fragment_data,
  output wire [3:0]    io_outputs_16_cmd_payload_fragment_mask,
  output wire [48:0]   io_outputs_16_cmd_payload_fragment_context,
  input  wire          io_outputs_16_rsp_valid,
  output wire          io_outputs_16_rsp_ready,
  input  wire          io_outputs_16_rsp_payload_last,
  input  wire [0:0]    io_outputs_16_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_outputs_16_rsp_payload_fragment_data,
  input  wire [48:0]   io_outputs_16_rsp_payload_fragment_context,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire       [0:0]    _zz_logic_noHitS0;
  wire       [6:0]    _zz_logic_noHitS0_1;
  wire                _zz_logic_input_ready;
  wire       [0:0]    _zz_logic_input_ready_1;
  wire       [9:0]    _zz_logic_input_ready_2;
  wire                _zz_logic_input_ready_3;
  wire       [0:0]    _zz_logic_input_ready_4;
  wire       [2:0]    _zz_logic_input_ready_5;
  wire       [3:0]    _zz_logic_rspPendingCounter;
  wire       [3:0]    _zz_logic_rspPendingCounter_1;
  wire       [0:0]    _zz_logic_rspPendingCounter_2;
  wire       [3:0]    _zz_logic_rspPendingCounter_3;
  wire       [0:0]    _zz_logic_rspPendingCounter_4;
  wire       [0:0]    _zz_logic_rspNoHitValid;
  wire       [6:0]    _zz_logic_rspNoHitValid_1;
  wire       [0:0]    _zz_io_input_rsp_valid;
  wire       [7:0]    _zz_io_input_rsp_valid_1;
  reg                 _zz_io_input_rsp_payload_last_5;
  reg        [0:0]    _zz_io_input_rsp_payload_fragment_opcode;
  reg        [31:0]   _zz_io_input_rsp_payload_fragment_data;
  reg        [48:0]   _zz_io_input_rsp_payload_fragment_context;
  wire                _zz_logic_cmdWait;
  wire                _zz_logic_cmdWait_1;
  wire                _zz_logic_cmdWait_2;
  wire                _zz_logic_cmdWait_3;
  wire                logic_input_valid;
  reg                 logic_input_ready;
  wire                logic_input_payload_last;
  wire       [0:0]    logic_input_payload_fragment_opcode;
  wire       [23:0]   logic_input_payload_fragment_address;
  wire       [1:0]    logic_input_payload_fragment_length;
  wire       [31:0]   logic_input_payload_fragment_data;
  wire       [3:0]    logic_input_payload_fragment_mask;
  wire       [48:0]   logic_input_payload_fragment_context;
  reg                 io_input_cmd_rValid;
  wire                logic_input_fire;
  reg                 io_input_cmd_rData_last;
  reg        [0:0]    io_input_cmd_rData_fragment_opcode;
  reg        [23:0]   io_input_cmd_rData_fragment_address;
  reg        [1:0]    io_input_cmd_rData_fragment_length;
  reg        [31:0]   io_input_cmd_rData_fragment_data;
  reg        [3:0]    io_input_cmd_rData_fragment_mask;
  reg        [48:0]   io_input_cmd_rData_fragment_context;
  wire                logic_hitsS0_0;
  wire                logic_hitsS0_1;
  wire                logic_hitsS0_2;
  wire                logic_hitsS0_3;
  wire                logic_hitsS0_4;
  wire                logic_hitsS0_5;
  wire                logic_hitsS0_6;
  wire                logic_hitsS0_7;
  wire                logic_hitsS0_8;
  wire                logic_hitsS0_9;
  wire                logic_hitsS0_10;
  wire                logic_hitsS0_11;
  wire                logic_hitsS0_12;
  wire                logic_hitsS0_13;
  wire                logic_hitsS0_14;
  wire                logic_hitsS0_15;
  wire                logic_hitsS0_16;
  wire                logic_noHitS0;
  wire                io_input_cmd_fire;
  reg                 logic_hitsS1_0;
  reg                 logic_hitsS1_1;
  reg                 logic_hitsS1_2;
  reg                 logic_hitsS1_3;
  reg                 logic_hitsS1_4;
  reg                 logic_hitsS1_5;
  reg                 logic_hitsS1_6;
  reg                 logic_hitsS1_7;
  reg                 logic_hitsS1_8;
  reg                 logic_hitsS1_9;
  reg                 logic_hitsS1_10;
  reg                 logic_hitsS1_11;
  reg                 logic_hitsS1_12;
  reg                 logic_hitsS1_13;
  reg                 logic_hitsS1_14;
  reg                 logic_hitsS1_15;
  reg                 logic_hitsS1_16;
  reg                 logic_noHitS1;
  wire                _zz_io_outputs_0_cmd_payload_last;
  wire                _zz_io_outputs_1_cmd_payload_last;
  wire                _zz_io_outputs_2_cmd_payload_last;
  wire                _zz_io_outputs_3_cmd_payload_last;
  wire                _zz_io_outputs_4_cmd_payload_last;
  wire                _zz_io_outputs_5_cmd_payload_last;
  wire                _zz_io_outputs_6_cmd_payload_last;
  wire                _zz_io_outputs_7_cmd_payload_last;
  wire                _zz_io_outputs_8_cmd_payload_last;
  wire                _zz_io_outputs_9_cmd_payload_last;
  wire                _zz_io_outputs_10_cmd_payload_last;
  wire                _zz_io_outputs_11_cmd_payload_last;
  wire                _zz_io_outputs_12_cmd_payload_last;
  wire                _zz_io_outputs_13_cmd_payload_last;
  wire                _zz_io_outputs_14_cmd_payload_last;
  wire                _zz_io_outputs_15_cmd_payload_last;
  wire                _zz_io_outputs_16_cmd_payload_last;
  reg        [3:0]    logic_rspPendingCounter;
  wire                io_input_rsp_fire;
  wire                logic_cmdWait;
  wire                when_BmbDecoder_l56;
  reg                 logic_rspHits_0;
  reg                 logic_rspHits_1;
  reg                 logic_rspHits_2;
  reg                 logic_rspHits_3;
  reg                 logic_rspHits_4;
  reg                 logic_rspHits_5;
  reg                 logic_rspHits_6;
  reg                 logic_rspHits_7;
  reg                 logic_rspHits_8;
  reg                 logic_rspHits_9;
  reg                 logic_rspHits_10;
  reg                 logic_rspHits_11;
  reg                 logic_rspHits_12;
  reg                 logic_rspHits_13;
  reg                 logic_rspHits_14;
  reg                 logic_rspHits_15;
  reg                 logic_rspHits_16;
  wire                logic_rspPending;
  wire                logic_rspNoHitValid;
  reg                 logic_rspNoHit_doIt;
  wire                when_BmbDecoder_l60;
  wire                when_BmbDecoder_l60_1;
  reg                 logic_rspNoHit_singleBeatRsp;
  reg        [48:0]   logic_rspNoHit_context;
  wire                _zz_io_input_rsp_payload_last;
  wire                _zz_io_input_rsp_payload_last_1;
  wire                _zz_io_input_rsp_payload_last_2;
  wire                _zz_io_input_rsp_payload_last_3;
  wire       [4:0]    _zz_io_input_rsp_payload_last_4;

  assign _zz_logic_rspPendingCounter = (logic_rspPendingCounter + _zz_logic_rspPendingCounter_1);
  assign _zz_logic_rspPendingCounter_2 = (logic_input_fire && logic_input_payload_last);
  assign _zz_logic_rspPendingCounter_1 = {3'd0, _zz_logic_rspPendingCounter_2};
  assign _zz_logic_rspPendingCounter_4 = (io_input_rsp_fire && io_input_rsp_payload_last);
  assign _zz_logic_rspPendingCounter_3 = {3'd0, _zz_logic_rspPendingCounter_4};
  assign _zz_logic_noHitS0 = logic_hitsS0_7;
  assign _zz_logic_noHitS0_1 = {logic_hitsS0_6,{logic_hitsS0_5,{logic_hitsS0_4,{logic_hitsS0_3,{logic_hitsS0_2,{logic_hitsS0_1,logic_hitsS0_0}}}}}};
  assign _zz_logic_input_ready = (logic_hitsS1_11 && io_outputs_11_cmd_ready);
  assign _zz_logic_input_ready_1 = (logic_hitsS1_10 && io_outputs_10_cmd_ready);
  assign _zz_logic_input_ready_2 = {(logic_hitsS1_9 && io_outputs_9_cmd_ready),{(logic_hitsS1_8 && io_outputs_8_cmd_ready),{(logic_hitsS1_7 && io_outputs_7_cmd_ready),{(logic_hitsS1_6 && io_outputs_6_cmd_ready),{(logic_hitsS1_5 && io_outputs_5_cmd_ready),{_zz_logic_input_ready_3,{_zz_logic_input_ready_4,_zz_logic_input_ready_5}}}}}}};
  assign _zz_logic_input_ready_3 = (logic_hitsS1_4 && io_outputs_4_cmd_ready);
  assign _zz_logic_input_ready_4 = (logic_hitsS1_3 && io_outputs_3_cmd_ready);
  assign _zz_logic_input_ready_5 = {(logic_hitsS1_2 && io_outputs_2_cmd_ready),{(logic_hitsS1_1 && io_outputs_1_cmd_ready),(logic_hitsS1_0 && io_outputs_0_cmd_ready)}};
  assign _zz_logic_rspNoHitValid = logic_rspHits_7;
  assign _zz_logic_rspNoHitValid_1 = {logic_rspHits_6,{logic_rspHits_5,{logic_rspHits_4,{logic_rspHits_3,{logic_rspHits_2,{logic_rspHits_1,logic_rspHits_0}}}}}};
  assign _zz_io_input_rsp_valid = io_outputs_8_rsp_valid;
  assign _zz_io_input_rsp_valid_1 = {io_outputs_7_rsp_valid,{io_outputs_6_rsp_valid,{io_outputs_5_rsp_valid,{io_outputs_4_rsp_valid,{io_outputs_3_rsp_valid,{io_outputs_2_rsp_valid,{io_outputs_1_rsp_valid,io_outputs_0_rsp_valid}}}}}}};
  assign _zz_logic_cmdWait = (((((((((_zz_logic_cmdWait_1 || _zz_logic_cmdWait_2) || (logic_hitsS1_2 != logic_rspHits_2)) || (logic_hitsS1_3 != logic_rspHits_3)) || (logic_hitsS1_4 != logic_rspHits_4)) || (logic_hitsS1_5 != logic_rspHits_5)) || (logic_hitsS1_6 != logic_rspHits_6)) || (logic_hitsS1_7 != logic_rspHits_7)) || (logic_hitsS1_8 != logic_rspHits_8)) || (logic_hitsS1_9 != logic_rspHits_9));
  assign _zz_logic_cmdWait_3 = (logic_hitsS1_10 != logic_rspHits_10);
  assign _zz_logic_cmdWait_1 = (logic_hitsS1_0 != logic_rspHits_0);
  assign _zz_logic_cmdWait_2 = (logic_hitsS1_1 != logic_rspHits_1);
  always @(*) begin
    case(_zz_io_input_rsp_payload_last_4)
      5'b00000 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_0_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_0_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_0_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_0_rsp_payload_fragment_context;
      end
      5'b00001 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_1_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_1_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_1_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_1_rsp_payload_fragment_context;
      end
      5'b00010 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_2_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_2_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_2_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_2_rsp_payload_fragment_context;
      end
      5'b00011 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_3_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_3_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_3_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_3_rsp_payload_fragment_context;
      end
      5'b00100 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_4_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_4_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_4_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_4_rsp_payload_fragment_context;
      end
      5'b00101 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_5_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_5_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_5_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_5_rsp_payload_fragment_context;
      end
      5'b00110 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_6_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_6_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_6_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_6_rsp_payload_fragment_context;
      end
      5'b00111 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_7_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_7_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_7_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_7_rsp_payload_fragment_context;
      end
      5'b01000 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_8_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_8_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_8_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_8_rsp_payload_fragment_context;
      end
      5'b01001 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_9_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_9_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_9_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_9_rsp_payload_fragment_context;
      end
      5'b01010 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_10_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_10_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_10_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_10_rsp_payload_fragment_context;
      end
      5'b01011 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_11_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_11_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_11_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_11_rsp_payload_fragment_context;
      end
      5'b01100 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_12_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_12_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_12_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_12_rsp_payload_fragment_context;
      end
      5'b01101 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_13_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_13_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_13_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_13_rsp_payload_fragment_context;
      end
      5'b01110 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_14_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_14_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_14_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_14_rsp_payload_fragment_context;
      end
      5'b01111 : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_15_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_15_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_15_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_15_rsp_payload_fragment_context;
      end
      default : begin
        _zz_io_input_rsp_payload_last_5 = io_outputs_16_rsp_payload_last;
        _zz_io_input_rsp_payload_fragment_opcode = io_outputs_16_rsp_payload_fragment_opcode;
        _zz_io_input_rsp_payload_fragment_data = io_outputs_16_rsp_payload_fragment_data;
        _zz_io_input_rsp_payload_fragment_context = io_outputs_16_rsp_payload_fragment_context;
      end
    endcase
  end

  assign logic_input_fire = (logic_input_valid && logic_input_ready);
  assign io_input_cmd_ready = (! io_input_cmd_rValid);
  assign logic_input_valid = io_input_cmd_rValid;
  assign logic_input_payload_last = io_input_cmd_rData_last;
  assign logic_input_payload_fragment_opcode = io_input_cmd_rData_fragment_opcode;
  assign logic_input_payload_fragment_address = io_input_cmd_rData_fragment_address;
  assign logic_input_payload_fragment_length = io_input_cmd_rData_fragment_length;
  assign logic_input_payload_fragment_data = io_input_cmd_rData_fragment_data;
  assign logic_input_payload_fragment_mask = io_input_cmd_rData_fragment_mask;
  assign logic_input_payload_fragment_context = io_input_cmd_rData_fragment_context;
  assign logic_noHitS0 = (! (|{logic_hitsS0_16,{logic_hitsS0_15,{logic_hitsS0_14,{logic_hitsS0_13,{logic_hitsS0_12,{logic_hitsS0_11,{logic_hitsS0_10,{logic_hitsS0_9,{logic_hitsS0_8,{_zz_logic_noHitS0,_zz_logic_noHitS0_1}}}}}}}}}}));
  assign io_input_cmd_fire = (io_input_cmd_valid && io_input_cmd_ready);
  assign logic_hitsS0_0 = ((io_input_cmd_payload_fragment_address & (~ 24'h3fffff)) == 24'hc00000);
  always @(*) begin
    io_outputs_0_cmd_valid = (logic_input_valid && logic_hitsS1_0);
    if(logic_cmdWait) begin
      io_outputs_0_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_0_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_0_cmd_payload_last = _zz_io_outputs_0_cmd_payload_last;
  assign io_outputs_0_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_0_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_0_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_0_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_0_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_0_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_1 = ((io_input_cmd_payload_fragment_address & (~ 24'h00ffff)) == 24'hb00000);
  always @(*) begin
    io_outputs_1_cmd_valid = (logic_input_valid && logic_hitsS1_1);
    if(logic_cmdWait) begin
      io_outputs_1_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_1_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_1_cmd_payload_last = _zz_io_outputs_1_cmd_payload_last;
  assign io_outputs_1_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_1_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_1_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_1_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_1_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_1_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_2 = ((io_input_cmd_payload_fragment_address & (~ 24'h00003f)) == 24'h010000);
  always @(*) begin
    io_outputs_2_cmd_valid = (logic_input_valid && logic_hitsS1_2);
    if(logic_cmdWait) begin
      io_outputs_2_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_2_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_2_cmd_payload_last = _zz_io_outputs_2_cmd_payload_last;
  assign io_outputs_2_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_2_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_2_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_2_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_2_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_2_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_3 = ((io_input_cmd_payload_fragment_address & (~ 24'h000fff)) == 24'h014000);
  always @(*) begin
    io_outputs_3_cmd_valid = (logic_input_valid && logic_hitsS1_3);
    if(logic_cmdWait) begin
      io_outputs_3_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_3_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_3_cmd_payload_last = _zz_io_outputs_3_cmd_payload_last;
  assign io_outputs_3_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_3_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_3_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_3_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_3_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_3_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_4 = ((io_input_cmd_payload_fragment_address & (~ 24'h000fff)) == 24'h015000);
  always @(*) begin
    io_outputs_4_cmd_valid = (logic_input_valid && logic_hitsS1_4);
    if(logic_cmdWait) begin
      io_outputs_4_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_4_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_4_cmd_payload_last = _zz_io_outputs_4_cmd_payload_last;
  assign io_outputs_4_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_4_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_4_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_4_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_4_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_4_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_5 = ((io_input_cmd_payload_fragment_address & (~ 24'h0000ff)) == 24'h017000);
  always @(*) begin
    io_outputs_5_cmd_valid = (logic_input_valid && logic_hitsS1_5);
    if(logic_cmdWait) begin
      io_outputs_5_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_5_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_5_cmd_payload_last = _zz_io_outputs_5_cmd_payload_last;
  assign io_outputs_5_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_5_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_5_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_5_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_5_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_5_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_6 = ((io_input_cmd_payload_fragment_address & (~ 24'h0000ff)) == 24'h019000);
  always @(*) begin
    io_outputs_6_cmd_valid = (logic_input_valid && logic_hitsS1_6);
    if(logic_cmdWait) begin
      io_outputs_6_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_6_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_6_cmd_payload_last = _zz_io_outputs_6_cmd_payload_last;
  assign io_outputs_6_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_6_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_6_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_6_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_6_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_6_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_7 = ((io_input_cmd_payload_fragment_address & (~ 24'h0000ff)) == 24'h018000);
  always @(*) begin
    io_outputs_7_cmd_valid = (logic_input_valid && logic_hitsS1_7);
    if(logic_cmdWait) begin
      io_outputs_7_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_7_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_7_cmd_payload_last = _zz_io_outputs_7_cmd_payload_last;
  assign io_outputs_7_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_7_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_7_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_7_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_7_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_7_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_8 = ((io_input_cmd_payload_fragment_address & (~ 24'h000fff)) == 24'h01b000);
  always @(*) begin
    io_outputs_8_cmd_valid = (logic_input_valid && logic_hitsS1_8);
    if(logic_cmdWait) begin
      io_outputs_8_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_8_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_8_cmd_payload_last = _zz_io_outputs_8_cmd_payload_last;
  assign io_outputs_8_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_8_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_8_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_8_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_8_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_8_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_9 = ((io_input_cmd_payload_fragment_address & (~ 24'h000fff)) == 24'h01a000);
  always @(*) begin
    io_outputs_9_cmd_valid = (logic_input_valid && logic_hitsS1_9);
    if(logic_cmdWait) begin
      io_outputs_9_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_9_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_9_cmd_payload_last = _zz_io_outputs_9_cmd_payload_last;
  assign io_outputs_9_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_9_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_9_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_9_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_9_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_9_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_10 = ((io_input_cmd_payload_fragment_address & (~ 24'h0000ff)) == 24'h016000);
  always @(*) begin
    io_outputs_10_cmd_valid = (logic_input_valid && logic_hitsS1_10);
    if(logic_cmdWait) begin
      io_outputs_10_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_10_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_10_cmd_payload_last = _zz_io_outputs_10_cmd_payload_last;
  assign io_outputs_10_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_10_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_10_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_10_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_10_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_10_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_11 = ((io_input_cmd_payload_fragment_address & (~ 24'h0000ff)) == 24'h01c000);
  always @(*) begin
    io_outputs_11_cmd_valid = (logic_input_valid && logic_hitsS1_11);
    if(logic_cmdWait) begin
      io_outputs_11_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_11_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_11_cmd_payload_last = _zz_io_outputs_11_cmd_payload_last;
  assign io_outputs_11_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_11_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_11_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_11_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_11_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_11_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_12 = ((io_input_cmd_payload_fragment_address & (~ 24'h00ffff)) == 24'h120000);
  always @(*) begin
    io_outputs_12_cmd_valid = (logic_input_valid && logic_hitsS1_12);
    if(logic_cmdWait) begin
      io_outputs_12_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_12_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_12_cmd_payload_last = _zz_io_outputs_12_cmd_payload_last;
  assign io_outputs_12_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_12_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_12_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_12_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_12_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_12_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_13 = ((io_input_cmd_payload_fragment_address & (~ 24'h00ffff)) == 24'h110000);
  always @(*) begin
    io_outputs_13_cmd_valid = (logic_input_valid && logic_hitsS1_13);
    if(logic_cmdWait) begin
      io_outputs_13_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_13_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_13_cmd_payload_last = _zz_io_outputs_13_cmd_payload_last;
  assign io_outputs_13_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_13_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_13_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_13_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_13_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_13_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_14 = ((io_input_cmd_payload_fragment_address & (~ 24'h00ffff)) == 24'h140000);
  always @(*) begin
    io_outputs_14_cmd_valid = (logic_input_valid && logic_hitsS1_14);
    if(logic_cmdWait) begin
      io_outputs_14_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_14_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_14_cmd_payload_last = _zz_io_outputs_14_cmd_payload_last;
  assign io_outputs_14_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_14_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_14_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_14_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_14_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_14_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_15 = ((io_input_cmd_payload_fragment_address & (~ 24'h00ffff)) == 24'h100000);
  always @(*) begin
    io_outputs_15_cmd_valid = (logic_input_valid && logic_hitsS1_15);
    if(logic_cmdWait) begin
      io_outputs_15_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_15_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_15_cmd_payload_last = _zz_io_outputs_15_cmd_payload_last;
  assign io_outputs_15_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_15_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_15_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_15_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_15_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_15_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  assign logic_hitsS0_16 = ((io_input_cmd_payload_fragment_address & (~ 24'h00ffff)) == 24'h130000);
  always @(*) begin
    io_outputs_16_cmd_valid = (logic_input_valid && logic_hitsS1_16);
    if(logic_cmdWait) begin
      io_outputs_16_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_16_cmd_payload_last = logic_input_payload_last;
  assign io_outputs_16_cmd_payload_last = _zz_io_outputs_16_cmd_payload_last;
  assign io_outputs_16_cmd_payload_fragment_opcode = logic_input_payload_fragment_opcode;
  assign io_outputs_16_cmd_payload_fragment_address = logic_input_payload_fragment_address;
  assign io_outputs_16_cmd_payload_fragment_length = logic_input_payload_fragment_length;
  assign io_outputs_16_cmd_payload_fragment_data = logic_input_payload_fragment_data;
  assign io_outputs_16_cmd_payload_fragment_mask = logic_input_payload_fragment_mask;
  assign io_outputs_16_cmd_payload_fragment_context = logic_input_payload_fragment_context;
  always @(*) begin
    logic_input_ready = ((|{(logic_hitsS1_16 && io_outputs_16_cmd_ready),{(logic_hitsS1_15 && io_outputs_15_cmd_ready),{(logic_hitsS1_14 && io_outputs_14_cmd_ready),{(logic_hitsS1_13 && io_outputs_13_cmd_ready),{(logic_hitsS1_12 && io_outputs_12_cmd_ready),{_zz_logic_input_ready,{_zz_logic_input_ready_1,_zz_logic_input_ready_2}}}}}}}) || logic_noHitS1);
    if(logic_cmdWait) begin
      logic_input_ready = 1'b0;
    end
  end

  assign io_input_rsp_fire = (io_input_rsp_valid && io_input_rsp_ready);
  assign when_BmbDecoder_l56 = (logic_input_valid && (! logic_cmdWait));
  assign logic_rspPending = (logic_rspPendingCounter != 4'b0000);
  assign logic_rspNoHitValid = (! (|{logic_rspHits_16,{logic_rspHits_15,{logic_rspHits_14,{logic_rspHits_13,{logic_rspHits_12,{logic_rspHits_11,{logic_rspHits_10,{logic_rspHits_9,{logic_rspHits_8,{_zz_logic_rspNoHitValid,_zz_logic_rspNoHitValid_1}}}}}}}}}}));
  assign when_BmbDecoder_l60 = (io_input_rsp_fire && io_input_rsp_payload_last);
  assign when_BmbDecoder_l60_1 = ((logic_input_fire && logic_noHitS1) && logic_input_payload_last);
  always @(*) begin
    io_input_rsp_valid = ((|{io_outputs_16_rsp_valid,{io_outputs_15_rsp_valid,{io_outputs_14_rsp_valid,{io_outputs_13_rsp_valid,{io_outputs_12_rsp_valid,{io_outputs_11_rsp_valid,{io_outputs_10_rsp_valid,{io_outputs_9_rsp_valid,{_zz_io_input_rsp_valid,_zz_io_input_rsp_valid_1}}}}}}}}}) || (logic_rspPending && logic_rspNoHitValid));
    if(logic_rspNoHit_doIt) begin
      io_input_rsp_valid = 1'b1;
    end
  end

  assign _zz_io_input_rsp_payload_last = (((((((logic_rspHits_1 || logic_rspHits_3) || logic_rspHits_5) || logic_rspHits_7) || logic_rspHits_9) || logic_rspHits_11) || logic_rspHits_13) || logic_rspHits_15);
  assign _zz_io_input_rsp_payload_last_1 = (((((((logic_rspHits_2 || logic_rspHits_3) || logic_rspHits_6) || logic_rspHits_7) || logic_rspHits_10) || logic_rspHits_11) || logic_rspHits_14) || logic_rspHits_15);
  assign _zz_io_input_rsp_payload_last_2 = (((((((logic_rspHits_4 || logic_rspHits_5) || logic_rspHits_6) || logic_rspHits_7) || logic_rspHits_12) || logic_rspHits_13) || logic_rspHits_14) || logic_rspHits_15);
  assign _zz_io_input_rsp_payload_last_3 = (((((((logic_rspHits_8 || logic_rspHits_9) || logic_rspHits_10) || logic_rspHits_11) || logic_rspHits_12) || logic_rspHits_13) || logic_rspHits_14) || logic_rspHits_15);
  assign _zz_io_input_rsp_payload_last_4 = {logic_rspHits_16,{_zz_io_input_rsp_payload_last_3,{_zz_io_input_rsp_payload_last_2,{_zz_io_input_rsp_payload_last_1,_zz_io_input_rsp_payload_last}}}};
  always @(*) begin
    io_input_rsp_payload_last = _zz_io_input_rsp_payload_last_5;
    if(logic_rspNoHit_doIt) begin
      io_input_rsp_payload_last = 1'b1;
    end
  end

  always @(*) begin
    io_input_rsp_payload_fragment_opcode = _zz_io_input_rsp_payload_fragment_opcode;
    if(logic_rspNoHit_doIt) begin
      io_input_rsp_payload_fragment_opcode = 1'b1;
    end
  end

  assign io_input_rsp_payload_fragment_data = _zz_io_input_rsp_payload_fragment_data;
  always @(*) begin
    io_input_rsp_payload_fragment_context = _zz_io_input_rsp_payload_fragment_context;
    if(logic_rspNoHit_doIt) begin
      io_input_rsp_payload_fragment_context = logic_rspNoHit_context;
    end
  end

  assign io_outputs_0_rsp_ready = io_input_rsp_ready;
  assign io_outputs_1_rsp_ready = io_input_rsp_ready;
  assign io_outputs_2_rsp_ready = io_input_rsp_ready;
  assign io_outputs_3_rsp_ready = io_input_rsp_ready;
  assign io_outputs_4_rsp_ready = io_input_rsp_ready;
  assign io_outputs_5_rsp_ready = io_input_rsp_ready;
  assign io_outputs_6_rsp_ready = io_input_rsp_ready;
  assign io_outputs_7_rsp_ready = io_input_rsp_ready;
  assign io_outputs_8_rsp_ready = io_input_rsp_ready;
  assign io_outputs_9_rsp_ready = io_input_rsp_ready;
  assign io_outputs_10_rsp_ready = io_input_rsp_ready;
  assign io_outputs_11_rsp_ready = io_input_rsp_ready;
  assign io_outputs_12_rsp_ready = io_input_rsp_ready;
  assign io_outputs_13_rsp_ready = io_input_rsp_ready;
  assign io_outputs_14_rsp_ready = io_input_rsp_ready;
  assign io_outputs_15_rsp_ready = io_input_rsp_ready;
  assign io_outputs_16_rsp_ready = io_input_rsp_ready;
  assign logic_cmdWait = ((logic_rspPending && ((((((((_zz_logic_cmdWait || _zz_logic_cmdWait_3) || (logic_hitsS1_11 != logic_rspHits_11)) || (logic_hitsS1_12 != logic_rspHits_12)) || (logic_hitsS1_13 != logic_rspHits_13)) || (logic_hitsS1_14 != logic_rspHits_14)) || (logic_hitsS1_15 != logic_rspHits_15)) || (logic_hitsS1_16 != logic_rspHits_16)) || logic_rspNoHitValid)) || (logic_rspPendingCounter == 4'b1000));
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      io_input_cmd_rValid <= 1'b0;
      logic_rspPendingCounter <= 4'b0000;
      logic_rspNoHit_doIt <= 1'b0;
    end else begin
      if(io_input_cmd_valid) begin
        io_input_cmd_rValid <= 1'b1;
      end
      if(logic_input_fire) begin
        io_input_cmd_rValid <= 1'b0;
      end
      logic_rspPendingCounter <= (_zz_logic_rspPendingCounter - _zz_logic_rspPendingCounter_3);
      if(when_BmbDecoder_l60) begin
        logic_rspNoHit_doIt <= 1'b0;
      end
      if(when_BmbDecoder_l60_1) begin
        logic_rspNoHit_doIt <= 1'b1;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(io_input_cmd_ready) begin
      io_input_cmd_rData_last <= io_input_cmd_payload_last;
      io_input_cmd_rData_fragment_opcode <= io_input_cmd_payload_fragment_opcode;
      io_input_cmd_rData_fragment_address <= io_input_cmd_payload_fragment_address;
      io_input_cmd_rData_fragment_length <= io_input_cmd_payload_fragment_length;
      io_input_cmd_rData_fragment_data <= io_input_cmd_payload_fragment_data;
      io_input_cmd_rData_fragment_mask <= io_input_cmd_payload_fragment_mask;
      io_input_cmd_rData_fragment_context <= io_input_cmd_payload_fragment_context;
    end
    if(io_input_cmd_fire) begin
      logic_hitsS1_0 <= logic_hitsS0_0;
      logic_hitsS1_1 <= logic_hitsS0_1;
      logic_hitsS1_2 <= logic_hitsS0_2;
      logic_hitsS1_3 <= logic_hitsS0_3;
      logic_hitsS1_4 <= logic_hitsS0_4;
      logic_hitsS1_5 <= logic_hitsS0_5;
      logic_hitsS1_6 <= logic_hitsS0_6;
      logic_hitsS1_7 <= logic_hitsS0_7;
      logic_hitsS1_8 <= logic_hitsS0_8;
      logic_hitsS1_9 <= logic_hitsS0_9;
      logic_hitsS1_10 <= logic_hitsS0_10;
      logic_hitsS1_11 <= logic_hitsS0_11;
      logic_hitsS1_12 <= logic_hitsS0_12;
      logic_hitsS1_13 <= logic_hitsS0_13;
      logic_hitsS1_14 <= logic_hitsS0_14;
      logic_hitsS1_15 <= logic_hitsS0_15;
      logic_hitsS1_16 <= logic_hitsS0_16;
    end
    if(io_input_cmd_fire) begin
      logic_noHitS1 <= logic_noHitS0;
    end
    if(when_BmbDecoder_l56) begin
      logic_rspHits_0 <= logic_hitsS1_0;
      logic_rspHits_1 <= logic_hitsS1_1;
      logic_rspHits_2 <= logic_hitsS1_2;
      logic_rspHits_3 <= logic_hitsS1_3;
      logic_rspHits_4 <= logic_hitsS1_4;
      logic_rspHits_5 <= logic_hitsS1_5;
      logic_rspHits_6 <= logic_hitsS1_6;
      logic_rspHits_7 <= logic_hitsS1_7;
      logic_rspHits_8 <= logic_hitsS1_8;
      logic_rspHits_9 <= logic_hitsS1_9;
      logic_rspHits_10 <= logic_hitsS1_10;
      logic_rspHits_11 <= logic_hitsS1_11;
      logic_rspHits_12 <= logic_hitsS1_12;
      logic_rspHits_13 <= logic_hitsS1_13;
      logic_rspHits_14 <= logic_hitsS1_14;
      logic_rspHits_15 <= logic_hitsS1_15;
      logic_rspHits_16 <= logic_hitsS1_16;
    end
    if(logic_input_fire) begin
      logic_rspNoHit_singleBeatRsp <= (logic_input_payload_fragment_opcode == 1'b1);
    end
    if(logic_input_fire) begin
      logic_rspNoHit_context <= logic_input_payload_fragment_context;
    end
  end


endmodule

module BmbUnburstify_1 (
  input  wire          io_input_cmd_valid,
  output reg           io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [63:0]   io_input_cmd_payload_fragment_data,
  input  wire [7:0]    io_input_cmd_payload_fragment_mask,
  input  wire [43:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire [43:0]   io_input_rsp_payload_fragment_context,
  output reg           io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output reg  [0:0]    io_output_cmd_payload_fragment_opcode,
  output reg  [31:0]   io_output_cmd_payload_fragment_address,
  output reg  [2:0]    io_output_cmd_payload_fragment_length,
  output wire [63:0]   io_output_cmd_payload_fragment_data,
  output wire [7:0]    io_output_cmd_payload_fragment_mask,
  output wire [47:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output reg           io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_output_rsp_payload_fragment_data,
  input  wire [47:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [2:0]    _zz_buffer_last;
  wire       [0:0]    _zz_buffer_last_1;
  wire       [11:0]   _zz_buffer_addressIncr;
  wire                doResult;
  reg                 buffer_valid;
  reg        [0:0]    buffer_opcode;
  reg        [1:0]    buffer_source;
  reg        [31:0]   buffer_address;
  reg        [43:0]   buffer_context;
  reg        [2:0]    buffer_beat;
  wire                buffer_last;
  wire       [31:0]   buffer_addressIncr;
  wire                buffer_isWrite;
  wire                io_output_cmd_fire;
  wire       [2:0]    cmdTransferBeatCount;
  wire                requireBuffer;
  reg                 cmdContext_drop;
  reg                 cmdContext_last;
  reg        [1:0]    cmdContext_source;
  reg        [43:0]   cmdContext_context;
  wire                rspContext_drop;
  wire                rspContext_last;
  wire       [1:0]    rspContext_source;
  wire       [43:0]   rspContext_context;
  wire       [47:0]   _zz_rspContext_drop;
  wire                when_Stream_l445;
  reg                 io_output_rsp_thrown_valid;
  wire                io_output_rsp_thrown_ready;
  wire                io_output_rsp_thrown_payload_last;
  wire       [0:0]    io_output_rsp_thrown_payload_fragment_opcode;
  wire       [63:0]   io_output_rsp_thrown_payload_fragment_data;
  wire       [47:0]   io_output_rsp_thrown_payload_fragment_context;

  assign _zz_buffer_last_1 = 1'b1;
  assign _zz_buffer_last = {2'd0, _zz_buffer_last_1};
  assign _zz_buffer_addressIncr = (buffer_address[11 : 0] + 12'h008);
  assign buffer_last = (buffer_beat == _zz_buffer_last);
  assign buffer_addressIncr = {buffer_address[31 : 12],(_zz_buffer_addressIncr & (~ 12'h007))};
  assign buffer_isWrite = (buffer_opcode == 1'b1);
  assign io_output_cmd_fire = (io_output_cmd_valid && io_output_cmd_ready);
  assign cmdTransferBeatCount = io_input_cmd_payload_fragment_length[5 : 3];
  assign requireBuffer = (cmdTransferBeatCount != 3'b000);
  assign io_output_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_output_cmd_payload_last = 1'b1;
  assign io_output_cmd_payload_fragment_context = {cmdContext_context,{cmdContext_source,{cmdContext_last,cmdContext_drop}}};
  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_payload_fragment_address = buffer_addressIncr;
    end else begin
      io_output_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
      if(requireBuffer) begin
        io_output_cmd_payload_fragment_address[2 : 0] = 3'b000;
      end
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_payload_fragment_opcode = buffer_opcode;
    end else begin
      io_output_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_payload_fragment_length = 3'b111;
    end else begin
      if(requireBuffer) begin
        io_output_cmd_payload_fragment_length = 3'b111;
      end else begin
        io_output_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length[2:0];
      end
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_context = buffer_context;
    end else begin
      cmdContext_context = io_input_cmd_payload_fragment_context;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_source = buffer_source;
    end else begin
      cmdContext_source = io_input_cmd_payload_fragment_source;
    end
  end

  always @(*) begin
    io_input_cmd_ready = 1'b0;
    if(buffer_valid) begin
      io_input_cmd_ready = (buffer_isWrite && io_output_cmd_ready);
    end else begin
      io_input_cmd_ready = io_output_cmd_ready;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_valid = (! (buffer_isWrite && (! io_input_cmd_valid)));
    end else begin
      io_output_cmd_valid = io_input_cmd_valid;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_last = buffer_last;
    end else begin
      cmdContext_last = (! requireBuffer);
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_drop = buffer_isWrite;
    end else begin
      cmdContext_drop = (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
  end

  assign _zz_rspContext_drop = io_output_rsp_payload_fragment_context;
  assign rspContext_drop = _zz_rspContext_drop[0];
  assign rspContext_last = _zz_rspContext_drop[1];
  assign rspContext_source = _zz_rspContext_drop[3 : 2];
  assign rspContext_context = _zz_rspContext_drop[47 : 4];
  assign when_Stream_l445 = (! (rspContext_last || (! rspContext_drop)));
  always @(*) begin
    io_output_rsp_thrown_valid = io_output_rsp_valid;
    if(when_Stream_l445) begin
      io_output_rsp_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    io_output_rsp_ready = io_output_rsp_thrown_ready;
    if(when_Stream_l445) begin
      io_output_rsp_ready = 1'b1;
    end
  end

  assign io_output_rsp_thrown_payload_last = io_output_rsp_payload_last;
  assign io_output_rsp_thrown_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_output_rsp_thrown_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_output_rsp_thrown_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign io_input_rsp_valid = io_output_rsp_thrown_valid;
  assign io_output_rsp_thrown_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = rspContext_last;
  assign io_input_rsp_payload_fragment_source = rspContext_source;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = rspContext_context;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      buffer_valid <= 1'b0;
    end else begin
      if(io_output_cmd_fire) begin
        if(buffer_last) begin
          buffer_valid <= 1'b0;
        end
      end
      if(!buffer_valid) begin
        buffer_valid <= (requireBuffer && io_output_cmd_fire);
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_output_cmd_fire) begin
      buffer_beat <= (buffer_beat - 3'b001);
      buffer_address[11 : 0] <= buffer_addressIncr[11 : 0];
    end
    if(!buffer_valid) begin
      buffer_opcode <= io_input_cmd_payload_fragment_opcode;
      buffer_source <= io_input_cmd_payload_fragment_source;
      buffer_address <= io_input_cmd_payload_fragment_address;
      buffer_context <= io_input_cmd_payload_fragment_context;
      buffer_beat <= cmdTransferBeatCount;
    end
  end


endmodule

module BmbCcToggle (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [1:0]    io_input_cmd_payload_fragment_length,
  input  wire [31:0]   io_input_cmd_payload_fragment_data,
  input  wire [3:0]    io_input_cmd_payload_fragment_mask,
  input  wire [48:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [31:0]   io_input_rsp_payload_fragment_data,
  output wire [48:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [1:0]    io_output_cmd_payload_fragment_length,
  output wire [31:0]   io_output_cmd_payload_fragment_data,
  output wire [3:0]    io_output_cmd_payload_fragment_mask,
  output wire [48:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_output_rsp_payload_fragment_data,
  input  wire [48:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset,
  input  wire          io_peripheralClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1,
  input  wire          peripheralCd_logic_outputReset,
  input  wire          system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1
);

  wire                io_input_cmd_ccToggle_io_input_ready;
  wire                io_input_cmd_ccToggle_io_output_valid;
  wire                io_input_cmd_ccToggle_io_output_payload_last;
  wire       [0:0]    io_input_cmd_ccToggle_io_output_payload_fragment_opcode;
  wire       [31:0]   io_input_cmd_ccToggle_io_output_payload_fragment_address;
  wire       [1:0]    io_input_cmd_ccToggle_io_output_payload_fragment_length;
  wire       [31:0]   io_input_cmd_ccToggle_io_output_payload_fragment_data;
  wire       [3:0]    io_input_cmd_ccToggle_io_output_payload_fragment_mask;
  wire       [48:0]   io_input_cmd_ccToggle_io_output_payload_fragment_context;
  wire                io_output_rsp_ccToggle_io_input_ready;
  wire                io_output_rsp_ccToggle_io_output_valid;
  wire                io_output_rsp_ccToggle_io_output_payload_last;
  wire       [0:0]    io_output_rsp_ccToggle_io_output_payload_fragment_opcode;
  wire       [31:0]   io_output_rsp_ccToggle_io_output_payload_fragment_data;
  wire       [48:0]   io_output_rsp_ccToggle_io_output_payload_fragment_context;

  StreamCCByToggle io_input_cmd_ccToggle (
    .io_input_valid                                                                  (io_input_cmd_valid                                                             ), //i
    .io_input_ready                                                                  (io_input_cmd_ccToggle_io_input_ready                                           ), //o
    .io_input_payload_last                                                           (io_input_cmd_payload_last                                                      ), //i
    .io_input_payload_fragment_opcode                                                (io_input_cmd_payload_fragment_opcode                                           ), //i
    .io_input_payload_fragment_address                                               (io_input_cmd_payload_fragment_address[31:0]                                    ), //i
    .io_input_payload_fragment_length                                                (io_input_cmd_payload_fragment_length[1:0]                                      ), //i
    .io_input_payload_fragment_data                                                  (io_input_cmd_payload_fragment_data[31:0]                                       ), //i
    .io_input_payload_fragment_mask                                                  (io_input_cmd_payload_fragment_mask[3:0]                                        ), //i
    .io_input_payload_fragment_context                                               (io_input_cmd_payload_fragment_context[48:0]                                    ), //i
    .io_output_valid                                                                 (io_input_cmd_ccToggle_io_output_valid                                          ), //o
    .io_output_ready                                                                 (io_output_cmd_ready                                                            ), //i
    .io_output_payload_last                                                          (io_input_cmd_ccToggle_io_output_payload_last                                   ), //o
    .io_output_payload_fragment_opcode                                               (io_input_cmd_ccToggle_io_output_payload_fragment_opcode                        ), //o
    .io_output_payload_fragment_address                                              (io_input_cmd_ccToggle_io_output_payload_fragment_address[31:0]                 ), //o
    .io_output_payload_fragment_length                                               (io_input_cmd_ccToggle_io_output_payload_fragment_length[1:0]                   ), //o
    .io_output_payload_fragment_data                                                 (io_input_cmd_ccToggle_io_output_payload_fragment_data[31:0]                    ), //o
    .io_output_payload_fragment_mask                                                 (io_input_cmd_ccToggle_io_output_payload_fragment_mask[3:0]                     ), //o
    .io_output_payload_fragment_context                                              (io_input_cmd_ccToggle_io_output_payload_fragment_context[48:0]                 ), //o
    .io_systemClk                                                                    (io_systemClk                                                                   ), //i
    .systemCd_logic_outputReset                                                      (systemCd_logic_outputReset                                                     ), //i
    .io_peripheralClk                                                                (io_peripheralClk                                                               ), //i
    .system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1)  //i
  );
  StreamCCByToggle_1 io_output_rsp_ccToggle (
    .io_input_valid                                                                      (io_output_rsp_valid                                                                ), //i
    .io_input_ready                                                                      (io_output_rsp_ccToggle_io_input_ready                                              ), //o
    .io_input_payload_last                                                               (io_output_rsp_payload_last                                                         ), //i
    .io_input_payload_fragment_opcode                                                    (io_output_rsp_payload_fragment_opcode                                              ), //i
    .io_input_payload_fragment_data                                                      (io_output_rsp_payload_fragment_data[31:0]                                          ), //i
    .io_input_payload_fragment_context                                                   (io_output_rsp_payload_fragment_context[48:0]                                       ), //i
    .io_output_valid                                                                     (io_output_rsp_ccToggle_io_output_valid                                             ), //o
    .io_output_ready                                                                     (io_input_rsp_ready                                                                 ), //i
    .io_output_payload_last                                                              (io_output_rsp_ccToggle_io_output_payload_last                                      ), //o
    .io_output_payload_fragment_opcode                                                   (io_output_rsp_ccToggle_io_output_payload_fragment_opcode                           ), //o
    .io_output_payload_fragment_data                                                     (io_output_rsp_ccToggle_io_output_payload_fragment_data[31:0]                       ), //o
    .io_output_payload_fragment_context                                                  (io_output_rsp_ccToggle_io_output_payload_fragment_context[48:0]                    ), //o
    .io_peripheralClk                                                                    (io_peripheralClk                                                                   ), //i
    .peripheralCd_logic_outputReset                                                      (peripheralCd_logic_outputReset                                                     ), //i
    .io_systemClk                                                                        (io_systemClk                                                                       ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //i
  );
  assign io_input_cmd_ready = io_input_cmd_ccToggle_io_input_ready;
  assign io_output_cmd_valid = io_input_cmd_ccToggle_io_output_valid;
  assign io_output_cmd_payload_last = io_input_cmd_ccToggle_io_output_payload_last;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_ccToggle_io_output_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_ccToggle_io_output_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_ccToggle_io_output_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = io_input_cmd_ccToggle_io_output_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = io_input_cmd_ccToggle_io_output_payload_fragment_mask;
  assign io_output_cmd_payload_fragment_context = io_input_cmd_ccToggle_io_output_payload_fragment_context;
  assign io_output_rsp_ready = io_output_rsp_ccToggle_io_input_ready;
  assign io_input_rsp_valid = io_output_rsp_ccToggle_io_output_valid;
  assign io_input_rsp_payload_last = io_output_rsp_ccToggle_io_output_payload_last;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_ccToggle_io_output_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_ccToggle_io_output_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = io_output_rsp_ccToggle_io_output_payload_fragment_context;

endmodule

module BmbUnburstify (
  input  wire          io_input_cmd_valid,
  output reg           io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [31:0]   io_input_cmd_payload_fragment_data,
  input  wire [3:0]    io_input_cmd_payload_fragment_mask,
  input  wire [44:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [31:0]   io_input_rsp_payload_fragment_data,
  output wire [44:0]   io_input_rsp_payload_fragment_context,
  output reg           io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output reg  [0:0]    io_output_cmd_payload_fragment_opcode,
  output reg  [31:0]   io_output_cmd_payload_fragment_address,
  output reg  [1:0]    io_output_cmd_payload_fragment_length,
  output wire [31:0]   io_output_cmd_payload_fragment_data,
  output wire [3:0]    io_output_cmd_payload_fragment_mask,
  output wire [48:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output reg           io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_output_rsp_payload_fragment_data,
  input  wire [48:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [3:0]    _zz_buffer_last;
  wire       [0:0]    _zz_buffer_last_1;
  wire       [11:0]   _zz_buffer_addressIncr;
  wire                doResult;
  reg                 buffer_valid;
  reg        [0:0]    buffer_opcode;
  reg        [1:0]    buffer_source;
  reg        [31:0]   buffer_address;
  reg        [44:0]   buffer_context;
  reg        [3:0]    buffer_beat;
  wire                buffer_last;
  wire       [31:0]   buffer_addressIncr;
  wire                buffer_isWrite;
  wire                io_output_cmd_fire;
  wire       [3:0]    cmdTransferBeatCount;
  wire                requireBuffer;
  reg                 cmdContext_drop;
  reg                 cmdContext_last;
  reg        [1:0]    cmdContext_source;
  reg        [44:0]   cmdContext_context;
  wire                rspContext_drop;
  wire                rspContext_last;
  wire       [1:0]    rspContext_source;
  wire       [44:0]   rspContext_context;
  wire       [48:0]   _zz_rspContext_drop;
  wire                when_Stream_l445;
  reg                 io_output_rsp_thrown_valid;
  wire                io_output_rsp_thrown_ready;
  wire                io_output_rsp_thrown_payload_last;
  wire       [0:0]    io_output_rsp_thrown_payload_fragment_opcode;
  wire       [31:0]   io_output_rsp_thrown_payload_fragment_data;
  wire       [48:0]   io_output_rsp_thrown_payload_fragment_context;

  assign _zz_buffer_last_1 = 1'b1;
  assign _zz_buffer_last = {3'd0, _zz_buffer_last_1};
  assign _zz_buffer_addressIncr = (buffer_address[11 : 0] + 12'h004);
  assign buffer_last = (buffer_beat == _zz_buffer_last);
  assign buffer_addressIncr = {buffer_address[31 : 12],(_zz_buffer_addressIncr & (~ 12'h003))};
  assign buffer_isWrite = (buffer_opcode == 1'b1);
  assign io_output_cmd_fire = (io_output_cmd_valid && io_output_cmd_ready);
  assign cmdTransferBeatCount = io_input_cmd_payload_fragment_length[5 : 2];
  assign requireBuffer = (cmdTransferBeatCount != 4'b0000);
  assign io_output_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_output_cmd_payload_last = 1'b1;
  assign io_output_cmd_payload_fragment_context = {cmdContext_context,{cmdContext_source,{cmdContext_last,cmdContext_drop}}};
  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_payload_fragment_address = buffer_addressIncr;
    end else begin
      io_output_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
      if(requireBuffer) begin
        io_output_cmd_payload_fragment_address[1 : 0] = 2'b00;
      end
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_payload_fragment_opcode = buffer_opcode;
    end else begin
      io_output_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_payload_fragment_length = 2'b11;
    end else begin
      if(requireBuffer) begin
        io_output_cmd_payload_fragment_length = 2'b11;
      end else begin
        io_output_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length[1:0];
      end
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_context = buffer_context;
    end else begin
      cmdContext_context = io_input_cmd_payload_fragment_context;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_source = buffer_source;
    end else begin
      cmdContext_source = io_input_cmd_payload_fragment_source;
    end
  end

  always @(*) begin
    io_input_cmd_ready = 1'b0;
    if(buffer_valid) begin
      io_input_cmd_ready = (buffer_isWrite && io_output_cmd_ready);
    end else begin
      io_input_cmd_ready = io_output_cmd_ready;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      io_output_cmd_valid = (! (buffer_isWrite && (! io_input_cmd_valid)));
    end else begin
      io_output_cmd_valid = io_input_cmd_valid;
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_last = buffer_last;
    end else begin
      cmdContext_last = (! requireBuffer);
    end
  end

  always @(*) begin
    if(buffer_valid) begin
      cmdContext_drop = buffer_isWrite;
    end else begin
      cmdContext_drop = (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
  end

  assign _zz_rspContext_drop = io_output_rsp_payload_fragment_context;
  assign rspContext_drop = _zz_rspContext_drop[0];
  assign rspContext_last = _zz_rspContext_drop[1];
  assign rspContext_source = _zz_rspContext_drop[3 : 2];
  assign rspContext_context = _zz_rspContext_drop[48 : 4];
  assign when_Stream_l445 = (! (rspContext_last || (! rspContext_drop)));
  always @(*) begin
    io_output_rsp_thrown_valid = io_output_rsp_valid;
    if(when_Stream_l445) begin
      io_output_rsp_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    io_output_rsp_ready = io_output_rsp_thrown_ready;
    if(when_Stream_l445) begin
      io_output_rsp_ready = 1'b1;
    end
  end

  assign io_output_rsp_thrown_payload_last = io_output_rsp_payload_last;
  assign io_output_rsp_thrown_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_output_rsp_thrown_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_output_rsp_thrown_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign io_input_rsp_valid = io_output_rsp_thrown_valid;
  assign io_output_rsp_thrown_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = rspContext_last;
  assign io_input_rsp_payload_fragment_source = rspContext_source;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = rspContext_context;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      buffer_valid <= 1'b0;
    end else begin
      if(io_output_cmd_fire) begin
        if(buffer_last) begin
          buffer_valid <= 1'b0;
        end
      end
      if(!buffer_valid) begin
        buffer_valid <= (requireBuffer && io_output_cmd_fire);
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_output_cmd_fire) begin
      buffer_beat <= (buffer_beat - 4'b0001);
      buffer_address[11 : 0] <= buffer_addressIncr[11 : 0];
    end
    if(!buffer_valid) begin
      buffer_opcode <= io_input_cmd_payload_fragment_opcode;
      buffer_source <= io_input_cmd_payload_fragment_source;
      buffer_address <= io_input_cmd_payload_fragment_address;
      buffer_context <= io_input_cmd_payload_fragment_context;
      buffer_beat <= cmdTransferBeatCount;
    end
  end


endmodule

//BmbDownSizerBridge_1 replaced by BmbDownSizerBridge

module BmbOnChipRam (
  input  wire          io_bus_cmd_valid,
  output wire          io_bus_cmd_ready,
  input  wire          io_bus_cmd_payload_last,
  input  wire [0:0]    io_bus_cmd_payload_fragment_opcode,
  input  wire [10:0]   io_bus_cmd_payload_fragment_address,
  input  wire [2:0]    io_bus_cmd_payload_fragment_length,
  input  wire [63:0]   io_bus_cmd_payload_fragment_data,
  input  wire [7:0]    io_bus_cmd_payload_fragment_mask,
  input  wire [47:0]   io_bus_cmd_payload_fragment_context,
  output wire          io_bus_rsp_valid,
  input  wire          io_bus_rsp_ready,
  output wire          io_bus_rsp_payload_last,
  output wire [0:0]    io_bus_rsp_payload_fragment_opcode,
  output wire [63:0]   io_bus_rsp_payload_fragment_data,
  output wire [47:0]   io_bus_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg        [63:0]   ram_spinal_port0;
  wire                enabled;
  wire                io_bus_rsp_isStall;
  reg                 io_bus_cmd_valid_regNextWhen;
  reg        [47:0]   io_bus_cmd_payload_fragment_context_regNextWhen;
  wire       [7:0]    address;
  wire       [63:0]   data;
  wire                io_bus_cmd_fire;
  wire                enable;
  wire                write;
  wire       [7:0]    mask;
  wire       [63:0]   _zz_io_bus_rsp_payload_fragment_data;
  reg [7:0] ram_symbol0 [0:255];
  reg [7:0] ram_symbol1 [0:255];
  reg [7:0] ram_symbol2 [0:255];
  reg [7:0] ram_symbol3 [0:255];
  reg [7:0] ram_symbol4 [0:255];
  reg [7:0] ram_symbol5 [0:255];
  reg [7:0] ram_symbol6 [0:255];
  reg [7:0] ram_symbol7 [0:255];
  reg [7:0] _zz_ramsymbol_read;
  reg [7:0] _zz_ramsymbol_read_1;
  reg [7:0] _zz_ramsymbol_read_2;
  reg [7:0] _zz_ramsymbol_read_3;
  reg [7:0] _zz_ramsymbol_read_4;
  reg [7:0] _zz_ramsymbol_read_5;
  reg [7:0] _zz_ramsymbol_read_6;
  reg [7:0] _zz_ramsymbol_read_7;

  initial begin
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol0.bin",ram_symbol0);
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol1.bin",ram_symbol1);
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol2.bin",ram_symbol2);
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol3.bin",ram_symbol3);
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol4.bin",ram_symbol4);
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol5.bin",ram_symbol5);
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol6.bin",ram_symbol6);
    $readmemb("EfxSapphireSoc.v_toplevel_system_ramA_logic_ram_symbol7.bin",ram_symbol7);
  end
  always @(*) begin
    ram_spinal_port0 = {_zz_ramsymbol_read_7, _zz_ramsymbol_read_6, _zz_ramsymbol_read_5, _zz_ramsymbol_read_4, _zz_ramsymbol_read_3, _zz_ramsymbol_read_2, _zz_ramsymbol_read_1, _zz_ramsymbol_read};
  end
  always @(posedge io_systemClk) begin
    if(enable) begin
      _zz_ramsymbol_read <= ram_symbol0[address];
      _zz_ramsymbol_read_1 <= ram_symbol1[address];
      _zz_ramsymbol_read_2 <= ram_symbol2[address];
      _zz_ramsymbol_read_3 <= ram_symbol3[address];
      _zz_ramsymbol_read_4 <= ram_symbol4[address];
      _zz_ramsymbol_read_5 <= ram_symbol5[address];
      _zz_ramsymbol_read_6 <= ram_symbol6[address];
      _zz_ramsymbol_read_7 <= ram_symbol7[address];
    end
  end

  always @(posedge io_systemClk) begin
    if(mask[0] && enable && write ) begin
      ram_symbol0[address] <= _zz_io_bus_rsp_payload_fragment_data[7 : 0];
    end
    if(mask[1] && enable && write ) begin
      ram_symbol1[address] <= _zz_io_bus_rsp_payload_fragment_data[15 : 8];
    end
    if(mask[2] && enable && write ) begin
      ram_symbol2[address] <= _zz_io_bus_rsp_payload_fragment_data[23 : 16];
    end
    if(mask[3] && enable && write ) begin
      ram_symbol3[address] <= _zz_io_bus_rsp_payload_fragment_data[31 : 24];
    end
    if(mask[4] && enable && write ) begin
      ram_symbol4[address] <= _zz_io_bus_rsp_payload_fragment_data[39 : 32];
    end
    if(mask[5] && enable && write ) begin
      ram_symbol5[address] <= _zz_io_bus_rsp_payload_fragment_data[47 : 40];
    end
    if(mask[6] && enable && write ) begin
      ram_symbol6[address] <= _zz_io_bus_rsp_payload_fragment_data[55 : 48];
    end
    if(mask[7] && enable && write ) begin
      ram_symbol7[address] <= _zz_io_bus_rsp_payload_fragment_data[63 : 56];
    end
  end

  assign enabled = 1'b1;
  assign io_bus_rsp_isStall = (io_bus_rsp_valid && (! io_bus_rsp_ready));
  assign io_bus_cmd_ready = (! io_bus_rsp_isStall);
  assign io_bus_rsp_valid = io_bus_cmd_valid_regNextWhen;
  assign io_bus_rsp_payload_fragment_context = io_bus_cmd_payload_fragment_context_regNextWhen;
  assign address = (io_bus_cmd_payload_fragment_address >>> 2'd3);
  assign data = io_bus_cmd_payload_fragment_data;
  assign io_bus_cmd_fire = (io_bus_cmd_valid && io_bus_cmd_ready);
  assign enable = (io_bus_cmd_fire && enabled);
  assign write = (io_bus_cmd_payload_fragment_opcode == 1'b1);
  assign mask = io_bus_cmd_payload_fragment_mask;
  assign _zz_io_bus_rsp_payload_fragment_data = data;
  assign io_bus_rsp_payload_fragment_data = ram_spinal_port0;
  assign io_bus_rsp_payload_fragment_opcode = 1'b0;
  assign io_bus_rsp_payload_last = 1'b1;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      io_bus_cmd_valid_regNextWhen <= 1'b0;
    end else begin
      if(io_bus_cmd_ready) begin
        io_bus_cmd_valid_regNextWhen <= io_bus_cmd_valid;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_bus_cmd_ready) begin
      io_bus_cmd_payload_fragment_context_regNextWhen <= io_bus_cmd_payload_fragment_context;
    end
  end


endmodule

module BmbCcFifo_1 (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [31:0]   io_input_cmd_payload_fragment_data,
  input  wire [3:0]    io_input_cmd_payload_fragment_mask,
  input  wire [44:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [31:0]   io_input_rsp_payload_fragment_data,
  output wire [44:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [1:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output wire [31:0]   io_output_cmd_payload_fragment_data,
  output wire [3:0]    io_output_cmd_payload_fragment_mask,
  output wire [44:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [1:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_output_rsp_payload_fragment_data,
  input  wire [44:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset,
  output wire          system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1,
  output wire          system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1
);

  wire                io_input_cmd_queue_io_push_ready;
  wire                io_input_cmd_queue_io_pop_valid;
  wire                io_input_cmd_queue_io_pop_payload_last;
  wire       [1:0]    io_input_cmd_queue_io_pop_payload_fragment_source;
  wire       [0:0]    io_input_cmd_queue_io_pop_payload_fragment_opcode;
  wire       [31:0]   io_input_cmd_queue_io_pop_payload_fragment_address;
  wire       [5:0]    io_input_cmd_queue_io_pop_payload_fragment_length;
  wire       [31:0]   io_input_cmd_queue_io_pop_payload_fragment_data;
  wire       [3:0]    io_input_cmd_queue_io_pop_payload_fragment_mask;
  wire       [44:0]   io_input_cmd_queue_io_pop_payload_fragment_context;
  wire       [4:0]    io_input_cmd_queue_io_pushOccupancy;
  wire       [4:0]    io_input_cmd_queue_io_popOccupancy;
  wire                io_input_cmd_queue_system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1;
  wire                io_output_rsp_queue_io_push_ready;
  wire                io_output_rsp_queue_io_pop_valid;
  wire                io_output_rsp_queue_io_pop_payload_last;
  wire       [1:0]    io_output_rsp_queue_io_pop_payload_fragment_source;
  wire       [0:0]    io_output_rsp_queue_io_pop_payload_fragment_opcode;
  wire       [31:0]   io_output_rsp_queue_io_pop_payload_fragment_data;
  wire       [44:0]   io_output_rsp_queue_io_pop_payload_fragment_context;
  wire       [4:0]    io_output_rsp_queue_io_pushOccupancy;
  wire       [4:0]    io_output_rsp_queue_io_popOccupancy;
  wire                io_output_rsp_queue_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1;

  StreamFifoCC_12 io_input_cmd_queue (
    .io_push_valid                                                                   (io_input_cmd_valid                                                                                ), //i
    .io_push_ready                                                                   (io_input_cmd_queue_io_push_ready                                                                  ), //o
    .io_push_payload_last                                                            (io_input_cmd_payload_last                                                                         ), //i
    .io_push_payload_fragment_source                                                 (io_input_cmd_payload_fragment_source[1:0]                                                         ), //i
    .io_push_payload_fragment_opcode                                                 (io_input_cmd_payload_fragment_opcode                                                              ), //i
    .io_push_payload_fragment_address                                                (io_input_cmd_payload_fragment_address[31:0]                                                       ), //i
    .io_push_payload_fragment_length                                                 (io_input_cmd_payload_fragment_length[5:0]                                                         ), //i
    .io_push_payload_fragment_data                                                   (io_input_cmd_payload_fragment_data[31:0]                                                          ), //i
    .io_push_payload_fragment_mask                                                   (io_input_cmd_payload_fragment_mask[3:0]                                                           ), //i
    .io_push_payload_fragment_context                                                (io_input_cmd_payload_fragment_context[44:0]                                                       ), //i
    .io_pop_valid                                                                    (io_input_cmd_queue_io_pop_valid                                                                   ), //o
    .io_pop_ready                                                                    (io_output_cmd_ready                                                                               ), //i
    .io_pop_payload_last                                                             (io_input_cmd_queue_io_pop_payload_last                                                            ), //o
    .io_pop_payload_fragment_source                                                  (io_input_cmd_queue_io_pop_payload_fragment_source[1:0]                                            ), //o
    .io_pop_payload_fragment_opcode                                                  (io_input_cmd_queue_io_pop_payload_fragment_opcode                                                 ), //o
    .io_pop_payload_fragment_address                                                 (io_input_cmd_queue_io_pop_payload_fragment_address[31:0]                                          ), //o
    .io_pop_payload_fragment_length                                                  (io_input_cmd_queue_io_pop_payload_fragment_length[5:0]                                            ), //o
    .io_pop_payload_fragment_data                                                    (io_input_cmd_queue_io_pop_payload_fragment_data[31:0]                                             ), //o
    .io_pop_payload_fragment_mask                                                    (io_input_cmd_queue_io_pop_payload_fragment_mask[3:0]                                              ), //o
    .io_pop_payload_fragment_context                                                 (io_input_cmd_queue_io_pop_payload_fragment_context[44:0]                                          ), //o
    .io_pushOccupancy                                                                (io_input_cmd_queue_io_pushOccupancy[4:0]                                                          ), //o
    .io_popOccupancy                                                                 (io_input_cmd_queue_io_popOccupancy[4:0]                                                           ), //o
    .io_systemClk                                                                    (io_systemClk                                                                                      ), //i
    .systemCd_logic_outputReset                                                      (systemCd_logic_outputReset                                                                        ), //i
    .io_peripheralClk                                                                (io_peripheralClk                                                                                  ), //i
    .system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1 (io_input_cmd_queue_system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1)  //o
  );
  StreamFifoCC_13 io_output_rsp_queue (
    .io_push_valid                                                                       (io_output_rsp_valid                                                                                    ), //i
    .io_push_ready                                                                       (io_output_rsp_queue_io_push_ready                                                                      ), //o
    .io_push_payload_last                                                                (io_output_rsp_payload_last                                                                             ), //i
    .io_push_payload_fragment_source                                                     (io_output_rsp_payload_fragment_source[1:0]                                                             ), //i
    .io_push_payload_fragment_opcode                                                     (io_output_rsp_payload_fragment_opcode                                                                  ), //i
    .io_push_payload_fragment_data                                                       (io_output_rsp_payload_fragment_data[31:0]                                                              ), //i
    .io_push_payload_fragment_context                                                    (io_output_rsp_payload_fragment_context[44:0]                                                           ), //i
    .io_pop_valid                                                                        (io_output_rsp_queue_io_pop_valid                                                                       ), //o
    .io_pop_ready                                                                        (io_input_rsp_ready                                                                                     ), //i
    .io_pop_payload_last                                                                 (io_output_rsp_queue_io_pop_payload_last                                                                ), //o
    .io_pop_payload_fragment_source                                                      (io_output_rsp_queue_io_pop_payload_fragment_source[1:0]                                                ), //o
    .io_pop_payload_fragment_opcode                                                      (io_output_rsp_queue_io_pop_payload_fragment_opcode                                                     ), //o
    .io_pop_payload_fragment_data                                                        (io_output_rsp_queue_io_pop_payload_fragment_data[31:0]                                                 ), //o
    .io_pop_payload_fragment_context                                                     (io_output_rsp_queue_io_pop_payload_fragment_context[44:0]                                              ), //o
    .io_pushOccupancy                                                                    (io_output_rsp_queue_io_pushOccupancy[4:0]                                                              ), //o
    .io_popOccupancy                                                                     (io_output_rsp_queue_io_popOccupancy[4:0]                                                               ), //o
    .io_peripheralClk                                                                    (io_peripheralClk                                                                                       ), //i
    .peripheralCd_logic_outputReset                                                      (peripheralCd_logic_outputReset                                                                         ), //i
    .io_systemClk                                                                        (io_systemClk                                                                                           ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (io_output_rsp_queue_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //o
  );
  assign io_input_cmd_ready = io_input_cmd_queue_io_push_ready;
  assign io_output_cmd_valid = io_input_cmd_queue_io_pop_valid;
  assign io_output_cmd_payload_last = io_input_cmd_queue_io_pop_payload_last;
  assign io_output_cmd_payload_fragment_source = io_input_cmd_queue_io_pop_payload_fragment_source;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_queue_io_pop_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_queue_io_pop_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_queue_io_pop_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = io_input_cmd_queue_io_pop_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = io_input_cmd_queue_io_pop_payload_fragment_mask;
  assign io_output_cmd_payload_fragment_context = io_input_cmd_queue_io_pop_payload_fragment_context;
  assign io_output_rsp_ready = io_output_rsp_queue_io_push_ready;
  assign io_input_rsp_valid = io_output_rsp_queue_io_pop_valid;
  assign io_input_rsp_payload_last = io_output_rsp_queue_io_pop_payload_last;
  assign io_input_rsp_payload_fragment_source = io_output_rsp_queue_io_pop_payload_fragment_source;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_queue_io_pop_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_queue_io_pop_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = io_output_rsp_queue_io_pop_payload_fragment_context;
  assign system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1 = io_input_cmd_queue_system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1;
  assign system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 = io_output_rsp_queue_system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1;

endmodule

module BmbDownSizerBridge (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [63:0]   io_input_cmd_payload_fragment_data,
  input  wire [7:0]    io_input_cmd_payload_fragment_mask,
  input  wire [43:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire [43:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [1:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output wire [31:0]   io_output_cmd_payload_fragment_data,
  output wire [3:0]    io_output_cmd_payload_fragment_mask,
  output wire [44:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output reg           io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [1:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [31:0]   io_output_rsp_payload_fragment_data,
  input  wire [44:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg        [31:0]   _zz_io_output_cmd_payload_fragment_data;
  reg        [3:0]    _zz_io_output_cmd_payload_fragment_mask;
  wire       [31:0]   _zz_io_output_cmd_payload_last;
  wire       [31:0]   _zz_io_output_cmd_payload_last_1;
  wire       [0:0]    cmdArea_context_sel;
  wire       [43:0]   cmdArea_context_context;
  wire                io_output_cmd_fire;
  reg                 cmdArea_writeLogic_locked;
  reg        [0:0]    cmdArea_writeLogic_counter;
  wire       [0:0]    cmdArea_writeLogic_sel;
  wire       [0:0]    rspArea_context_sel;
  wire       [43:0]   rspArea_context_context;
  wire       [44:0]   _zz_rspArea_context_sel;
  wire                io_output_rsp_fire;
  reg                 rspArea_readLogic_locked;
  reg        [0:0]    rspArea_readLogic_counter;
  wire       [0:0]    rspArea_readLogic_sel;
  reg        [31:0]   rspArea_readLogic_buffers_0;
  reg        [31:0]   rspArea_readLogic_words_0;
  wire       [31:0]   rspArea_readLogic_words_1;
  wire                when_BmbDownSizerBridge_l97;
  wire                when_BmbDownSizerBridge_l106;
  wire                when_BmbDownSizerBridge_l114;

  assign _zz_io_output_cmd_payload_last = (io_input_cmd_payload_fragment_address + _zz_io_output_cmd_payload_last_1);
  assign _zz_io_output_cmd_payload_last_1 = {26'd0, io_input_cmd_payload_fragment_length};
  always @(*) begin
    case(cmdArea_writeLogic_sel)
      1'b0 : begin
        _zz_io_output_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data[31 : 0];
        _zz_io_output_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask[3 : 0];
      end
      default : begin
        _zz_io_output_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data[63 : 32];
        _zz_io_output_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask[7 : 4];
      end
    endcase
  end

  assign cmdArea_context_context = io_input_cmd_payload_fragment_context;
  assign cmdArea_context_sel = io_input_cmd_payload_fragment_address[2 : 2];
  assign io_output_cmd_valid = io_input_cmd_valid;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_output_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_output_cmd_payload_fragment_context = {cmdArea_context_context,cmdArea_context_sel};
  assign io_output_cmd_fire = (io_output_cmd_valid && io_output_cmd_ready);
  assign cmdArea_writeLogic_sel = (cmdArea_writeLogic_locked ? cmdArea_writeLogic_counter : io_input_cmd_payload_fragment_address[2 : 2]);
  assign io_output_cmd_payload_fragment_data = _zz_io_output_cmd_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = _zz_io_output_cmd_payload_fragment_mask;
  assign io_output_cmd_payload_last = (io_input_cmd_payload_last && ((io_input_cmd_payload_fragment_opcode == 1'b0) || (cmdArea_writeLogic_sel == _zz_io_output_cmd_payload_last[2 : 2])));
  assign io_input_cmd_ready = (io_output_cmd_ready && ((cmdArea_writeLogic_sel == 1'b1) || io_output_cmd_payload_last));
  assign _zz_rspArea_context_sel = io_output_rsp_payload_fragment_context;
  assign rspArea_context_sel = _zz_rspArea_context_sel[0 : 0];
  assign rspArea_context_context = _zz_rspArea_context_sel[44 : 1];
  assign io_input_rsp_payload_last = io_output_rsp_payload_last;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_source = io_output_rsp_payload_fragment_source;
  assign io_input_rsp_payload_fragment_context = rspArea_context_context;
  always @(*) begin
    io_output_rsp_ready = io_input_rsp_ready;
    if(when_BmbDownSizerBridge_l114) begin
      io_output_rsp_ready = 1'b1;
    end
  end

  assign io_output_rsp_fire = (io_output_rsp_valid && io_output_rsp_ready);
  assign rspArea_readLogic_sel = (rspArea_readLogic_locked ? rspArea_readLogic_counter : rspArea_context_sel);
  assign when_BmbDownSizerBridge_l97 = (rspArea_readLogic_sel == 1'b0);
  always @(*) begin
    rspArea_readLogic_words_0 = rspArea_readLogic_buffers_0;
    if(when_BmbDownSizerBridge_l106) begin
      rspArea_readLogic_words_0 = io_output_rsp_payload_fragment_data;
    end
  end

  assign when_BmbDownSizerBridge_l106 = (io_input_rsp_payload_last && (rspArea_readLogic_sel == 1'b0));
  assign rspArea_readLogic_words_1 = io_output_rsp_payload_fragment_data;
  assign io_input_rsp_valid = (io_output_rsp_valid && (io_output_rsp_payload_last || (rspArea_readLogic_sel == 1'b1)));
  assign io_input_rsp_payload_fragment_data = {rspArea_readLogic_words_1,rspArea_readLogic_words_0};
  assign when_BmbDownSizerBridge_l114 = (! io_input_rsp_valid);
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      cmdArea_writeLogic_locked <= 1'b0;
      rspArea_readLogic_locked <= 1'b0;
    end else begin
      if(io_output_cmd_fire) begin
        cmdArea_writeLogic_locked <= (! io_output_cmd_payload_last);
      end
      if(io_output_rsp_fire) begin
        rspArea_readLogic_locked <= (! io_output_rsp_payload_last);
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_output_cmd_fire) begin
      cmdArea_writeLogic_counter <= (cmdArea_writeLogic_sel + 1'b1);
    end
    if(io_output_rsp_fire) begin
      rspArea_readLogic_counter <= (rspArea_readLogic_sel + 1'b1);
      if(when_BmbDownSizerBridge_l97) begin
        rspArea_readLogic_buffers_0 <= io_output_rsp_payload_fragment_data;
      end
    end
  end


endmodule

module BmbUpSizerBridge (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [63:0]   io_input_cmd_payload_fragment_data,
  input  wire [7:0]    io_input_cmd_payload_fragment_mask,
  input  wire [43:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output reg           io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire [43:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [1:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output reg  [127:0]  io_output_cmd_payload_fragment_data,
  output reg  [15:0]   io_output_cmd_payload_fragment_mask,
  output wire [45:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [1:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [127:0]  io_output_rsp_payload_fragment_data,
  input  wire [45:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [2:0]    _zz_cmdArea_context_selEnd;
  wire       [2:0]    _zz_cmdArea_context_selEnd_1;
  wire       [0:0]    _zz_cmdArea_context_selEnd_2;
  reg        [63:0]   _zz_io_input_rsp_payload_fragment_data;
  wire       [0:0]    cmdArea_selStart;
  wire       [0:0]    cmdArea_context_selStart;
  reg        [0:0]    cmdArea_context_selEnd;
  wire       [43:0]   cmdArea_context_context;
  wire                when_BmbUpSizerBridge_l53;
  reg        [63:0]   cmdArea_writeLogic_dataRegs_0;
  reg        [7:0]    cmdArea_writeLogic_maskRegs_0;
  reg        [0:0]    cmdArea_writeLogic_selReg;
  wire                io_input_cmd_fire;
  reg                 io_input_cmd_payload_first;
  wire       [0:0]    cmdArea_writeLogic_sel;
  wire       [63:0]   cmdArea_writeLogic_outputData_0;
  wire       [63:0]   cmdArea_writeLogic_outputData_1;
  wire       [7:0]    cmdArea_writeLogic_outputMask_0;
  wire       [7:0]    cmdArea_writeLogic_outputMask_1;
  wire                when_BmbUpSizerBridge_l85;
  wire                when_BmbUpSizerBridge_l95;
  wire                io_output_cmd_fire;
  wire                io_output_cmd_isStall;
  wire       [0:0]    rspArea_context_selStart;
  wire       [0:0]    rspArea_context_selEnd;
  wire       [43:0]   rspArea_context_context;
  wire       [45:0]   _zz_rspArea_context_selStart;
  reg        [0:0]    rspArea_readLogic_selReg;
  wire                io_input_rsp_fire;
  reg                 io_input_rsp_payload_first;
  wire       [0:0]    rspArea_readLogic_sel;
  wire                when_BmbUpSizerBridge_l133;

  assign _zz_cmdArea_context_selEnd = (_zz_cmdArea_context_selEnd_1 + io_input_cmd_payload_fragment_length[5 : 3]);
  assign _zz_cmdArea_context_selEnd_2 = io_input_cmd_payload_fragment_address[3 : 3];
  assign _zz_cmdArea_context_selEnd_1 = {2'd0, _zz_cmdArea_context_selEnd_2};
  always @(*) begin
    case(rspArea_readLogic_sel)
      1'b0 : _zz_io_input_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data[63 : 0];
      default : _zz_io_input_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data[127 : 64];
    endcase
  end

  assign cmdArea_selStart = io_input_cmd_payload_fragment_address[3 : 3];
  assign cmdArea_context_context = io_input_cmd_payload_fragment_context;
  assign cmdArea_context_selStart = cmdArea_selStart;
  always @(*) begin
    cmdArea_context_selEnd = _zz_cmdArea_context_selEnd[0:0];
    if(when_BmbUpSizerBridge_l53) begin
      cmdArea_context_selEnd = io_input_cmd_payload_fragment_address[3 : 3];
    end
  end

  assign when_BmbUpSizerBridge_l53 = (io_input_cmd_payload_fragment_opcode == 1'b1);
  assign io_output_cmd_payload_last = io_input_cmd_payload_last;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_output_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_output_cmd_payload_fragment_context = {cmdArea_context_context,{cmdArea_context_selEnd,cmdArea_context_selStart}};
  assign io_input_cmd_fire = (io_input_cmd_valid && io_input_cmd_ready);
  assign cmdArea_writeLogic_sel = (io_input_cmd_payload_first ? cmdArea_selStart : cmdArea_writeLogic_selReg);
  assign cmdArea_writeLogic_outputData_0 = io_output_cmd_payload_fragment_data[63 : 0];
  assign cmdArea_writeLogic_outputData_1 = io_output_cmd_payload_fragment_data[127 : 64];
  assign cmdArea_writeLogic_outputMask_0 = io_output_cmd_payload_fragment_mask[7 : 0];
  assign cmdArea_writeLogic_outputMask_1 = io_output_cmd_payload_fragment_mask[15 : 8];
  always @(*) begin
    io_output_cmd_payload_fragment_data[63 : 0] = io_input_cmd_payload_fragment_data;
    if(when_BmbUpSizerBridge_l85) begin
      io_output_cmd_payload_fragment_data[63 : 0] = cmdArea_writeLogic_dataRegs_0;
    end
    io_output_cmd_payload_fragment_data[127 : 64] = io_input_cmd_payload_fragment_data;
  end

  assign when_BmbUpSizerBridge_l85 = ((! io_input_cmd_payload_first) && (cmdArea_writeLogic_selReg != 1'b0));
  always @(*) begin
    io_output_cmd_payload_fragment_mask[7 : 0] = ((cmdArea_writeLogic_sel == 1'b0) ? io_input_cmd_payload_fragment_mask : cmdArea_writeLogic_maskRegs_0);
    io_output_cmd_payload_fragment_mask[15 : 8] = ((cmdArea_writeLogic_sel == 1'b1) ? io_input_cmd_payload_fragment_mask : 8'h0);
  end

  assign when_BmbUpSizerBridge_l95 = (io_input_cmd_valid && (cmdArea_writeLogic_sel == 1'b0));
  assign io_output_cmd_fire = (io_output_cmd_valid && io_output_cmd_ready);
  assign io_output_cmd_valid = (io_input_cmd_valid && ((cmdArea_writeLogic_sel == 1'b1) || io_input_cmd_payload_last));
  assign io_output_cmd_isStall = (io_output_cmd_valid && (! io_output_cmd_ready));
  assign io_input_cmd_ready = (! io_output_cmd_isStall);
  assign _zz_rspArea_context_selStart = io_output_rsp_payload_fragment_context;
  assign rspArea_context_selStart = _zz_rspArea_context_selStart[0 : 0];
  assign rspArea_context_selEnd = _zz_rspArea_context_selStart[1 : 1];
  assign rspArea_context_context = _zz_rspArea_context_selStart[45 : 2];
  assign io_input_rsp_valid = io_output_rsp_valid;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_source = io_output_rsp_payload_fragment_source;
  assign io_input_rsp_payload_fragment_context = rspArea_context_context;
  assign io_input_rsp_fire = (io_input_rsp_valid && io_input_rsp_ready);
  assign rspArea_readLogic_sel = (io_input_rsp_payload_first ? rspArea_context_selStart : rspArea_readLogic_selReg);
  always @(*) begin
    io_input_rsp_payload_last = (io_output_rsp_payload_last && (rspArea_readLogic_sel == rspArea_context_selEnd));
    if(when_BmbUpSizerBridge_l133) begin
      io_input_rsp_payload_last = 1'b0;
    end
  end

  assign io_output_rsp_ready = (io_input_rsp_ready && (io_input_rsp_payload_last || (rspArea_readLogic_sel == 1'b1)));
  assign when_BmbUpSizerBridge_l133 = (rspArea_context_selEnd != rspArea_readLogic_sel);
  assign io_input_rsp_payload_fragment_data = _zz_io_input_rsp_payload_fragment_data;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      cmdArea_writeLogic_maskRegs_0 <= 8'h0;
      io_input_cmd_payload_first <= 1'b1;
      io_input_rsp_payload_first <= 1'b1;
    end else begin
      if(io_input_cmd_fire) begin
        io_input_cmd_payload_first <= io_input_cmd_payload_last;
      end
      if(when_BmbUpSizerBridge_l95) begin
        cmdArea_writeLogic_maskRegs_0 <= io_input_cmd_payload_fragment_mask;
      end
      if(io_output_cmd_fire) begin
        cmdArea_writeLogic_maskRegs_0 <= 8'h0;
      end
      if(io_input_rsp_fire) begin
        io_input_rsp_payload_first <= io_input_rsp_payload_last;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_input_cmd_fire) begin
      cmdArea_writeLogic_selReg <= (cmdArea_writeLogic_sel + 1'b1);
    end
    if(!when_BmbUpSizerBridge_l85) begin
      cmdArea_writeLogic_dataRegs_0 <= io_input_cmd_payload_fragment_data;
    end
    rspArea_readLogic_selReg <= rspArea_readLogic_sel;
    if(io_input_rsp_fire) begin
      rspArea_readLogic_selReg <= (rspArea_readLogic_sel + 1'b1);
    end
  end


endmodule

module BmbDecoderPerSource (
  input  wire          io_input_cmd_valid,
  output reg           io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [63:0]   io_input_cmd_payload_fragment_data,
  input  wire [7:0]    io_input_cmd_payload_fragment_mask,
  input  wire [43:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire [43:0]   io_input_rsp_payload_fragment_context,
  output reg           io_outputs_0_cmd_valid,
  input  wire          io_outputs_0_cmd_ready,
  output wire          io_outputs_0_cmd_payload_last,
  output wire [1:0]    io_outputs_0_cmd_payload_fragment_source,
  output wire [0:0]    io_outputs_0_cmd_payload_fragment_opcode,
  output wire [31:0]   io_outputs_0_cmd_payload_fragment_address,
  output wire [5:0]    io_outputs_0_cmd_payload_fragment_length,
  output wire [63:0]   io_outputs_0_cmd_payload_fragment_data,
  output wire [7:0]    io_outputs_0_cmd_payload_fragment_mask,
  output wire [43:0]   io_outputs_0_cmd_payload_fragment_context,
  input  wire          io_outputs_0_rsp_valid,
  output wire          io_outputs_0_rsp_ready,
  input  wire          io_outputs_0_rsp_payload_last,
  input  wire [1:0]    io_outputs_0_rsp_payload_fragment_source,
  input  wire [0:0]    io_outputs_0_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_outputs_0_rsp_payload_fragment_data,
  input  wire [43:0]   io_outputs_0_rsp_payload_fragment_context,
  output reg           io_outputs_1_cmd_valid,
  input  wire          io_outputs_1_cmd_ready,
  output wire          io_outputs_1_cmd_payload_last,
  output wire [1:0]    io_outputs_1_cmd_payload_fragment_source,
  output wire [0:0]    io_outputs_1_cmd_payload_fragment_opcode,
  output wire [31:0]   io_outputs_1_cmd_payload_fragment_address,
  output wire [5:0]    io_outputs_1_cmd_payload_fragment_length,
  output wire [63:0]   io_outputs_1_cmd_payload_fragment_data,
  output wire [7:0]    io_outputs_1_cmd_payload_fragment_mask,
  output wire [43:0]   io_outputs_1_cmd_payload_fragment_context,
  input  wire          io_outputs_1_rsp_valid,
  output wire          io_outputs_1_rsp_ready,
  input  wire          io_outputs_1_rsp_payload_last,
  input  wire [1:0]    io_outputs_1_rsp_payload_fragment_source,
  input  wire [0:0]    io_outputs_1_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_outputs_1_rsp_payload_fragment_data,
  input  wire [43:0]   io_outputs_1_rsp_payload_fragment_context,
  output reg           io_outputs_2_cmd_valid,
  input  wire          io_outputs_2_cmd_ready,
  output wire          io_outputs_2_cmd_payload_last,
  output wire [1:0]    io_outputs_2_cmd_payload_fragment_source,
  output wire [0:0]    io_outputs_2_cmd_payload_fragment_opcode,
  output wire [31:0]   io_outputs_2_cmd_payload_fragment_address,
  output wire [5:0]    io_outputs_2_cmd_payload_fragment_length,
  output wire [63:0]   io_outputs_2_cmd_payload_fragment_data,
  output wire [7:0]    io_outputs_2_cmd_payload_fragment_mask,
  output wire [43:0]   io_outputs_2_cmd_payload_fragment_context,
  input  wire          io_outputs_2_rsp_valid,
  output wire          io_outputs_2_rsp_ready,
  input  wire          io_outputs_2_rsp_payload_last,
  input  wire [1:0]    io_outputs_2_rsp_payload_fragment_source,
  input  wire [0:0]    io_outputs_2_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_outputs_2_rsp_payload_fragment_data,
  input  wire [43:0]   io_outputs_2_rsp_payload_fragment_context,
  output reg           io_outputs_3_cmd_valid,
  input  wire          io_outputs_3_cmd_ready,
  output wire          io_outputs_3_cmd_payload_last,
  output wire [1:0]    io_outputs_3_cmd_payload_fragment_source,
  output wire [0:0]    io_outputs_3_cmd_payload_fragment_opcode,
  output wire [31:0]   io_outputs_3_cmd_payload_fragment_address,
  output wire [5:0]    io_outputs_3_cmd_payload_fragment_length,
  output wire [63:0]   io_outputs_3_cmd_payload_fragment_data,
  output wire [7:0]    io_outputs_3_cmd_payload_fragment_mask,
  output wire [43:0]   io_outputs_3_cmd_payload_fragment_context,
  input  wire          io_outputs_3_rsp_valid,
  output wire          io_outputs_3_rsp_ready,
  input  wire          io_outputs_3_rsp_payload_last,
  input  wire [1:0]    io_outputs_3_rsp_payload_fragment_source,
  input  wire [0:0]    io_outputs_3_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_outputs_3_rsp_payload_fragment_data,
  input  wire [43:0]   io_outputs_3_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg                 bmbErrorSlave_1_io_input_cmd_valid;
  wire                bmbErrorSlave_1_io_input_cmd_ready;
  wire                bmbErrorSlave_1_io_input_rsp_valid;
  wire                bmbErrorSlave_1_io_input_rsp_payload_last;
  wire       [1:0]    bmbErrorSlave_1_io_input_rsp_payload_fragment_source;
  wire       [0:0]    bmbErrorSlave_1_io_input_rsp_payload_fragment_opcode;
  wire       [63:0]   bmbErrorSlave_1_io_input_rsp_payload_fragment_data;
  wire       [43:0]   bmbErrorSlave_1_io_input_rsp_payload_fragment_context;
  wire                streamArbiter_10_io_inputs_0_ready;
  wire                streamArbiter_10_io_inputs_1_ready;
  wire                streamArbiter_10_io_inputs_2_ready;
  wire                streamArbiter_10_io_inputs_3_ready;
  wire                streamArbiter_10_io_inputs_4_ready;
  wire                streamArbiter_10_io_output_valid;
  wire                streamArbiter_10_io_output_payload_last;
  wire       [1:0]    streamArbiter_10_io_output_payload_fragment_source;
  wire       [0:0]    streamArbiter_10_io_output_payload_fragment_opcode;
  wire       [63:0]   streamArbiter_10_io_output_payload_fragment_data;
  wire       [43:0]   streamArbiter_10_io_output_payload_fragment_context;
  wire       [2:0]    streamArbiter_10_io_chosen;
  wire       [4:0]    streamArbiter_10_io_chosenOH;
  wire       [5:0]    _zz_logic_sources_0_rspPendingCounter;
  wire       [5:0]    _zz_logic_sources_0_rspPendingCounter_1;
  wire       [0:0]    _zz_logic_sources_0_rspPendingCounter_2;
  wire       [5:0]    _zz_logic_sources_0_rspPendingCounter_3;
  wire       [0:0]    _zz_logic_sources_0_rspPendingCounter_4;
  wire       [5:0]    _zz_logic_sources_1_rspPendingCounter;
  wire       [5:0]    _zz_logic_sources_1_rspPendingCounter_1;
  wire       [0:0]    _zz_logic_sources_1_rspPendingCounter_2;
  wire       [5:0]    _zz_logic_sources_1_rspPendingCounter_3;
  wire       [0:0]    _zz_logic_sources_1_rspPendingCounter_4;
  wire       [5:0]    _zz_logic_sources_2_rspPendingCounter;
  wire       [5:0]    _zz_logic_sources_2_rspPendingCounter_1;
  wire       [0:0]    _zz_logic_sources_2_rspPendingCounter_2;
  wire       [5:0]    _zz_logic_sources_2_rspPendingCounter_3;
  wire       [0:0]    _zz_logic_sources_2_rspPendingCounter_4;
  wire       [5:0]    _zz_logic_sources_3_rspPendingCounter;
  wire       [5:0]    _zz_logic_sources_3_rspPendingCounter_1;
  wire       [0:0]    _zz_logic_sources_3_rspPendingCounter_2;
  wire       [5:0]    _zz_logic_sources_3_rspPendingCounter_3;
  wire       [0:0]    _zz_logic_sources_3_rspPendingCounter_4;
  wire                logic_hits_0;
  wire                logic_hits_1;
  wire                logic_hits_2;
  wire                logic_hits_3;
  wire                logic_hits_4;
  wire                _zz_io_outputs_0_cmd_payload_last;
  wire                _zz_io_outputs_1_cmd_payload_last;
  wire                _zz_io_outputs_2_cmd_payload_last;
  wire                _zz_io_outputs_3_cmd_payload_last;
  wire                _zz_io_input_cmd_payload_last;
  wire                logic_sources_0_hit;
  wire                io_input_cmd_fire;
  wire                when_BmbDecoder_l187;
  reg                 logic_sources_0_rspHits_0;
  reg                 logic_sources_0_rspHits_1;
  reg                 logic_sources_0_rspHits_2;
  reg                 logic_sources_0_rspHits_3;
  reg                 logic_sources_0_rspHits_4;
  reg        [5:0]    logic_sources_0_rspPendingCounter;
  wire                io_input_rsp_fire;
  wire                logic_sources_0_rspPending;
  wire                logic_sources_0_full;
  wire                logic_sources_0_cmdWait;
  wire                logic_sources_1_hit;
  wire                when_BmbDecoder_l187_1;
  reg                 logic_sources_1_rspHits_0;
  reg                 logic_sources_1_rspHits_1;
  reg                 logic_sources_1_rspHits_2;
  reg                 logic_sources_1_rspHits_3;
  reg                 logic_sources_1_rspHits_4;
  reg        [5:0]    logic_sources_1_rspPendingCounter;
  wire                logic_sources_1_rspPending;
  wire                logic_sources_1_full;
  wire                logic_sources_1_cmdWait;
  wire                logic_sources_2_hit;
  wire                when_BmbDecoder_l187_2;
  reg                 logic_sources_2_rspHits_0;
  reg                 logic_sources_2_rspHits_1;
  reg                 logic_sources_2_rspHits_2;
  reg                 logic_sources_2_rspHits_3;
  reg                 logic_sources_2_rspHits_4;
  reg        [5:0]    logic_sources_2_rspPendingCounter;
  wire                logic_sources_2_rspPending;
  wire                logic_sources_2_full;
  wire                logic_sources_2_cmdWait;
  wire                logic_sources_3_hit;
  wire                when_BmbDecoder_l187_3;
  reg                 logic_sources_3_rspHits_0;
  reg                 logic_sources_3_rspHits_1;
  reg                 logic_sources_3_rspHits_2;
  reg                 logic_sources_3_rspHits_3;
  reg                 logic_sources_3_rspHits_4;
  reg        [5:0]    logic_sources_3_rspPendingCounter;
  wire                logic_sources_3_rspPending;
  wire                logic_sources_3_full;
  wire                logic_sources_3_cmdWait;
  wire                when_BmbDecoder_l196;
  wire                streamArbiter_10_io_output_combStage_valid;
  wire                streamArbiter_10_io_output_combStage_ready;
  wire                streamArbiter_10_io_output_combStage_payload_last;
  wire       [1:0]    streamArbiter_10_io_output_combStage_payload_fragment_source;
  wire       [0:0]    streamArbiter_10_io_output_combStage_payload_fragment_opcode;
  wire       [63:0]   streamArbiter_10_io_output_combStage_payload_fragment_data;
  wire       [43:0]   streamArbiter_10_io_output_combStage_payload_fragment_context;

  assign _zz_logic_sources_0_rspPendingCounter = (logic_sources_0_rspPendingCounter + _zz_logic_sources_0_rspPendingCounter_1);
  assign _zz_logic_sources_0_rspPendingCounter_2 = ((io_input_cmd_fire && io_input_cmd_payload_last) && (io_input_cmd_payload_fragment_source == 2'b00));
  assign _zz_logic_sources_0_rspPendingCounter_1 = {5'd0, _zz_logic_sources_0_rspPendingCounter_2};
  assign _zz_logic_sources_0_rspPendingCounter_4 = ((io_input_rsp_fire && io_input_rsp_payload_last) && (io_input_rsp_payload_fragment_source == 2'b00));
  assign _zz_logic_sources_0_rspPendingCounter_3 = {5'd0, _zz_logic_sources_0_rspPendingCounter_4};
  assign _zz_logic_sources_1_rspPendingCounter = (logic_sources_1_rspPendingCounter + _zz_logic_sources_1_rspPendingCounter_1);
  assign _zz_logic_sources_1_rspPendingCounter_2 = ((io_input_cmd_fire && io_input_cmd_payload_last) && (io_input_cmd_payload_fragment_source == 2'b10));
  assign _zz_logic_sources_1_rspPendingCounter_1 = {5'd0, _zz_logic_sources_1_rspPendingCounter_2};
  assign _zz_logic_sources_1_rspPendingCounter_4 = ((io_input_rsp_fire && io_input_rsp_payload_last) && (io_input_rsp_payload_fragment_source == 2'b10));
  assign _zz_logic_sources_1_rspPendingCounter_3 = {5'd0, _zz_logic_sources_1_rspPendingCounter_4};
  assign _zz_logic_sources_2_rspPendingCounter = (logic_sources_2_rspPendingCounter + _zz_logic_sources_2_rspPendingCounter_1);
  assign _zz_logic_sources_2_rspPendingCounter_2 = ((io_input_cmd_fire && io_input_cmd_payload_last) && (io_input_cmd_payload_fragment_source == 2'b01));
  assign _zz_logic_sources_2_rspPendingCounter_1 = {5'd0, _zz_logic_sources_2_rspPendingCounter_2};
  assign _zz_logic_sources_2_rspPendingCounter_4 = ((io_input_rsp_fire && io_input_rsp_payload_last) && (io_input_rsp_payload_fragment_source == 2'b01));
  assign _zz_logic_sources_2_rspPendingCounter_3 = {5'd0, _zz_logic_sources_2_rspPendingCounter_4};
  assign _zz_logic_sources_3_rspPendingCounter = (logic_sources_3_rspPendingCounter + _zz_logic_sources_3_rspPendingCounter_1);
  assign _zz_logic_sources_3_rspPendingCounter_2 = ((io_input_cmd_fire && io_input_cmd_payload_last) && (io_input_cmd_payload_fragment_source == 2'b11));
  assign _zz_logic_sources_3_rspPendingCounter_1 = {5'd0, _zz_logic_sources_3_rspPendingCounter_2};
  assign _zz_logic_sources_3_rspPendingCounter_4 = ((io_input_rsp_fire && io_input_rsp_payload_last) && (io_input_rsp_payload_fragment_source == 2'b11));
  assign _zz_logic_sources_3_rspPendingCounter_3 = {5'd0, _zz_logic_sources_3_rspPendingCounter_4};
  BmbErrorSlave bmbErrorSlave_1 (
    .io_input_cmd_valid                    (bmbErrorSlave_1_io_input_cmd_valid                         ), //i
    .io_input_cmd_ready                    (bmbErrorSlave_1_io_input_cmd_ready                         ), //o
    .io_input_cmd_payload_last             (_zz_io_input_cmd_payload_last                              ), //i
    .io_input_cmd_payload_fragment_source  (io_input_cmd_payload_fragment_source[1:0]                  ), //i
    .io_input_cmd_payload_fragment_opcode  (io_input_cmd_payload_fragment_opcode                       ), //i
    .io_input_cmd_payload_fragment_address (io_input_cmd_payload_fragment_address[31:0]                ), //i
    .io_input_cmd_payload_fragment_length  (io_input_cmd_payload_fragment_length[5:0]                  ), //i
    .io_input_cmd_payload_fragment_data    (io_input_cmd_payload_fragment_data[63:0]                   ), //i
    .io_input_cmd_payload_fragment_mask    (io_input_cmd_payload_fragment_mask[7:0]                    ), //i
    .io_input_cmd_payload_fragment_context (io_input_cmd_payload_fragment_context[43:0]                ), //i
    .io_input_rsp_valid                    (bmbErrorSlave_1_io_input_rsp_valid                         ), //o
    .io_input_rsp_ready                    (streamArbiter_10_io_inputs_4_ready                         ), //i
    .io_input_rsp_payload_last             (bmbErrorSlave_1_io_input_rsp_payload_last                  ), //o
    .io_input_rsp_payload_fragment_source  (bmbErrorSlave_1_io_input_rsp_payload_fragment_source[1:0]  ), //o
    .io_input_rsp_payload_fragment_opcode  (bmbErrorSlave_1_io_input_rsp_payload_fragment_opcode       ), //o
    .io_input_rsp_payload_fragment_data    (bmbErrorSlave_1_io_input_rsp_payload_fragment_data[63:0]   ), //o
    .io_input_rsp_payload_fragment_context (bmbErrorSlave_1_io_input_rsp_payload_fragment_context[43:0]), //o
    .io_systemClk                          (io_systemClk                                               ), //i
    .systemCd_logic_outputReset            (systemCd_logic_outputReset                                 )  //i
  );
  StreamArbiter_9 streamArbiter_10 (
    .io_inputs_0_valid                    (io_outputs_0_rsp_valid                                     ), //i
    .io_inputs_0_ready                    (streamArbiter_10_io_inputs_0_ready                         ), //o
    .io_inputs_0_payload_last             (io_outputs_0_rsp_payload_last                              ), //i
    .io_inputs_0_payload_fragment_source  (io_outputs_0_rsp_payload_fragment_source[1:0]              ), //i
    .io_inputs_0_payload_fragment_opcode  (io_outputs_0_rsp_payload_fragment_opcode                   ), //i
    .io_inputs_0_payload_fragment_data    (io_outputs_0_rsp_payload_fragment_data[63:0]               ), //i
    .io_inputs_0_payload_fragment_context (io_outputs_0_rsp_payload_fragment_context[43:0]            ), //i
    .io_inputs_1_valid                    (io_outputs_1_rsp_valid                                     ), //i
    .io_inputs_1_ready                    (streamArbiter_10_io_inputs_1_ready                         ), //o
    .io_inputs_1_payload_last             (io_outputs_1_rsp_payload_last                              ), //i
    .io_inputs_1_payload_fragment_source  (io_outputs_1_rsp_payload_fragment_source[1:0]              ), //i
    .io_inputs_1_payload_fragment_opcode  (io_outputs_1_rsp_payload_fragment_opcode                   ), //i
    .io_inputs_1_payload_fragment_data    (io_outputs_1_rsp_payload_fragment_data[63:0]               ), //i
    .io_inputs_1_payload_fragment_context (io_outputs_1_rsp_payload_fragment_context[43:0]            ), //i
    .io_inputs_2_valid                    (io_outputs_2_rsp_valid                                     ), //i
    .io_inputs_2_ready                    (streamArbiter_10_io_inputs_2_ready                         ), //o
    .io_inputs_2_payload_last             (io_outputs_2_rsp_payload_last                              ), //i
    .io_inputs_2_payload_fragment_source  (io_outputs_2_rsp_payload_fragment_source[1:0]              ), //i
    .io_inputs_2_payload_fragment_opcode  (io_outputs_2_rsp_payload_fragment_opcode                   ), //i
    .io_inputs_2_payload_fragment_data    (io_outputs_2_rsp_payload_fragment_data[63:0]               ), //i
    .io_inputs_2_payload_fragment_context (io_outputs_2_rsp_payload_fragment_context[43:0]            ), //i
    .io_inputs_3_valid                    (io_outputs_3_rsp_valid                                     ), //i
    .io_inputs_3_ready                    (streamArbiter_10_io_inputs_3_ready                         ), //o
    .io_inputs_3_payload_last             (io_outputs_3_rsp_payload_last                              ), //i
    .io_inputs_3_payload_fragment_source  (io_outputs_3_rsp_payload_fragment_source[1:0]              ), //i
    .io_inputs_3_payload_fragment_opcode  (io_outputs_3_rsp_payload_fragment_opcode                   ), //i
    .io_inputs_3_payload_fragment_data    (io_outputs_3_rsp_payload_fragment_data[63:0]               ), //i
    .io_inputs_3_payload_fragment_context (io_outputs_3_rsp_payload_fragment_context[43:0]            ), //i
    .io_inputs_4_valid                    (bmbErrorSlave_1_io_input_rsp_valid                         ), //i
    .io_inputs_4_ready                    (streamArbiter_10_io_inputs_4_ready                         ), //o
    .io_inputs_4_payload_last             (bmbErrorSlave_1_io_input_rsp_payload_last                  ), //i
    .io_inputs_4_payload_fragment_source  (bmbErrorSlave_1_io_input_rsp_payload_fragment_source[1:0]  ), //i
    .io_inputs_4_payload_fragment_opcode  (bmbErrorSlave_1_io_input_rsp_payload_fragment_opcode       ), //i
    .io_inputs_4_payload_fragment_data    (bmbErrorSlave_1_io_input_rsp_payload_fragment_data[63:0]   ), //i
    .io_inputs_4_payload_fragment_context (bmbErrorSlave_1_io_input_rsp_payload_fragment_context[43:0]), //i
    .io_output_valid                      (streamArbiter_10_io_output_valid                           ), //o
    .io_output_ready                      (streamArbiter_10_io_output_combStage_ready                 ), //i
    .io_output_payload_last               (streamArbiter_10_io_output_payload_last                    ), //o
    .io_output_payload_fragment_source    (streamArbiter_10_io_output_payload_fragment_source[1:0]    ), //o
    .io_output_payload_fragment_opcode    (streamArbiter_10_io_output_payload_fragment_opcode         ), //o
    .io_output_payload_fragment_data      (streamArbiter_10_io_output_payload_fragment_data[63:0]     ), //o
    .io_output_payload_fragment_context   (streamArbiter_10_io_output_payload_fragment_context[43:0]  ), //o
    .io_chosen                            (streamArbiter_10_io_chosen[2:0]                            ), //o
    .io_chosenOH                          (streamArbiter_10_io_chosenOH[4:0]                          ), //o
    .io_systemClk                         (io_systemClk                                               ), //i
    .systemCd_logic_outputReset           (systemCd_logic_outputReset                                 )  //i
  );
  assign logic_hits_0 = ((io_input_cmd_payload_fragment_address & (~ 32'h000007ff)) == 32'hf9000000);
  always @(*) begin
    io_outputs_0_cmd_valid = (io_input_cmd_valid && logic_hits_0);
    if(when_BmbDecoder_l196) begin
      io_outputs_0_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_0_cmd_payload_last = io_input_cmd_payload_last;
  assign io_outputs_0_cmd_payload_last = _zz_io_outputs_0_cmd_payload_last;
  assign io_outputs_0_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_outputs_0_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_outputs_0_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_outputs_0_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_outputs_0_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_outputs_0_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_outputs_0_cmd_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign logic_hits_1 = ((io_input_cmd_payload_fragment_address & (~ 32'h00ffffff)) == 32'hf8000000);
  always @(*) begin
    io_outputs_1_cmd_valid = (io_input_cmd_valid && logic_hits_1);
    if(when_BmbDecoder_l196) begin
      io_outputs_1_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_1_cmd_payload_last = io_input_cmd_payload_last;
  assign io_outputs_1_cmd_payload_last = _zz_io_outputs_1_cmd_payload_last;
  assign io_outputs_1_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_outputs_1_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_outputs_1_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_outputs_1_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_outputs_1_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_outputs_1_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_outputs_1_cmd_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign logic_hits_2 = ((32'h00001000 <= io_input_cmd_payload_fragment_address) && (io_input_cmd_payload_fragment_address < 32'he0001000));
  always @(*) begin
    io_outputs_2_cmd_valid = (io_input_cmd_valid && logic_hits_2);
    if(when_BmbDecoder_l196) begin
      io_outputs_2_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_2_cmd_payload_last = io_input_cmd_payload_last;
  assign io_outputs_2_cmd_payload_last = _zz_io_outputs_2_cmd_payload_last;
  assign io_outputs_2_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_outputs_2_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_outputs_2_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_outputs_2_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_outputs_2_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_outputs_2_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_outputs_2_cmd_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign logic_hits_3 = ((io_input_cmd_payload_fragment_address & (~ 32'h00ffffff)) == 32'he1000000);
  always @(*) begin
    io_outputs_3_cmd_valid = (io_input_cmd_valid && logic_hits_3);
    if(when_BmbDecoder_l196) begin
      io_outputs_3_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_outputs_3_cmd_payload_last = io_input_cmd_payload_last;
  assign io_outputs_3_cmd_payload_last = _zz_io_outputs_3_cmd_payload_last;
  assign io_outputs_3_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_outputs_3_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_outputs_3_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_outputs_3_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_outputs_3_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_outputs_3_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_outputs_3_cmd_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign logic_hits_4 = (! (|{logic_hits_3,{logic_hits_2,{logic_hits_1,logic_hits_0}}}));
  always @(*) begin
    bmbErrorSlave_1_io_input_cmd_valid = (io_input_cmd_valid && logic_hits_4);
    if(when_BmbDecoder_l196) begin
      bmbErrorSlave_1_io_input_cmd_valid = 1'b0;
    end
  end

  assign _zz_io_input_cmd_payload_last = io_input_cmd_payload_last;
  always @(*) begin
    io_input_cmd_ready = (|{(logic_hits_4 && bmbErrorSlave_1_io_input_cmd_ready),{(logic_hits_3 && io_outputs_3_cmd_ready),{(logic_hits_2 && io_outputs_2_cmd_ready),{(logic_hits_1 && io_outputs_1_cmd_ready),(logic_hits_0 && io_outputs_0_cmd_ready)}}}});
    if(when_BmbDecoder_l196) begin
      io_input_cmd_ready = 1'b0;
    end
  end

  assign logic_sources_0_hit = (io_input_cmd_payload_fragment_source == 2'b00);
  assign io_input_cmd_fire = (io_input_cmd_valid && io_input_cmd_ready);
  assign when_BmbDecoder_l187 = (io_input_cmd_fire && logic_sources_0_hit);
  assign io_input_rsp_fire = (io_input_rsp_valid && io_input_rsp_ready);
  assign logic_sources_0_rspPending = (logic_sources_0_rspPendingCounter != 6'h0);
  assign logic_sources_0_full = (logic_sources_0_rspPendingCounter == 6'h3f);
  assign logic_sources_0_cmdWait = (logic_sources_0_hit && ((logic_sources_0_rspPending && (((((logic_hits_0 != logic_sources_0_rspHits_0) || (logic_hits_1 != logic_sources_0_rspHits_1)) || (logic_hits_2 != logic_sources_0_rspHits_2)) || (logic_hits_3 != logic_sources_0_rspHits_3)) || (logic_hits_4 != logic_sources_0_rspHits_4))) || logic_sources_0_full));
  assign logic_sources_1_hit = (io_input_cmd_payload_fragment_source == 2'b10);
  assign when_BmbDecoder_l187_1 = (io_input_cmd_fire && logic_sources_1_hit);
  assign logic_sources_1_rspPending = (logic_sources_1_rspPendingCounter != 6'h0);
  assign logic_sources_1_full = (logic_sources_1_rspPendingCounter == 6'h3f);
  assign logic_sources_1_cmdWait = (logic_sources_1_hit && ((logic_sources_1_rspPending && (((((logic_hits_0 != logic_sources_1_rspHits_0) || (logic_hits_1 != logic_sources_1_rspHits_1)) || (logic_hits_2 != logic_sources_1_rspHits_2)) || (logic_hits_3 != logic_sources_1_rspHits_3)) || (logic_hits_4 != logic_sources_1_rspHits_4))) || logic_sources_1_full));
  assign logic_sources_2_hit = (io_input_cmd_payload_fragment_source == 2'b01);
  assign when_BmbDecoder_l187_2 = (io_input_cmd_fire && logic_sources_2_hit);
  assign logic_sources_2_rspPending = (logic_sources_2_rspPendingCounter != 6'h0);
  assign logic_sources_2_full = (logic_sources_2_rspPendingCounter == 6'h3f);
  assign logic_sources_2_cmdWait = (logic_sources_2_hit && ((logic_sources_2_rspPending && (((((logic_hits_0 != logic_sources_2_rspHits_0) || (logic_hits_1 != logic_sources_2_rspHits_1)) || (logic_hits_2 != logic_sources_2_rspHits_2)) || (logic_hits_3 != logic_sources_2_rspHits_3)) || (logic_hits_4 != logic_sources_2_rspHits_4))) || logic_sources_2_full));
  assign logic_sources_3_hit = (io_input_cmd_payload_fragment_source == 2'b11);
  assign when_BmbDecoder_l187_3 = (io_input_cmd_fire && logic_sources_3_hit);
  assign logic_sources_3_rspPending = (logic_sources_3_rspPendingCounter != 6'h0);
  assign logic_sources_3_full = (logic_sources_3_rspPendingCounter == 6'h3f);
  assign logic_sources_3_cmdWait = (logic_sources_3_hit && ((logic_sources_3_rspPending && (((((logic_hits_0 != logic_sources_3_rspHits_0) || (logic_hits_1 != logic_sources_3_rspHits_1)) || (logic_hits_2 != logic_sources_3_rspHits_2)) || (logic_hits_3 != logic_sources_3_rspHits_3)) || (logic_hits_4 != logic_sources_3_rspHits_4))) || logic_sources_3_full));
  assign when_BmbDecoder_l196 = (|{logic_sources_3_cmdWait,{logic_sources_2_cmdWait,{logic_sources_1_cmdWait,logic_sources_0_cmdWait}}});
  assign io_outputs_0_rsp_ready = streamArbiter_10_io_inputs_0_ready;
  assign io_outputs_1_rsp_ready = streamArbiter_10_io_inputs_1_ready;
  assign io_outputs_2_rsp_ready = streamArbiter_10_io_inputs_2_ready;
  assign io_outputs_3_rsp_ready = streamArbiter_10_io_inputs_3_ready;
  assign streamArbiter_10_io_output_combStage_valid = streamArbiter_10_io_output_valid;
  assign streamArbiter_10_io_output_combStage_payload_last = streamArbiter_10_io_output_payload_last;
  assign streamArbiter_10_io_output_combStage_payload_fragment_source = streamArbiter_10_io_output_payload_fragment_source;
  assign streamArbiter_10_io_output_combStage_payload_fragment_opcode = streamArbiter_10_io_output_payload_fragment_opcode;
  assign streamArbiter_10_io_output_combStage_payload_fragment_data = streamArbiter_10_io_output_payload_fragment_data;
  assign streamArbiter_10_io_output_combStage_payload_fragment_context = streamArbiter_10_io_output_payload_fragment_context;
  assign io_input_rsp_valid = streamArbiter_10_io_output_combStage_valid;
  assign streamArbiter_10_io_output_combStage_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = streamArbiter_10_io_output_combStage_payload_last;
  assign io_input_rsp_payload_fragment_source = streamArbiter_10_io_output_combStage_payload_fragment_source;
  assign io_input_rsp_payload_fragment_opcode = streamArbiter_10_io_output_combStage_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = streamArbiter_10_io_output_combStage_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = streamArbiter_10_io_output_combStage_payload_fragment_context;
  always @(posedge io_systemClk) begin
    if(when_BmbDecoder_l187) begin
      logic_sources_0_rspHits_0 <= logic_hits_0;
      logic_sources_0_rspHits_1 <= logic_hits_1;
      logic_sources_0_rspHits_2 <= logic_hits_2;
      logic_sources_0_rspHits_3 <= logic_hits_3;
      logic_sources_0_rspHits_4 <= logic_hits_4;
    end
    if(when_BmbDecoder_l187_1) begin
      logic_sources_1_rspHits_0 <= logic_hits_0;
      logic_sources_1_rspHits_1 <= logic_hits_1;
      logic_sources_1_rspHits_2 <= logic_hits_2;
      logic_sources_1_rspHits_3 <= logic_hits_3;
      logic_sources_1_rspHits_4 <= logic_hits_4;
    end
    if(when_BmbDecoder_l187_2) begin
      logic_sources_2_rspHits_0 <= logic_hits_0;
      logic_sources_2_rspHits_1 <= logic_hits_1;
      logic_sources_2_rspHits_2 <= logic_hits_2;
      logic_sources_2_rspHits_3 <= logic_hits_3;
      logic_sources_2_rspHits_4 <= logic_hits_4;
    end
    if(when_BmbDecoder_l187_3) begin
      logic_sources_3_rspHits_0 <= logic_hits_0;
      logic_sources_3_rspHits_1 <= logic_hits_1;
      logic_sources_3_rspHits_2 <= logic_hits_2;
      logic_sources_3_rspHits_3 <= logic_hits_3;
      logic_sources_3_rspHits_4 <= logic_hits_4;
    end
  end

  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      logic_sources_0_rspPendingCounter <= 6'h0;
      logic_sources_1_rspPendingCounter <= 6'h0;
      logic_sources_2_rspPendingCounter <= 6'h0;
      logic_sources_3_rspPendingCounter <= 6'h0;
    end else begin
      logic_sources_0_rspPendingCounter <= (_zz_logic_sources_0_rspPendingCounter - _zz_logic_sources_0_rspPendingCounter_3);
      logic_sources_1_rspPendingCounter <= (_zz_logic_sources_1_rspPendingCounter - _zz_logic_sources_1_rspPendingCounter_3);
      logic_sources_2_rspPendingCounter <= (_zz_logic_sources_2_rspPendingCounter - _zz_logic_sources_2_rspPendingCounter_3);
      logic_sources_3_rspPendingCounter <= (_zz_logic_sources_3_rspPendingCounter - _zz_logic_sources_3_rspPendingCounter_3);
    end
  end


endmodule

module BmbToAxi4SharedBridge_1 (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [31:0]   io_input_cmd_payload_fragment_data,
  input  wire [3:0]    io_input_cmd_payload_fragment_mask,
  input  wire [44:0]   io_input_cmd_payload_fragment_context,
  output reg           io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output reg           io_input_rsp_payload_last,
  output reg  [1:0]    io_input_rsp_payload_fragment_source,
  output reg  [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [31:0]   io_input_rsp_payload_fragment_data,
  output reg  [44:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_arw_valid,
  input  wire          io_output_arw_ready,
  output wire [31:0]   io_output_arw_payload_addr,
  output wire [7:0]    io_output_arw_payload_len,
  output wire [2:0]    io_output_arw_payload_size,
  output wire [3:0]    io_output_arw_payload_cache,
  output wire [2:0]    io_output_arw_payload_prot,
  output wire          io_output_arw_payload_write,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [31:0]   io_output_w_payload_data,
  output wire [3:0]    io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [31:0]   io_output_r_payload_data,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire                writeCmdInfo_fifo_io_pop_ready;
  wire                readCmdInfo_fifo_io_pop_ready;
  wire                writeCmdInfo_fifo_io_push_ready;
  wire                writeCmdInfo_fifo_io_pop_valid;
  wire       [1:0]    writeCmdInfo_fifo_io_pop_payload_source;
  wire       [44:0]   writeCmdInfo_fifo_io_pop_payload_context;
  wire       [3:0]    writeCmdInfo_fifo_io_occupancy;
  wire       [3:0]    writeCmdInfo_fifo_io_availability;
  wire                readCmdInfo_fifo_io_push_ready;
  wire                readCmdInfo_fifo_io_pop_valid;
  wire       [1:0]    readCmdInfo_fifo_io_pop_payload_source;
  wire       [44:0]   readCmdInfo_fifo_io_pop_payload_context;
  wire       [3:0]    readCmdInfo_fifo_io_occupancy;
  wire       [3:0]    readCmdInfo_fifo_io_availability;
  wire       [3:0]    _zz_io_output_arw_payload_len;
  reg                 pendingWrite;
  reg        [2:0]    pendingCounter;
  wire                io_input_cmd_fire;
  wire                when_Utils_l706;
  wire                io_input_rsp_fire;
  wire                when_Utils_l709;
  reg                 states_0_counter_incrementIt;
  reg                 states_0_counter_decrementIt;
  wire       [2:0]    states_0_counter_valueNext;
  reg        [2:0]    states_0_counter_value;
  wire                states_0_counter_mayOverflow;
  wire                states_0_counter_willOverflowIfInc;
  wire                states_0_counter_willOverflow;
  reg        [2:0]    states_0_counter_finalIncrement;
  wire                when_Utils_l735;
  wire                when_Utils_l737;
  wire                when_BmbToAxi4Bridge_l45;
  reg                 states_0_write;
  wire                when_BmbToAxi4Bridge_l47;
  wire                when_Utils_l706_1;
  wire                when_Utils_l709_1;
  reg                 states_1_counter_incrementIt;
  reg                 states_1_counter_decrementIt;
  wire       [2:0]    states_1_counter_valueNext;
  reg        [2:0]    states_1_counter_value;
  wire                states_1_counter_mayOverflow;
  wire                states_1_counter_willOverflowIfInc;
  wire                states_1_counter_willOverflow;
  reg        [2:0]    states_1_counter_finalIncrement;
  wire                when_Utils_l735_1;
  wire                when_Utils_l737_1;
  wire                when_BmbToAxi4Bridge_l45_1;
  reg                 states_1_write;
  wire                when_BmbToAxi4Bridge_l47_1;
  wire                when_Utils_l706_2;
  wire                when_Utils_l709_2;
  reg                 states_2_counter_incrementIt;
  reg                 states_2_counter_decrementIt;
  wire       [2:0]    states_2_counter_valueNext;
  reg        [2:0]    states_2_counter_value;
  wire                states_2_counter_mayOverflow;
  wire                states_2_counter_willOverflowIfInc;
  wire                states_2_counter_willOverflow;
  reg        [2:0]    states_2_counter_finalIncrement;
  wire                when_Utils_l735_2;
  wire                when_Utils_l737_2;
  wire                when_BmbToAxi4Bridge_l45_2;
  reg                 states_2_write;
  wire                when_BmbToAxi4Bridge_l47_2;
  wire                when_Utils_l706_3;
  wire                when_Utils_l709_3;
  reg                 states_3_counter_incrementIt;
  reg                 states_3_counter_decrementIt;
  wire       [2:0]    states_3_counter_valueNext;
  reg        [2:0]    states_3_counter_value;
  wire                states_3_counter_mayOverflow;
  wire                states_3_counter_willOverflowIfInc;
  wire                states_3_counter_willOverflow;
  reg        [2:0]    states_3_counter_finalIncrement;
  wire                when_Utils_l735_3;
  wire                when_Utils_l737_3;
  wire                when_BmbToAxi4Bridge_l45_3;
  reg                 states_3_write;
  wire                when_BmbToAxi4Bridge_l47_3;
  wire                hazard;
  wire                _zz_io_input_cmd_ready;
  wire                _zz_cmdFork_valid;
  reg                 _zz_io_input_cmd_ready_1;
  wire                _zz_cmdFork_payload_last;
  wire       [1:0]    _zz_cmdFork_payload_fragment_source;
  wire       [0:0]    _zz_cmdFork_payload_fragment_opcode;
  wire       [31:0]   _zz_cmdFork_payload_fragment_address;
  wire       [5:0]    _zz_cmdFork_payload_fragment_length;
  wire       [31:0]   _zz_cmdFork_payload_fragment_data;
  wire       [3:0]    _zz_cmdFork_payload_fragment_mask;
  wire       [44:0]   _zz_cmdFork_payload_fragment_context;
  wire                cmdFork_valid;
  reg                 cmdFork_ready;
  wire                cmdFork_payload_last;
  wire       [1:0]    cmdFork_payload_fragment_source;
  wire       [0:0]    cmdFork_payload_fragment_opcode;
  wire       [31:0]   cmdFork_payload_fragment_address;
  wire       [5:0]    cmdFork_payload_fragment_length;
  wire       [31:0]   cmdFork_payload_fragment_data;
  wire       [3:0]    cmdFork_payload_fragment_mask;
  wire       [44:0]   cmdFork_payload_fragment_context;
  wire                dataFork_valid;
  reg                 dataFork_ready;
  wire                dataFork_payload_last;
  wire       [1:0]    dataFork_payload_fragment_source;
  wire       [0:0]    dataFork_payload_fragment_opcode;
  wire       [31:0]   dataFork_payload_fragment_address;
  wire       [5:0]    dataFork_payload_fragment_length;
  wire       [31:0]   dataFork_payload_fragment_data;
  wire       [3:0]    dataFork_payload_fragment_mask;
  wire       [44:0]   dataFork_payload_fragment_context;
  reg                 _zz_cmdFork_valid_1;
  reg                 _zz_dataFork_valid;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdFork_fire;
  wire                dataFork_fire;
  reg                 io_input_cmd_payload_first;
  wire                when_Stream_l445;
  reg                 cmdStage_valid;
  wire                cmdStage_ready;
  wire                cmdStage_payload_last;
  wire       [1:0]    cmdStage_payload_fragment_source;
  wire       [0:0]    cmdStage_payload_fragment_opcode;
  wire       [31:0]   cmdStage_payload_fragment_address;
  wire       [5:0]    cmdStage_payload_fragment_length;
  wire       [31:0]   cmdStage_payload_fragment_data;
  wire       [3:0]    cmdStage_payload_fragment_mask;
  wire       [44:0]   cmdStage_payload_fragment_context;
  wire                when_Stream_l445_1;
  reg                 dataStage_valid;
  wire                dataStage_ready;
  wire                dataStage_payload_last;
  wire       [1:0]    dataStage_payload_fragment_source;
  wire       [0:0]    dataStage_payload_fragment_opcode;
  wire       [31:0]   dataStage_payload_fragment_address;
  wire       [5:0]    dataStage_payload_fragment_length;
  wire       [31:0]   dataStage_payload_fragment_data;
  wire       [3:0]    dataStage_payload_fragment_mask;
  wire       [44:0]   dataStage_payload_fragment_context;
  wire                writeCmdInfo_valid;
  wire                writeCmdInfo_ready;
  wire       [1:0]    writeCmdInfo_payload_source;
  wire       [44:0]   writeCmdInfo_payload_context;
  wire                readCmdInfo_valid;
  wire                readCmdInfo_ready;
  wire       [1:0]    readCmdInfo_payload_source;
  wire       [44:0]   readCmdInfo_payload_context;
  wire                cmdStage_fire;
  wire                writeRspInfo_valid;
  wire                writeRspInfo_ready;
  wire       [1:0]    writeRspInfo_payload_source;
  wire       [44:0]   writeRspInfo_payload_context;
  reg                 writeCmdInfo_fifo_io_pop_rValid;
  wire                writeRspInfo_fire;
  reg        [1:0]    writeCmdInfo_fifo_io_pop_rData_source;
  reg        [44:0]   writeCmdInfo_fifo_io_pop_rData_context;
  wire                readRspInfo_valid;
  wire                readRspInfo_ready;
  wire       [1:0]    readRspInfo_payload_source;
  wire       [44:0]   readRspInfo_payload_context;
  reg                 readCmdInfo_fifo_io_pop_rValid;
  wire                readRspInfo_fire;
  reg        [1:0]    readCmdInfo_fifo_io_pop_rData_source;
  reg        [44:0]   readCmdInfo_fifo_io_pop_rData_context;
  wire                _zz_io_output_arw_valid;
  reg                 rspSelLock;
  wire                when_BmbToAxi4Bridge_l87;
  wire                io_output_r_fire;
  wire                io_output_b_fire;
  wire                when_BmbToAxi4Bridge_l87_1;
  wire                when_BmbToAxi4Bridge_l88;
  reg                 rspSelReadLast;
  wire                rspSelRead;
  wire                when_BmbToAxi4Bridge_l108;

  assign _zz_io_output_arw_payload_len = io_input_cmd_payload_fragment_length[5 : 2];
  StreamFifo_7 writeCmdInfo_fifo (
    .io_push_valid                  (writeCmdInfo_valid                            ), //i
    .io_push_ready                  (writeCmdInfo_fifo_io_push_ready               ), //o
    .io_push_payload_source         (writeCmdInfo_payload_source[1:0]              ), //i
    .io_push_payload_context        (writeCmdInfo_payload_context[44:0]            ), //i
    .io_pop_valid                   (writeCmdInfo_fifo_io_pop_valid                ), //o
    .io_pop_ready                   (writeCmdInfo_fifo_io_pop_ready                ), //i
    .io_pop_payload_source          (writeCmdInfo_fifo_io_pop_payload_source[1:0]  ), //o
    .io_pop_payload_context         (writeCmdInfo_fifo_io_pop_payload_context[44:0]), //o
    .io_flush                       (1'b0                                          ), //i
    .io_occupancy                   (writeCmdInfo_fifo_io_occupancy[3:0]           ), //o
    .io_availability                (writeCmdInfo_fifo_io_availability[3:0]        ), //o
    .io_peripheralClk               (io_peripheralClk                              ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                )  //i
  );
  StreamFifo_7 readCmdInfo_fifo (
    .io_push_valid                  (readCmdInfo_valid                            ), //i
    .io_push_ready                  (readCmdInfo_fifo_io_push_ready               ), //o
    .io_push_payload_source         (readCmdInfo_payload_source[1:0]              ), //i
    .io_push_payload_context        (readCmdInfo_payload_context[44:0]            ), //i
    .io_pop_valid                   (readCmdInfo_fifo_io_pop_valid                ), //o
    .io_pop_ready                   (readCmdInfo_fifo_io_pop_ready                ), //i
    .io_pop_payload_source          (readCmdInfo_fifo_io_pop_payload_source[1:0]  ), //o
    .io_pop_payload_context         (readCmdInfo_fifo_io_pop_payload_context[44:0]), //o
    .io_flush                       (1'b0                                         ), //i
    .io_occupancy                   (readCmdInfo_fifo_io_occupancy[3:0]           ), //o
    .io_availability                (readCmdInfo_fifo_io_availability[3:0]        ), //o
    .io_peripheralClk               (io_peripheralClk                             ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset               )  //i
  );
  always @(*) begin
    pendingWrite = 1'bx;
    if(when_BmbToAxi4Bridge_l47) begin
      pendingWrite = states_0_write;
    end
    if(when_BmbToAxi4Bridge_l47_1) begin
      pendingWrite = states_1_write;
    end
    if(when_BmbToAxi4Bridge_l47_2) begin
      pendingWrite = states_2_write;
    end
    if(when_BmbToAxi4Bridge_l47_3) begin
      pendingWrite = states_3_write;
    end
  end

  always @(*) begin
    pendingCounter = 3'bxxx;
    if(when_BmbToAxi4Bridge_l47) begin
      pendingCounter = states_0_counter_value;
    end
    if(when_BmbToAxi4Bridge_l47_1) begin
      pendingCounter = states_1_counter_value;
    end
    if(when_BmbToAxi4Bridge_l47_2) begin
      pendingCounter = states_2_counter_value;
    end
    if(when_BmbToAxi4Bridge_l47_3) begin
      pendingCounter = states_3_counter_value;
    end
  end

  assign io_input_cmd_fire = (io_input_cmd_valid && io_input_cmd_ready);
  assign when_Utils_l706 = (((io_input_cmd_payload_fragment_source == 2'b00) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign io_input_rsp_fire = (io_input_rsp_valid && io_input_rsp_ready);
  assign when_Utils_l709 = (((io_input_rsp_payload_fragment_source == 2'b00) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_0_counter_incrementIt = 1'b0;
    if(when_Utils_l706) begin
      states_0_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_0_counter_decrementIt = 1'b0;
    if(when_Utils_l709) begin
      states_0_counter_decrementIt = 1'b1;
    end
  end

  assign states_0_counter_mayOverflow = (states_0_counter_value == 3'b111);
  assign states_0_counter_willOverflowIfInc = (states_0_counter_mayOverflow && (! states_0_counter_decrementIt));
  assign states_0_counter_willOverflow = (states_0_counter_willOverflowIfInc && states_0_counter_incrementIt);
  assign when_Utils_l735 = (states_0_counter_incrementIt && (! states_0_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735) begin
      states_0_counter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l737) begin
        states_0_counter_finalIncrement = 3'b111;
      end else begin
        states_0_counter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l737 = ((! states_0_counter_incrementIt) && states_0_counter_decrementIt);
  assign states_0_counter_valueNext = (states_0_counter_value + states_0_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45 = ((io_input_cmd_payload_fragment_source == 2'b00) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47 = (io_input_cmd_payload_fragment_source == 2'b00);
  assign when_Utils_l706_1 = (((io_input_cmd_payload_fragment_source == 2'b10) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign when_Utils_l709_1 = (((io_input_rsp_payload_fragment_source == 2'b10) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_1_counter_incrementIt = 1'b0;
    if(when_Utils_l706_1) begin
      states_1_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_1_counter_decrementIt = 1'b0;
    if(when_Utils_l709_1) begin
      states_1_counter_decrementIt = 1'b1;
    end
  end

  assign states_1_counter_mayOverflow = (states_1_counter_value == 3'b111);
  assign states_1_counter_willOverflowIfInc = (states_1_counter_mayOverflow && (! states_1_counter_decrementIt));
  assign states_1_counter_willOverflow = (states_1_counter_willOverflowIfInc && states_1_counter_incrementIt);
  assign when_Utils_l735_1 = (states_1_counter_incrementIt && (! states_1_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_1) begin
      states_1_counter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l737_1) begin
        states_1_counter_finalIncrement = 3'b111;
      end else begin
        states_1_counter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l737_1 = ((! states_1_counter_incrementIt) && states_1_counter_decrementIt);
  assign states_1_counter_valueNext = (states_1_counter_value + states_1_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45_1 = ((io_input_cmd_payload_fragment_source == 2'b10) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47_1 = (io_input_cmd_payload_fragment_source == 2'b10);
  assign when_Utils_l706_2 = (((io_input_cmd_payload_fragment_source == 2'b01) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign when_Utils_l709_2 = (((io_input_rsp_payload_fragment_source == 2'b01) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_2_counter_incrementIt = 1'b0;
    if(when_Utils_l706_2) begin
      states_2_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_2_counter_decrementIt = 1'b0;
    if(when_Utils_l709_2) begin
      states_2_counter_decrementIt = 1'b1;
    end
  end

  assign states_2_counter_mayOverflow = (states_2_counter_value == 3'b111);
  assign states_2_counter_willOverflowIfInc = (states_2_counter_mayOverflow && (! states_2_counter_decrementIt));
  assign states_2_counter_willOverflow = (states_2_counter_willOverflowIfInc && states_2_counter_incrementIt);
  assign when_Utils_l735_2 = (states_2_counter_incrementIt && (! states_2_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_2) begin
      states_2_counter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l737_2) begin
        states_2_counter_finalIncrement = 3'b111;
      end else begin
        states_2_counter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l737_2 = ((! states_2_counter_incrementIt) && states_2_counter_decrementIt);
  assign states_2_counter_valueNext = (states_2_counter_value + states_2_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45_2 = ((io_input_cmd_payload_fragment_source == 2'b01) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47_2 = (io_input_cmd_payload_fragment_source == 2'b01);
  assign when_Utils_l706_3 = (((io_input_cmd_payload_fragment_source == 2'b11) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign when_Utils_l709_3 = (((io_input_rsp_payload_fragment_source == 2'b11) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_3_counter_incrementIt = 1'b0;
    if(when_Utils_l706_3) begin
      states_3_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_3_counter_decrementIt = 1'b0;
    if(when_Utils_l709_3) begin
      states_3_counter_decrementIt = 1'b1;
    end
  end

  assign states_3_counter_mayOverflow = (states_3_counter_value == 3'b111);
  assign states_3_counter_willOverflowIfInc = (states_3_counter_mayOverflow && (! states_3_counter_decrementIt));
  assign states_3_counter_willOverflow = (states_3_counter_willOverflowIfInc && states_3_counter_incrementIt);
  assign when_Utils_l735_3 = (states_3_counter_incrementIt && (! states_3_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_3) begin
      states_3_counter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l737_3) begin
        states_3_counter_finalIncrement = 3'b111;
      end else begin
        states_3_counter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l737_3 = ((! states_3_counter_incrementIt) && states_3_counter_decrementIt);
  assign states_3_counter_valueNext = (states_3_counter_value + states_3_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45_3 = ((io_input_cmd_payload_fragment_source == 2'b11) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47_3 = (io_input_cmd_payload_fragment_source == 2'b11);
  assign hazard = ((((io_input_cmd_payload_fragment_opcode == 1'b1) != pendingWrite) && (pendingCounter != 3'b000)) || (pendingCounter == 3'b111));
  assign _zz_io_input_cmd_ready = (! hazard);
  assign _zz_cmdFork_valid = (io_input_cmd_valid && _zz_io_input_cmd_ready);
  assign io_input_cmd_ready = (_zz_io_input_cmd_ready_1 && _zz_io_input_cmd_ready);
  assign _zz_cmdFork_payload_last = io_input_cmd_payload_last;
  assign _zz_cmdFork_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign _zz_cmdFork_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign _zz_cmdFork_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign _zz_cmdFork_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign _zz_cmdFork_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign _zz_cmdFork_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign _zz_cmdFork_payload_fragment_context = io_input_cmd_payload_fragment_context;
  always @(*) begin
    _zz_io_input_cmd_ready_1 = 1'b1;
    if(when_Stream_l1063) begin
      _zz_io_input_cmd_ready_1 = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      _zz_io_input_cmd_ready_1 = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdFork_ready) && _zz_cmdFork_valid_1);
  assign when_Stream_l1063_1 = ((! dataFork_ready) && _zz_dataFork_valid);
  assign cmdFork_valid = (_zz_cmdFork_valid && _zz_cmdFork_valid_1);
  assign cmdFork_payload_last = _zz_cmdFork_payload_last;
  assign cmdFork_payload_fragment_source = _zz_cmdFork_payload_fragment_source;
  assign cmdFork_payload_fragment_opcode = _zz_cmdFork_payload_fragment_opcode;
  assign cmdFork_payload_fragment_address = _zz_cmdFork_payload_fragment_address;
  assign cmdFork_payload_fragment_length = _zz_cmdFork_payload_fragment_length;
  assign cmdFork_payload_fragment_data = _zz_cmdFork_payload_fragment_data;
  assign cmdFork_payload_fragment_mask = _zz_cmdFork_payload_fragment_mask;
  assign cmdFork_payload_fragment_context = _zz_cmdFork_payload_fragment_context;
  assign cmdFork_fire = (cmdFork_valid && cmdFork_ready);
  assign dataFork_valid = (_zz_cmdFork_valid && _zz_dataFork_valid);
  assign dataFork_payload_last = _zz_cmdFork_payload_last;
  assign dataFork_payload_fragment_source = _zz_cmdFork_payload_fragment_source;
  assign dataFork_payload_fragment_opcode = _zz_cmdFork_payload_fragment_opcode;
  assign dataFork_payload_fragment_address = _zz_cmdFork_payload_fragment_address;
  assign dataFork_payload_fragment_length = _zz_cmdFork_payload_fragment_length;
  assign dataFork_payload_fragment_data = _zz_cmdFork_payload_fragment_data;
  assign dataFork_payload_fragment_mask = _zz_cmdFork_payload_fragment_mask;
  assign dataFork_payload_fragment_context = _zz_cmdFork_payload_fragment_context;
  assign dataFork_fire = (dataFork_valid && dataFork_ready);
  assign when_Stream_l445 = (! io_input_cmd_payload_first);
  always @(*) begin
    cmdStage_valid = cmdFork_valid;
    if(when_Stream_l445) begin
      cmdStage_valid = 1'b0;
    end
  end

  always @(*) begin
    cmdFork_ready = cmdStage_ready;
    if(when_Stream_l445) begin
      cmdFork_ready = 1'b1;
    end
  end

  assign cmdStage_payload_last = cmdFork_payload_last;
  assign cmdStage_payload_fragment_source = cmdFork_payload_fragment_source;
  assign cmdStage_payload_fragment_opcode = cmdFork_payload_fragment_opcode;
  assign cmdStage_payload_fragment_address = cmdFork_payload_fragment_address;
  assign cmdStage_payload_fragment_length = cmdFork_payload_fragment_length;
  assign cmdStage_payload_fragment_data = cmdFork_payload_fragment_data;
  assign cmdStage_payload_fragment_mask = cmdFork_payload_fragment_mask;
  assign cmdStage_payload_fragment_context = cmdFork_payload_fragment_context;
  assign when_Stream_l445_1 = (! (dataFork_payload_fragment_opcode == 1'b1));
  always @(*) begin
    dataStage_valid = dataFork_valid;
    if(when_Stream_l445_1) begin
      dataStage_valid = 1'b0;
    end
  end

  always @(*) begin
    dataFork_ready = dataStage_ready;
    if(when_Stream_l445_1) begin
      dataFork_ready = 1'b1;
    end
  end

  assign dataStage_payload_last = dataFork_payload_last;
  assign dataStage_payload_fragment_source = dataFork_payload_fragment_source;
  assign dataStage_payload_fragment_opcode = dataFork_payload_fragment_opcode;
  assign dataStage_payload_fragment_address = dataFork_payload_fragment_address;
  assign dataStage_payload_fragment_length = dataFork_payload_fragment_length;
  assign dataStage_payload_fragment_data = dataFork_payload_fragment_data;
  assign dataStage_payload_fragment_mask = dataFork_payload_fragment_mask;
  assign dataStage_payload_fragment_context = dataFork_payload_fragment_context;
  assign cmdStage_fire = (cmdStage_valid && cmdStage_ready);
  assign writeCmdInfo_valid = (cmdStage_fire && (cmdStage_payload_fragment_opcode == 1'b1));
  assign writeCmdInfo_payload_source = cmdStage_payload_fragment_source;
  assign writeCmdInfo_payload_context = cmdStage_payload_fragment_context;
  assign readCmdInfo_valid = (cmdStage_fire && (cmdStage_payload_fragment_opcode == 1'b0));
  assign readCmdInfo_payload_source = cmdStage_payload_fragment_source;
  assign readCmdInfo_payload_context = cmdStage_payload_fragment_context;
  assign writeCmdInfo_ready = writeCmdInfo_fifo_io_push_ready;
  assign writeRspInfo_fire = (writeRspInfo_valid && writeRspInfo_ready);
  assign writeCmdInfo_fifo_io_pop_ready = (! writeCmdInfo_fifo_io_pop_rValid);
  assign writeRspInfo_valid = writeCmdInfo_fifo_io_pop_rValid;
  assign writeRspInfo_payload_source = writeCmdInfo_fifo_io_pop_rData_source;
  assign writeRspInfo_payload_context = writeCmdInfo_fifo_io_pop_rData_context;
  assign readCmdInfo_ready = readCmdInfo_fifo_io_push_ready;
  assign readRspInfo_fire = (readRspInfo_valid && readRspInfo_ready);
  assign readCmdInfo_fifo_io_pop_ready = (! readCmdInfo_fifo_io_pop_rValid);
  assign readRspInfo_valid = readCmdInfo_fifo_io_pop_rValid;
  assign readRspInfo_payload_source = readCmdInfo_fifo_io_pop_rData_source;
  assign readRspInfo_payload_context = readCmdInfo_fifo_io_pop_rData_context;
  assign _zz_io_output_arw_valid = (! ((! writeCmdInfo_ready) || (! readCmdInfo_ready)));
  assign cmdStage_ready = (io_output_arw_ready && _zz_io_output_arw_valid);
  assign io_output_arw_valid = (cmdStage_valid && _zz_io_output_arw_valid);
  assign io_output_arw_payload_write = (io_input_cmd_payload_fragment_opcode == 1'b1);
  assign io_output_arw_payload_addr = io_input_cmd_payload_fragment_address;
  assign io_output_arw_payload_len = {4'd0, _zz_io_output_arw_payload_len};
  assign io_output_arw_payload_size = 3'b010;
  assign io_output_arw_payload_prot = 3'b010;
  assign io_output_arw_payload_cache = 4'b1111;
  assign io_output_w_valid = dataStage_valid;
  assign dataStage_ready = io_output_w_ready;
  assign io_output_w_payload_data = dataStage_payload_fragment_data;
  assign io_output_w_payload_strb = dataStage_payload_fragment_mask;
  assign io_output_w_payload_last = dataStage_payload_last;
  assign when_BmbToAxi4Bridge_l87 = (io_output_r_valid || io_output_b_valid);
  assign io_output_r_fire = (io_output_r_valid && io_output_r_ready);
  assign io_output_b_fire = (io_output_b_valid && io_output_b_ready);
  assign when_BmbToAxi4Bridge_l87_1 = ((io_output_r_fire && io_output_r_payload_last) || io_output_b_fire);
  assign when_BmbToAxi4Bridge_l88 = (! rspSelLock);
  assign rspSelRead = (rspSelLock ? rspSelReadLast : io_output_r_valid);
  assign io_output_b_ready = ((io_input_rsp_ready && (! rspSelRead)) && writeRspInfo_valid);
  assign io_output_r_ready = ((io_input_rsp_ready && rspSelRead) && readRspInfo_valid);
  assign writeRspInfo_ready = ((io_input_rsp_fire && io_input_rsp_payload_last) && (! rspSelRead));
  assign readRspInfo_ready = ((io_input_rsp_fire && io_input_rsp_payload_last) && rspSelRead);
  assign io_input_rsp_payload_fragment_data = io_output_r_payload_data;
  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_valid = (io_output_r_valid && readRspInfo_valid);
    end else begin
      io_input_rsp_valid = (io_output_b_valid && writeRspInfo_valid);
    end
  end

  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_payload_last = io_output_r_payload_last;
    end else begin
      io_input_rsp_payload_last = 1'b1;
    end
  end

  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_payload_fragment_source = readRspInfo_payload_source;
    end else begin
      io_input_rsp_payload_fragment_source = writeRspInfo_payload_source;
    end
  end

  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_payload_fragment_context = readRspInfo_payload_context;
    end else begin
      io_input_rsp_payload_fragment_context = writeRspInfo_payload_context;
    end
  end

  assign when_BmbToAxi4Bridge_l108 = (rspSelRead ? (io_output_r_payload_resp == 2'b00) : (io_output_b_payload_resp == 2'b00));
  always @(*) begin
    if(when_BmbToAxi4Bridge_l108) begin
      io_input_rsp_payload_fragment_opcode = 1'b0;
    end else begin
      io_input_rsp_payload_fragment_opcode = 1'b1;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      states_0_counter_value <= 3'b000;
      states_1_counter_value <= 3'b000;
      states_2_counter_value <= 3'b000;
      states_3_counter_value <= 3'b000;
      _zz_cmdFork_valid_1 <= 1'b1;
      _zz_dataFork_valid <= 1'b1;
      io_input_cmd_payload_first <= 1'b1;
      writeCmdInfo_fifo_io_pop_rValid <= 1'b0;
      readCmdInfo_fifo_io_pop_rValid <= 1'b0;
      rspSelLock <= 1'b0;
    end else begin
      states_0_counter_value <= states_0_counter_valueNext;
      states_1_counter_value <= states_1_counter_valueNext;
      states_2_counter_value <= states_2_counter_valueNext;
      states_3_counter_value <= states_3_counter_valueNext;
      if(cmdFork_fire) begin
        _zz_cmdFork_valid_1 <= 1'b0;
      end
      if(dataFork_fire) begin
        _zz_dataFork_valid <= 1'b0;
      end
      if(_zz_io_input_cmd_ready_1) begin
        _zz_cmdFork_valid_1 <= 1'b1;
        _zz_dataFork_valid <= 1'b1;
      end
      if(io_input_cmd_fire) begin
        io_input_cmd_payload_first <= io_input_cmd_payload_last;
      end
      if(writeCmdInfo_fifo_io_pop_valid) begin
        writeCmdInfo_fifo_io_pop_rValid <= 1'b1;
      end
      if(writeRspInfo_fire) begin
        writeCmdInfo_fifo_io_pop_rValid <= 1'b0;
      end
      if(readCmdInfo_fifo_io_pop_valid) begin
        readCmdInfo_fifo_io_pop_rValid <= 1'b1;
      end
      if(readRspInfo_fire) begin
        readCmdInfo_fifo_io_pop_rValid <= 1'b0;
      end
      if(when_BmbToAxi4Bridge_l87) begin
        rspSelLock <= 1'b1;
      end
      if(when_BmbToAxi4Bridge_l87_1) begin
        rspSelLock <= 1'b0;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(when_BmbToAxi4Bridge_l45) begin
      states_0_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(when_BmbToAxi4Bridge_l45_1) begin
      states_1_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(when_BmbToAxi4Bridge_l45_2) begin
      states_2_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(when_BmbToAxi4Bridge_l45_3) begin
      states_3_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(writeCmdInfo_fifo_io_pop_ready) begin
      writeCmdInfo_fifo_io_pop_rData_source <= writeCmdInfo_fifo_io_pop_payload_source;
      writeCmdInfo_fifo_io_pop_rData_context <= writeCmdInfo_fifo_io_pop_payload_context;
    end
    if(readCmdInfo_fifo_io_pop_ready) begin
      readCmdInfo_fifo_io_pop_rData_source <= readCmdInfo_fifo_io_pop_payload_source;
      readCmdInfo_fifo_io_pop_rData_context <= readCmdInfo_fifo_io_pop_payload_context;
    end
    if(when_BmbToAxi4Bridge_l88) begin
      rspSelReadLast <= io_output_r_valid;
    end
  end


endmodule

module StreamFifoLowLatency_1 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [7:0]    io_push_payload_len,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [7:0]    io_pop_payload_len,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_ddrAReset_reset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [7:0]    fifo_io_pop_payload_len;
  wire       [2:0]    fifo_io_occupancy;
  wire       [2:0]    fifo_io_availability;

  StreamFifo_6 fifo (
    .io_push_valid                       (io_push_valid                      ), //i
    .io_push_ready                       (fifo_io_push_ready                 ), //o
    .io_push_payload_len                 (io_push_payload_len[7:0]           ), //i
    .io_pop_valid                        (fifo_io_pop_valid                  ), //o
    .io_pop_ready                        (io_pop_ready                       ), //i
    .io_pop_payload_len                  (fifo_io_pop_payload_len[7:0]       ), //o
    .io_flush                            (io_flush                           ), //i
    .io_occupancy                        (fifo_io_occupancy[2:0]             ), //o
    .io_availability                     (fifo_io_availability[2:0]          ), //o
    .io_memoryClk                        (io_memoryClk                       ), //i
    .system_ddr_ddrLogic_ddrAReset_reset (system_ddr_ddrLogic_ddrAReset_reset)  //i
  );
  assign io_push_ready = fifo_io_push_ready;
  assign io_pop_valid = fifo_io_pop_valid;
  assign io_pop_payload_len = fifo_io_pop_payload_len;
  assign io_occupancy = fifo_io_occupancy;
  assign io_availability = fifo_io_availability;

endmodule

module Axi4Upsizer_1 (
  input  wire          io_input_aw_valid,
  output wire          io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [3:0]    io_input_aw_payload_region,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire [0:0]    io_input_aw_payload_lock,
  input  wire [3:0]    io_input_aw_payload_cache,
  input  wire [3:0]    io_input_aw_payload_qos,
  input  wire [2:0]    io_input_aw_payload_prot,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [63:0]   io_input_w_payload_data,
  input  wire [7:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output wire [3:0]    io_input_b_payload_id,
  output wire [1:0]    io_input_b_payload_resp,
  input  wire          io_input_ar_valid,
  output wire          io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [3:0]    io_input_ar_payload_region,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  input  wire [0:0]    io_input_ar_payload_lock,
  input  wire [3:0]    io_input_ar_payload_cache,
  input  wire [3:0]    io_input_ar_payload_qos,
  input  wire [2:0]    io_input_ar_payload_prot,
  output wire          io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [63:0]   io_input_r_payload_data,
  output wire [3:0]    io_input_r_payload_id,
  output wire [1:0]    io_input_r_payload_resp,
  output wire          io_input_r_payload_last,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [3:0]    io_output_aw_payload_id,
  output wire [3:0]    io_output_aw_payload_region,
  output wire [7:0]    io_output_aw_payload_len,
  output wire [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire [0:0]    io_output_aw_payload_lock,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [3:0]    io_output_aw_payload_qos,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [127:0]  io_output_w_payload_data,
  output wire [15:0]   io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [3:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [3:0]    io_output_ar_payload_id,
  output wire [3:0]    io_output_ar_payload_region,
  output wire [7:0]    io_output_ar_payload_len,
  output wire [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  output wire [0:0]    io_output_ar_payload_lock,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [3:0]    io_output_ar_payload_qos,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [127:0]  io_output_r_payload_data,
  input  wire [3:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                readOnly_io_input_ar_ready;
  wire                readOnly_io_input_r_valid;
  wire       [63:0]   readOnly_io_input_r_payload_data;
  wire       [3:0]    readOnly_io_input_r_payload_id;
  wire       [1:0]    readOnly_io_input_r_payload_resp;
  wire                readOnly_io_input_r_payload_last;
  wire                readOnly_io_output_ar_valid;
  wire       [31:0]   readOnly_io_output_ar_payload_addr;
  wire       [3:0]    readOnly_io_output_ar_payload_id;
  wire       [3:0]    readOnly_io_output_ar_payload_region;
  wire       [7:0]    readOnly_io_output_ar_payload_len;
  wire       [2:0]    readOnly_io_output_ar_payload_size;
  wire       [1:0]    readOnly_io_output_ar_payload_burst;
  wire       [0:0]    readOnly_io_output_ar_payload_lock;
  wire       [3:0]    readOnly_io_output_ar_payload_cache;
  wire       [3:0]    readOnly_io_output_ar_payload_qos;
  wire       [2:0]    readOnly_io_output_ar_payload_prot;
  wire                readOnly_io_output_r_ready;
  wire                writeOnly_io_input_aw_ready;
  wire                writeOnly_io_input_w_ready;
  wire                writeOnly_io_input_b_valid;
  wire       [3:0]    writeOnly_io_input_b_payload_id;
  wire       [1:0]    writeOnly_io_input_b_payload_resp;
  wire                writeOnly_io_output_aw_valid;
  wire       [31:0]   writeOnly_io_output_aw_payload_addr;
  wire       [3:0]    writeOnly_io_output_aw_payload_id;
  wire       [3:0]    writeOnly_io_output_aw_payload_region;
  wire       [7:0]    writeOnly_io_output_aw_payload_len;
  wire       [2:0]    writeOnly_io_output_aw_payload_size;
  wire       [1:0]    writeOnly_io_output_aw_payload_burst;
  wire       [0:0]    writeOnly_io_output_aw_payload_lock;
  wire       [3:0]    writeOnly_io_output_aw_payload_cache;
  wire       [3:0]    writeOnly_io_output_aw_payload_qos;
  wire       [2:0]    writeOnly_io_output_aw_payload_prot;
  wire                writeOnly_io_output_w_valid;
  wire       [127:0]  writeOnly_io_output_w_payload_data;
  wire       [15:0]   writeOnly_io_output_w_payload_strb;
  wire                writeOnly_io_output_w_payload_last;
  wire                writeOnly_io_output_b_ready;

  Axi4ReadOnlyUpsizer_1 readOnly (
    .io_input_ar_valid           (io_input_ar_valid                        ), //i
    .io_input_ar_ready           (readOnly_io_input_ar_ready               ), //o
    .io_input_ar_payload_addr    (io_input_ar_payload_addr[31:0]           ), //i
    .io_input_ar_payload_id      (io_input_ar_payload_id[3:0]              ), //i
    .io_input_ar_payload_region  (io_input_ar_payload_region[3:0]          ), //i
    .io_input_ar_payload_len     (io_input_ar_payload_len[7:0]             ), //i
    .io_input_ar_payload_size    (io_input_ar_payload_size[2:0]            ), //i
    .io_input_ar_payload_burst   (io_input_ar_payload_burst[1:0]           ), //i
    .io_input_ar_payload_lock    (io_input_ar_payload_lock                 ), //i
    .io_input_ar_payload_cache   (io_input_ar_payload_cache[3:0]           ), //i
    .io_input_ar_payload_qos     (io_input_ar_payload_qos[3:0]             ), //i
    .io_input_ar_payload_prot    (io_input_ar_payload_prot[2:0]            ), //i
    .io_input_r_valid            (readOnly_io_input_r_valid                ), //o
    .io_input_r_ready            (io_input_r_ready                         ), //i
    .io_input_r_payload_data     (readOnly_io_input_r_payload_data[63:0]   ), //o
    .io_input_r_payload_id       (readOnly_io_input_r_payload_id[3:0]      ), //o
    .io_input_r_payload_resp     (readOnly_io_input_r_payload_resp[1:0]    ), //o
    .io_input_r_payload_last     (readOnly_io_input_r_payload_last         ), //o
    .io_output_ar_valid          (readOnly_io_output_ar_valid              ), //o
    .io_output_ar_ready          (io_output_ar_ready                       ), //i
    .io_output_ar_payload_addr   (readOnly_io_output_ar_payload_addr[31:0] ), //o
    .io_output_ar_payload_id     (readOnly_io_output_ar_payload_id[3:0]    ), //o
    .io_output_ar_payload_region (readOnly_io_output_ar_payload_region[3:0]), //o
    .io_output_ar_payload_len    (readOnly_io_output_ar_payload_len[7:0]   ), //o
    .io_output_ar_payload_size   (readOnly_io_output_ar_payload_size[2:0]  ), //o
    .io_output_ar_payload_burst  (readOnly_io_output_ar_payload_burst[1:0] ), //o
    .io_output_ar_payload_lock   (readOnly_io_output_ar_payload_lock       ), //o
    .io_output_ar_payload_cache  (readOnly_io_output_ar_payload_cache[3:0] ), //o
    .io_output_ar_payload_qos    (readOnly_io_output_ar_payload_qos[3:0]   ), //o
    .io_output_ar_payload_prot   (readOnly_io_output_ar_payload_prot[2:0]  ), //o
    .io_output_r_valid           (io_output_r_valid                        ), //i
    .io_output_r_ready           (readOnly_io_output_r_ready               ), //o
    .io_output_r_payload_data    (io_output_r_payload_data[127:0]          ), //i
    .io_output_r_payload_id      (io_output_r_payload_id[3:0]              ), //i
    .io_output_r_payload_resp    (io_output_r_payload_resp[1:0]            ), //i
    .io_output_r_payload_last    (io_output_r_payload_last                 ), //i
    .io_memoryClk                (io_memoryClk                             ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                  )  //i
  );
  Axi4WriteOnlyUpsizer_1 writeOnly (
    .io_input_aw_valid           (io_input_aw_valid                         ), //i
    .io_input_aw_ready           (writeOnly_io_input_aw_ready               ), //o
    .io_input_aw_payload_addr    (io_input_aw_payload_addr[31:0]            ), //i
    .io_input_aw_payload_id      (io_input_aw_payload_id[3:0]               ), //i
    .io_input_aw_payload_region  (io_input_aw_payload_region[3:0]           ), //i
    .io_input_aw_payload_len     (io_input_aw_payload_len[7:0]              ), //i
    .io_input_aw_payload_size    (io_input_aw_payload_size[2:0]             ), //i
    .io_input_aw_payload_burst   (io_input_aw_payload_burst[1:0]            ), //i
    .io_input_aw_payload_lock    (io_input_aw_payload_lock                  ), //i
    .io_input_aw_payload_cache   (io_input_aw_payload_cache[3:0]            ), //i
    .io_input_aw_payload_qos     (io_input_aw_payload_qos[3:0]              ), //i
    .io_input_aw_payload_prot    (io_input_aw_payload_prot[2:0]             ), //i
    .io_input_w_valid            (io_input_w_valid                          ), //i
    .io_input_w_ready            (writeOnly_io_input_w_ready                ), //o
    .io_input_w_payload_data     (io_input_w_payload_data[63:0]             ), //i
    .io_input_w_payload_strb     (io_input_w_payload_strb[7:0]              ), //i
    .io_input_w_payload_last     (io_input_w_payload_last                   ), //i
    .io_input_b_valid            (writeOnly_io_input_b_valid                ), //o
    .io_input_b_ready            (io_input_b_ready                          ), //i
    .io_input_b_payload_id       (writeOnly_io_input_b_payload_id[3:0]      ), //o
    .io_input_b_payload_resp     (writeOnly_io_input_b_payload_resp[1:0]    ), //o
    .io_output_aw_valid          (writeOnly_io_output_aw_valid              ), //o
    .io_output_aw_ready          (io_output_aw_ready                        ), //i
    .io_output_aw_payload_addr   (writeOnly_io_output_aw_payload_addr[31:0] ), //o
    .io_output_aw_payload_id     (writeOnly_io_output_aw_payload_id[3:0]    ), //o
    .io_output_aw_payload_region (writeOnly_io_output_aw_payload_region[3:0]), //o
    .io_output_aw_payload_len    (writeOnly_io_output_aw_payload_len[7:0]   ), //o
    .io_output_aw_payload_size   (writeOnly_io_output_aw_payload_size[2:0]  ), //o
    .io_output_aw_payload_burst  (writeOnly_io_output_aw_payload_burst[1:0] ), //o
    .io_output_aw_payload_lock   (writeOnly_io_output_aw_payload_lock       ), //o
    .io_output_aw_payload_cache  (writeOnly_io_output_aw_payload_cache[3:0] ), //o
    .io_output_aw_payload_qos    (writeOnly_io_output_aw_payload_qos[3:0]   ), //o
    .io_output_aw_payload_prot   (writeOnly_io_output_aw_payload_prot[2:0]  ), //o
    .io_output_w_valid           (writeOnly_io_output_w_valid               ), //o
    .io_output_w_ready           (io_output_w_ready                         ), //i
    .io_output_w_payload_data    (writeOnly_io_output_w_payload_data[127:0] ), //o
    .io_output_w_payload_strb    (writeOnly_io_output_w_payload_strb[15:0]  ), //o
    .io_output_w_payload_last    (writeOnly_io_output_w_payload_last        ), //o
    .io_output_b_valid           (io_output_b_valid                         ), //i
    .io_output_b_ready           (writeOnly_io_output_b_ready               ), //o
    .io_output_b_payload_id      (io_output_b_payload_id[3:0]               ), //i
    .io_output_b_payload_resp    (io_output_b_payload_resp[1:0]             ), //i
    .io_memoryClk                (io_memoryClk                              ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                   )  //i
  );
  assign io_input_ar_ready = readOnly_io_input_ar_ready;
  assign io_input_r_valid = readOnly_io_input_r_valid;
  assign io_input_r_payload_data = readOnly_io_input_r_payload_data;
  assign io_input_r_payload_id = readOnly_io_input_r_payload_id;
  assign io_input_r_payload_resp = readOnly_io_input_r_payload_resp;
  assign io_input_r_payload_last = readOnly_io_input_r_payload_last;
  assign io_input_aw_ready = writeOnly_io_input_aw_ready;
  assign io_input_w_ready = writeOnly_io_input_w_ready;
  assign io_input_b_valid = writeOnly_io_input_b_valid;
  assign io_input_b_payload_id = writeOnly_io_input_b_payload_id;
  assign io_input_b_payload_resp = writeOnly_io_input_b_payload_resp;
  assign io_output_ar_valid = readOnly_io_output_ar_valid;
  assign io_output_ar_payload_addr = readOnly_io_output_ar_payload_addr;
  assign io_output_ar_payload_id = readOnly_io_output_ar_payload_id;
  assign io_output_ar_payload_region = readOnly_io_output_ar_payload_region;
  assign io_output_ar_payload_len = readOnly_io_output_ar_payload_len;
  assign io_output_ar_payload_size = readOnly_io_output_ar_payload_size;
  assign io_output_ar_payload_burst = readOnly_io_output_ar_payload_burst;
  assign io_output_ar_payload_lock = readOnly_io_output_ar_payload_lock;
  assign io_output_ar_payload_cache = readOnly_io_output_ar_payload_cache;
  assign io_output_ar_payload_qos = readOnly_io_output_ar_payload_qos;
  assign io_output_ar_payload_prot = readOnly_io_output_ar_payload_prot;
  assign io_output_r_ready = readOnly_io_output_r_ready;
  assign io_output_aw_valid = writeOnly_io_output_aw_valid;
  assign io_output_aw_payload_addr = writeOnly_io_output_aw_payload_addr;
  assign io_output_aw_payload_id = writeOnly_io_output_aw_payload_id;
  assign io_output_aw_payload_region = writeOnly_io_output_aw_payload_region;
  assign io_output_aw_payload_len = writeOnly_io_output_aw_payload_len;
  assign io_output_aw_payload_size = writeOnly_io_output_aw_payload_size;
  assign io_output_aw_payload_burst = writeOnly_io_output_aw_payload_burst;
  assign io_output_aw_payload_lock = writeOnly_io_output_aw_payload_lock;
  assign io_output_aw_payload_cache = writeOnly_io_output_aw_payload_cache;
  assign io_output_aw_payload_qos = writeOnly_io_output_aw_payload_qos;
  assign io_output_aw_payload_prot = writeOnly_io_output_aw_payload_prot;
  assign io_output_w_valid = writeOnly_io_output_w_valid;
  assign io_output_w_payload_data = writeOnly_io_output_w_payload_data;
  assign io_output_w_payload_strb = writeOnly_io_output_w_payload_strb;
  assign io_output_w_payload_last = writeOnly_io_output_w_payload_last;
  assign io_output_b_ready = writeOnly_io_output_b_ready;

endmodule

module Axi4CC_1 (
  input  wire          io_input_aw_valid,
  output wire          io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [3:0]    io_input_aw_payload_region,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire [0:0]    io_input_aw_payload_lock,
  input  wire [3:0]    io_input_aw_payload_cache,
  input  wire [3:0]    io_input_aw_payload_qos,
  input  wire [2:0]    io_input_aw_payload_prot,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [63:0]   io_input_w_payload_data,
  input  wire [7:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output wire [3:0]    io_input_b_payload_id,
  output wire [1:0]    io_input_b_payload_resp,
  input  wire          io_input_ar_valid,
  output wire          io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [3:0]    io_input_ar_payload_region,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  input  wire [0:0]    io_input_ar_payload_lock,
  input  wire [3:0]    io_input_ar_payload_cache,
  input  wire [3:0]    io_input_ar_payload_qos,
  input  wire [2:0]    io_input_ar_payload_prot,
  output wire          io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [63:0]   io_input_r_payload_data,
  output wire [3:0]    io_input_r_payload_id,
  output wire [1:0]    io_input_r_payload_resp,
  output wire          io_input_r_payload_last,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [3:0]    io_output_aw_payload_id,
  output wire [3:0]    io_output_aw_payload_region,
  output wire [7:0]    io_output_aw_payload_len,
  output wire [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire [0:0]    io_output_aw_payload_lock,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [3:0]    io_output_aw_payload_qos,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [63:0]   io_output_w_payload_data,
  output wire [7:0]    io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [3:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [3:0]    io_output_ar_payload_id,
  output wire [3:0]    io_output_ar_payload_region,
  output wire [7:0]    io_output_ar_payload_len,
  output wire [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  output wire [0:0]    io_output_ar_payload_lock,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [3:0]    io_output_ar_payload_qos,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [63:0]   io_output_r_payload_data,
  input  wire [3:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_ddrMasters_0_clk,
  input  wire          io_ddrMasters_0_reset,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                io_input_ar_queue_io_push_ready;
  wire                io_input_ar_queue_io_pop_valid;
  wire       [31:0]   io_input_ar_queue_io_pop_payload_addr;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_id;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_region;
  wire       [7:0]    io_input_ar_queue_io_pop_payload_len;
  wire       [2:0]    io_input_ar_queue_io_pop_payload_size;
  wire       [1:0]    io_input_ar_queue_io_pop_payload_burst;
  wire       [0:0]    io_input_ar_queue_io_pop_payload_lock;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_cache;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_qos;
  wire       [2:0]    io_input_ar_queue_io_pop_payload_prot;
  wire       [4:0]    io_input_ar_queue_io_pushOccupancy;
  wire       [4:0]    io_input_ar_queue_io_popOccupancy;
  wire                io_input_ar_queue_system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1;
  wire                io_output_r_queue_io_push_ready;
  wire                io_output_r_queue_io_pop_valid;
  wire       [63:0]   io_output_r_queue_io_pop_payload_data;
  wire       [3:0]    io_output_r_queue_io_pop_payload_id;
  wire       [1:0]    io_output_r_queue_io_pop_payload_resp;
  wire                io_output_r_queue_io_pop_payload_last;
  wire       [4:0]    io_output_r_queue_io_pushOccupancy;
  wire       [4:0]    io_output_r_queue_io_popOccupancy;
  wire                io_output_r_queue_system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1;
  wire                io_input_aw_queue_io_push_ready;
  wire                io_input_aw_queue_io_pop_valid;
  wire       [31:0]   io_input_aw_queue_io_pop_payload_addr;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_id;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_region;
  wire       [7:0]    io_input_aw_queue_io_pop_payload_len;
  wire       [2:0]    io_input_aw_queue_io_pop_payload_size;
  wire       [1:0]    io_input_aw_queue_io_pop_payload_burst;
  wire       [0:0]    io_input_aw_queue_io_pop_payload_lock;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_cache;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_qos;
  wire       [2:0]    io_input_aw_queue_io_pop_payload_prot;
  wire       [4:0]    io_input_aw_queue_io_pushOccupancy;
  wire       [4:0]    io_input_aw_queue_io_popOccupancy;
  wire                io_input_w_queue_io_push_ready;
  wire                io_input_w_queue_io_pop_valid;
  wire       [63:0]   io_input_w_queue_io_pop_payload_data;
  wire       [7:0]    io_input_w_queue_io_pop_payload_strb;
  wire                io_input_w_queue_io_pop_payload_last;
  wire       [4:0]    io_input_w_queue_io_pushOccupancy;
  wire       [4:0]    io_input_w_queue_io_popOccupancy;
  wire                io_output_b_queue_io_push_ready;
  wire                io_output_b_queue_io_pop_valid;
  wire       [3:0]    io_output_b_queue_io_pop_payload_id;
  wire       [1:0]    io_output_b_queue_io_pop_payload_resp;
  wire       [4:0]    io_output_b_queue_io_pushOccupancy;
  wire       [4:0]    io_output_b_queue_io_popOccupancy;

  StreamFifoCC_7 io_input_ar_queue (
    .io_push_valid                                                                           (io_input_ar_valid                                                                                        ), //i
    .io_push_ready                                                                           (io_input_ar_queue_io_push_ready                                                                          ), //o
    .io_push_payload_addr                                                                    (io_input_ar_payload_addr[31:0]                                                                           ), //i
    .io_push_payload_id                                                                      (io_input_ar_payload_id[3:0]                                                                              ), //i
    .io_push_payload_region                                                                  (io_input_ar_payload_region[3:0]                                                                          ), //i
    .io_push_payload_len                                                                     (io_input_ar_payload_len[7:0]                                                                             ), //i
    .io_push_payload_size                                                                    (io_input_ar_payload_size[2:0]                                                                            ), //i
    .io_push_payload_burst                                                                   (io_input_ar_payload_burst[1:0]                                                                           ), //i
    .io_push_payload_lock                                                                    (io_input_ar_payload_lock                                                                                 ), //i
    .io_push_payload_cache                                                                   (io_input_ar_payload_cache[3:0]                                                                           ), //i
    .io_push_payload_qos                                                                     (io_input_ar_payload_qos[3:0]                                                                             ), //i
    .io_push_payload_prot                                                                    (io_input_ar_payload_prot[2:0]                                                                            ), //i
    .io_pop_valid                                                                            (io_input_ar_queue_io_pop_valid                                                                           ), //o
    .io_pop_ready                                                                            (io_output_ar_ready                                                                                       ), //i
    .io_pop_payload_addr                                                                     (io_input_ar_queue_io_pop_payload_addr[31:0]                                                              ), //o
    .io_pop_payload_id                                                                       (io_input_ar_queue_io_pop_payload_id[3:0]                                                                 ), //o
    .io_pop_payload_region                                                                   (io_input_ar_queue_io_pop_payload_region[3:0]                                                             ), //o
    .io_pop_payload_len                                                                      (io_input_ar_queue_io_pop_payload_len[7:0]                                                                ), //o
    .io_pop_payload_size                                                                     (io_input_ar_queue_io_pop_payload_size[2:0]                                                               ), //o
    .io_pop_payload_burst                                                                    (io_input_ar_queue_io_pop_payload_burst[1:0]                                                              ), //o
    .io_pop_payload_lock                                                                     (io_input_ar_queue_io_pop_payload_lock                                                                    ), //o
    .io_pop_payload_cache                                                                    (io_input_ar_queue_io_pop_payload_cache[3:0]                                                              ), //o
    .io_pop_payload_qos                                                                      (io_input_ar_queue_io_pop_payload_qos[3:0]                                                                ), //o
    .io_pop_payload_prot                                                                     (io_input_ar_queue_io_pop_payload_prot[2:0]                                                               ), //o
    .io_pushOccupancy                                                                        (io_input_ar_queue_io_pushOccupancy[4:0]                                                                  ), //o
    .io_popOccupancy                                                                         (io_input_ar_queue_io_popOccupancy[4:0]                                                                   ), //o
    .io_ddrMasters_0_clk                                                                     (io_ddrMasters_0_clk                                                                                      ), //i
    .io_ddrMasters_0_reset                                                                   (io_ddrMasters_0_reset                                                                                    ), //i
    .io_memoryClk                                                                            (io_memoryClk                                                                                             ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1 (io_input_ar_queue_system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1)  //o
  );
  StreamFifoCC_8 io_output_r_queue (
    .io_push_valid                                                                             (io_output_r_valid                                                                                          ), //i
    .io_push_ready                                                                             (io_output_r_queue_io_push_ready                                                                            ), //o
    .io_push_payload_data                                                                      (io_output_r_payload_data[63:0]                                                                             ), //i
    .io_push_payload_id                                                                        (io_output_r_payload_id[3:0]                                                                                ), //i
    .io_push_payload_resp                                                                      (io_output_r_payload_resp[1:0]                                                                              ), //i
    .io_push_payload_last                                                                      (io_output_r_payload_last                                                                                   ), //i
    .io_pop_valid                                                                              (io_output_r_queue_io_pop_valid                                                                             ), //o
    .io_pop_ready                                                                              (io_input_r_ready                                                                                           ), //i
    .io_pop_payload_data                                                                       (io_output_r_queue_io_pop_payload_data[63:0]                                                                ), //o
    .io_pop_payload_id                                                                         (io_output_r_queue_io_pop_payload_id[3:0]                                                                   ), //o
    .io_pop_payload_resp                                                                       (io_output_r_queue_io_pop_payload_resp[1:0]                                                                 ), //o
    .io_pop_payload_last                                                                       (io_output_r_queue_io_pop_payload_last                                                                      ), //o
    .io_pushOccupancy                                                                          (io_output_r_queue_io_pushOccupancy[4:0]                                                                    ), //o
    .io_popOccupancy                                                                           (io_output_r_queue_io_popOccupancy[4:0]                                                                     ), //o
    .io_memoryClk                                                                              (io_memoryClk                                                                                               ), //i
    .ddrCd_logic_outputReset                                                                   (ddrCd_logic_outputReset                                                                                    ), //i
    .io_ddrMasters_0_clk                                                                       (io_ddrMasters_0_clk                                                                                        ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 (io_output_r_queue_system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1)  //o
  );
  StreamFifoCC_9 io_input_aw_queue (
    .io_push_valid                                                                           (io_input_aw_valid                                                                                        ), //i
    .io_push_ready                                                                           (io_input_aw_queue_io_push_ready                                                                          ), //o
    .io_push_payload_addr                                                                    (io_input_aw_payload_addr[31:0]                                                                           ), //i
    .io_push_payload_id                                                                      (io_input_aw_payload_id[3:0]                                                                              ), //i
    .io_push_payload_region                                                                  (io_input_aw_payload_region[3:0]                                                                          ), //i
    .io_push_payload_len                                                                     (io_input_aw_payload_len[7:0]                                                                             ), //i
    .io_push_payload_size                                                                    (io_input_aw_payload_size[2:0]                                                                            ), //i
    .io_push_payload_burst                                                                   (io_input_aw_payload_burst[1:0]                                                                           ), //i
    .io_push_payload_lock                                                                    (io_input_aw_payload_lock                                                                                 ), //i
    .io_push_payload_cache                                                                   (io_input_aw_payload_cache[3:0]                                                                           ), //i
    .io_push_payload_qos                                                                     (io_input_aw_payload_qos[3:0]                                                                             ), //i
    .io_push_payload_prot                                                                    (io_input_aw_payload_prot[2:0]                                                                            ), //i
    .io_pop_valid                                                                            (io_input_aw_queue_io_pop_valid                                                                           ), //o
    .io_pop_ready                                                                            (io_output_aw_ready                                                                                       ), //i
    .io_pop_payload_addr                                                                     (io_input_aw_queue_io_pop_payload_addr[31:0]                                                              ), //o
    .io_pop_payload_id                                                                       (io_input_aw_queue_io_pop_payload_id[3:0]                                                                 ), //o
    .io_pop_payload_region                                                                   (io_input_aw_queue_io_pop_payload_region[3:0]                                                             ), //o
    .io_pop_payload_len                                                                      (io_input_aw_queue_io_pop_payload_len[7:0]                                                                ), //o
    .io_pop_payload_size                                                                     (io_input_aw_queue_io_pop_payload_size[2:0]                                                               ), //o
    .io_pop_payload_burst                                                                    (io_input_aw_queue_io_pop_payload_burst[1:0]                                                              ), //o
    .io_pop_payload_lock                                                                     (io_input_aw_queue_io_pop_payload_lock                                                                    ), //o
    .io_pop_payload_cache                                                                    (io_input_aw_queue_io_pop_payload_cache[3:0]                                                              ), //o
    .io_pop_payload_qos                                                                      (io_input_aw_queue_io_pop_payload_qos[3:0]                                                                ), //o
    .io_pop_payload_prot                                                                     (io_input_aw_queue_io_pop_payload_prot[2:0]                                                               ), //o
    .io_pushOccupancy                                                                        (io_input_aw_queue_io_pushOccupancy[4:0]                                                                  ), //o
    .io_popOccupancy                                                                         (io_input_aw_queue_io_popOccupancy[4:0]                                                                   ), //o
    .io_ddrMasters_0_clk                                                                     (io_ddrMasters_0_clk                                                                                      ), //i
    .io_ddrMasters_0_reset                                                                   (io_ddrMasters_0_reset                                                                                    ), //i
    .io_memoryClk                                                                            (io_memoryClk                                                                                             ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1 (io_input_ar_queue_system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1)  //i
  );
  StreamFifoCC_10 io_input_w_queue (
    .io_push_valid                                                                           (io_input_w_valid                                                                                         ), //i
    .io_push_ready                                                                           (io_input_w_queue_io_push_ready                                                                           ), //o
    .io_push_payload_data                                                                    (io_input_w_payload_data[63:0]                                                                            ), //i
    .io_push_payload_strb                                                                    (io_input_w_payload_strb[7:0]                                                                             ), //i
    .io_push_payload_last                                                                    (io_input_w_payload_last                                                                                  ), //i
    .io_pop_valid                                                                            (io_input_w_queue_io_pop_valid                                                                            ), //o
    .io_pop_ready                                                                            (io_output_w_ready                                                                                        ), //i
    .io_pop_payload_data                                                                     (io_input_w_queue_io_pop_payload_data[63:0]                                                               ), //o
    .io_pop_payload_strb                                                                     (io_input_w_queue_io_pop_payload_strb[7:0]                                                                ), //o
    .io_pop_payload_last                                                                     (io_input_w_queue_io_pop_payload_last                                                                     ), //o
    .io_pushOccupancy                                                                        (io_input_w_queue_io_pushOccupancy[4:0]                                                                   ), //o
    .io_popOccupancy                                                                         (io_input_w_queue_io_popOccupancy[4:0]                                                                    ), //o
    .io_ddrMasters_0_clk                                                                     (io_ddrMasters_0_clk                                                                                      ), //i
    .io_ddrMasters_0_reset                                                                   (io_ddrMasters_0_reset                                                                                    ), //i
    .io_memoryClk                                                                            (io_memoryClk                                                                                             ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1 (io_input_ar_queue_system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1)  //i
  );
  StreamFifoCC_11 io_output_b_queue (
    .io_push_valid                                                                             (io_output_b_valid                                                                                          ), //i
    .io_push_ready                                                                             (io_output_b_queue_io_push_ready                                                                            ), //o
    .io_push_payload_id                                                                        (io_output_b_payload_id[3:0]                                                                                ), //i
    .io_push_payload_resp                                                                      (io_output_b_payload_resp[1:0]                                                                              ), //i
    .io_pop_valid                                                                              (io_output_b_queue_io_pop_valid                                                                             ), //o
    .io_pop_ready                                                                              (io_input_b_ready                                                                                           ), //i
    .io_pop_payload_id                                                                         (io_output_b_queue_io_pop_payload_id[3:0]                                                                   ), //o
    .io_pop_payload_resp                                                                       (io_output_b_queue_io_pop_payload_resp[1:0]                                                                 ), //o
    .io_pushOccupancy                                                                          (io_output_b_queue_io_pushOccupancy[4:0]                                                                    ), //o
    .io_popOccupancy                                                                           (io_output_b_queue_io_popOccupancy[4:0]                                                                     ), //o
    .io_memoryClk                                                                              (io_memoryClk                                                                                               ), //i
    .ddrCd_logic_outputReset                                                                   (ddrCd_logic_outputReset                                                                                    ), //i
    .io_ddrMasters_0_clk                                                                       (io_ddrMasters_0_clk                                                                                        ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 (io_output_r_queue_system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1)  //i
  );
  assign io_input_ar_ready = io_input_ar_queue_io_push_ready;
  assign io_output_ar_valid = io_input_ar_queue_io_pop_valid;
  assign io_output_ar_payload_addr = io_input_ar_queue_io_pop_payload_addr;
  assign io_output_ar_payload_id = io_input_ar_queue_io_pop_payload_id;
  assign io_output_ar_payload_region = io_input_ar_queue_io_pop_payload_region;
  assign io_output_ar_payload_len = io_input_ar_queue_io_pop_payload_len;
  assign io_output_ar_payload_size = io_input_ar_queue_io_pop_payload_size;
  assign io_output_ar_payload_burst = io_input_ar_queue_io_pop_payload_burst;
  assign io_output_ar_payload_lock = io_input_ar_queue_io_pop_payload_lock;
  assign io_output_ar_payload_cache = io_input_ar_queue_io_pop_payload_cache;
  assign io_output_ar_payload_qos = io_input_ar_queue_io_pop_payload_qos;
  assign io_output_ar_payload_prot = io_input_ar_queue_io_pop_payload_prot;
  assign io_output_r_ready = io_output_r_queue_io_push_ready;
  assign io_input_r_valid = io_output_r_queue_io_pop_valid;
  assign io_input_r_payload_data = io_output_r_queue_io_pop_payload_data;
  assign io_input_r_payload_id = io_output_r_queue_io_pop_payload_id;
  assign io_input_r_payload_resp = io_output_r_queue_io_pop_payload_resp;
  assign io_input_r_payload_last = io_output_r_queue_io_pop_payload_last;
  assign io_input_aw_ready = io_input_aw_queue_io_push_ready;
  assign io_output_aw_valid = io_input_aw_queue_io_pop_valid;
  assign io_output_aw_payload_addr = io_input_aw_queue_io_pop_payload_addr;
  assign io_output_aw_payload_id = io_input_aw_queue_io_pop_payload_id;
  assign io_output_aw_payload_region = io_input_aw_queue_io_pop_payload_region;
  assign io_output_aw_payload_len = io_input_aw_queue_io_pop_payload_len;
  assign io_output_aw_payload_size = io_input_aw_queue_io_pop_payload_size;
  assign io_output_aw_payload_burst = io_input_aw_queue_io_pop_payload_burst;
  assign io_output_aw_payload_lock = io_input_aw_queue_io_pop_payload_lock;
  assign io_output_aw_payload_cache = io_input_aw_queue_io_pop_payload_cache;
  assign io_output_aw_payload_qos = io_input_aw_queue_io_pop_payload_qos;
  assign io_output_aw_payload_prot = io_input_aw_queue_io_pop_payload_prot;
  assign io_input_w_ready = io_input_w_queue_io_push_ready;
  assign io_output_w_valid = io_input_w_queue_io_pop_valid;
  assign io_output_w_payload_data = io_input_w_queue_io_pop_payload_data;
  assign io_output_w_payload_strb = io_input_w_queue_io_pop_payload_strb;
  assign io_output_w_payload_last = io_input_w_queue_io_pop_payload_last;
  assign io_output_b_ready = io_output_b_queue_io_push_ready;
  assign io_input_b_valid = io_output_b_queue_io_pop_valid;
  assign io_input_b_payload_id = io_output_b_queue_io_pop_payload_id;
  assign io_input_b_payload_resp = io_output_b_queue_io_pop_payload_resp;

endmodule

module BufferCC_67 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_ddrMasters_0_clk,
  input  wire          io_ddrMasters_0_reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_0_clk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

module Axi4Upsizer (
  input  wire          io_input_aw_valid,
  output wire          io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [3:0]    io_input_aw_payload_region,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire [0:0]    io_input_aw_payload_lock,
  input  wire [3:0]    io_input_aw_payload_cache,
  input  wire [3:0]    io_input_aw_payload_qos,
  input  wire [2:0]    io_input_aw_payload_prot,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [31:0]   io_input_w_payload_data,
  input  wire [3:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output wire [3:0]    io_input_b_payload_id,
  output wire [1:0]    io_input_b_payload_resp,
  input  wire          io_input_ar_valid,
  output wire          io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [3:0]    io_input_ar_payload_region,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  input  wire [0:0]    io_input_ar_payload_lock,
  input  wire [3:0]    io_input_ar_payload_cache,
  input  wire [3:0]    io_input_ar_payload_qos,
  input  wire [2:0]    io_input_ar_payload_prot,
  output wire          io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [31:0]   io_input_r_payload_data,
  output wire [3:0]    io_input_r_payload_id,
  output wire [1:0]    io_input_r_payload_resp,
  output wire          io_input_r_payload_last,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [3:0]    io_output_aw_payload_id,
  output wire [3:0]    io_output_aw_payload_region,
  output wire [7:0]    io_output_aw_payload_len,
  output wire [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire [0:0]    io_output_aw_payload_lock,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [3:0]    io_output_aw_payload_qos,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [127:0]  io_output_w_payload_data,
  output wire [15:0]   io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [3:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [3:0]    io_output_ar_payload_id,
  output wire [3:0]    io_output_ar_payload_region,
  output wire [7:0]    io_output_ar_payload_len,
  output wire [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  output wire [0:0]    io_output_ar_payload_lock,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [3:0]    io_output_ar_payload_qos,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [127:0]  io_output_r_payload_data,
  input  wire [3:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                readOnly_io_input_ar_ready;
  wire                readOnly_io_input_r_valid;
  wire       [31:0]   readOnly_io_input_r_payload_data;
  wire       [3:0]    readOnly_io_input_r_payload_id;
  wire       [1:0]    readOnly_io_input_r_payload_resp;
  wire                readOnly_io_input_r_payload_last;
  wire                readOnly_io_output_ar_valid;
  wire       [31:0]   readOnly_io_output_ar_payload_addr;
  wire       [3:0]    readOnly_io_output_ar_payload_id;
  wire       [3:0]    readOnly_io_output_ar_payload_region;
  wire       [7:0]    readOnly_io_output_ar_payload_len;
  wire       [2:0]    readOnly_io_output_ar_payload_size;
  wire       [1:0]    readOnly_io_output_ar_payload_burst;
  wire       [0:0]    readOnly_io_output_ar_payload_lock;
  wire       [3:0]    readOnly_io_output_ar_payload_cache;
  wire       [3:0]    readOnly_io_output_ar_payload_qos;
  wire       [2:0]    readOnly_io_output_ar_payload_prot;
  wire                readOnly_io_output_r_ready;
  wire                writeOnly_io_input_aw_ready;
  wire                writeOnly_io_input_w_ready;
  wire                writeOnly_io_input_b_valid;
  wire       [3:0]    writeOnly_io_input_b_payload_id;
  wire       [1:0]    writeOnly_io_input_b_payload_resp;
  wire                writeOnly_io_output_aw_valid;
  wire       [31:0]   writeOnly_io_output_aw_payload_addr;
  wire       [3:0]    writeOnly_io_output_aw_payload_id;
  wire       [3:0]    writeOnly_io_output_aw_payload_region;
  wire       [7:0]    writeOnly_io_output_aw_payload_len;
  wire       [2:0]    writeOnly_io_output_aw_payload_size;
  wire       [1:0]    writeOnly_io_output_aw_payload_burst;
  wire       [0:0]    writeOnly_io_output_aw_payload_lock;
  wire       [3:0]    writeOnly_io_output_aw_payload_cache;
  wire       [3:0]    writeOnly_io_output_aw_payload_qos;
  wire       [2:0]    writeOnly_io_output_aw_payload_prot;
  wire                writeOnly_io_output_w_valid;
  wire       [127:0]  writeOnly_io_output_w_payload_data;
  wire       [15:0]   writeOnly_io_output_w_payload_strb;
  wire                writeOnly_io_output_w_payload_last;
  wire                writeOnly_io_output_b_ready;

  Axi4ReadOnlyUpsizer readOnly (
    .io_input_ar_valid           (io_input_ar_valid                        ), //i
    .io_input_ar_ready           (readOnly_io_input_ar_ready               ), //o
    .io_input_ar_payload_addr    (io_input_ar_payload_addr[31:0]           ), //i
    .io_input_ar_payload_id      (io_input_ar_payload_id[3:0]              ), //i
    .io_input_ar_payload_region  (io_input_ar_payload_region[3:0]          ), //i
    .io_input_ar_payload_len     (io_input_ar_payload_len[7:0]             ), //i
    .io_input_ar_payload_size    (io_input_ar_payload_size[2:0]            ), //i
    .io_input_ar_payload_burst   (io_input_ar_payload_burst[1:0]           ), //i
    .io_input_ar_payload_lock    (io_input_ar_payload_lock                 ), //i
    .io_input_ar_payload_cache   (io_input_ar_payload_cache[3:0]           ), //i
    .io_input_ar_payload_qos     (io_input_ar_payload_qos[3:0]             ), //i
    .io_input_ar_payload_prot    (io_input_ar_payload_prot[2:0]            ), //i
    .io_input_r_valid            (readOnly_io_input_r_valid                ), //o
    .io_input_r_ready            (io_input_r_ready                         ), //i
    .io_input_r_payload_data     (readOnly_io_input_r_payload_data[31:0]   ), //o
    .io_input_r_payload_id       (readOnly_io_input_r_payload_id[3:0]      ), //o
    .io_input_r_payload_resp     (readOnly_io_input_r_payload_resp[1:0]    ), //o
    .io_input_r_payload_last     (readOnly_io_input_r_payload_last         ), //o
    .io_output_ar_valid          (readOnly_io_output_ar_valid              ), //o
    .io_output_ar_ready          (io_output_ar_ready                       ), //i
    .io_output_ar_payload_addr   (readOnly_io_output_ar_payload_addr[31:0] ), //o
    .io_output_ar_payload_id     (readOnly_io_output_ar_payload_id[3:0]    ), //o
    .io_output_ar_payload_region (readOnly_io_output_ar_payload_region[3:0]), //o
    .io_output_ar_payload_len    (readOnly_io_output_ar_payload_len[7:0]   ), //o
    .io_output_ar_payload_size   (readOnly_io_output_ar_payload_size[2:0]  ), //o
    .io_output_ar_payload_burst  (readOnly_io_output_ar_payload_burst[1:0] ), //o
    .io_output_ar_payload_lock   (readOnly_io_output_ar_payload_lock       ), //o
    .io_output_ar_payload_cache  (readOnly_io_output_ar_payload_cache[3:0] ), //o
    .io_output_ar_payload_qos    (readOnly_io_output_ar_payload_qos[3:0]   ), //o
    .io_output_ar_payload_prot   (readOnly_io_output_ar_payload_prot[2:0]  ), //o
    .io_output_r_valid           (io_output_r_valid                        ), //i
    .io_output_r_ready           (readOnly_io_output_r_ready               ), //o
    .io_output_r_payload_data    (io_output_r_payload_data[127:0]          ), //i
    .io_output_r_payload_id      (io_output_r_payload_id[3:0]              ), //i
    .io_output_r_payload_resp    (io_output_r_payload_resp[1:0]            ), //i
    .io_output_r_payload_last    (io_output_r_payload_last                 ), //i
    .io_memoryClk                (io_memoryClk                             ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                  )  //i
  );
  Axi4WriteOnlyUpsizer writeOnly (
    .io_input_aw_valid           (io_input_aw_valid                         ), //i
    .io_input_aw_ready           (writeOnly_io_input_aw_ready               ), //o
    .io_input_aw_payload_addr    (io_input_aw_payload_addr[31:0]            ), //i
    .io_input_aw_payload_id      (io_input_aw_payload_id[3:0]               ), //i
    .io_input_aw_payload_region  (io_input_aw_payload_region[3:0]           ), //i
    .io_input_aw_payload_len     (io_input_aw_payload_len[7:0]              ), //i
    .io_input_aw_payload_size    (io_input_aw_payload_size[2:0]             ), //i
    .io_input_aw_payload_burst   (io_input_aw_payload_burst[1:0]            ), //i
    .io_input_aw_payload_lock    (io_input_aw_payload_lock                  ), //i
    .io_input_aw_payload_cache   (io_input_aw_payload_cache[3:0]            ), //i
    .io_input_aw_payload_qos     (io_input_aw_payload_qos[3:0]              ), //i
    .io_input_aw_payload_prot    (io_input_aw_payload_prot[2:0]             ), //i
    .io_input_w_valid            (io_input_w_valid                          ), //i
    .io_input_w_ready            (writeOnly_io_input_w_ready                ), //o
    .io_input_w_payload_data     (io_input_w_payload_data[31:0]             ), //i
    .io_input_w_payload_strb     (io_input_w_payload_strb[3:0]              ), //i
    .io_input_w_payload_last     (io_input_w_payload_last                   ), //i
    .io_input_b_valid            (writeOnly_io_input_b_valid                ), //o
    .io_input_b_ready            (io_input_b_ready                          ), //i
    .io_input_b_payload_id       (writeOnly_io_input_b_payload_id[3:0]      ), //o
    .io_input_b_payload_resp     (writeOnly_io_input_b_payload_resp[1:0]    ), //o
    .io_output_aw_valid          (writeOnly_io_output_aw_valid              ), //o
    .io_output_aw_ready          (io_output_aw_ready                        ), //i
    .io_output_aw_payload_addr   (writeOnly_io_output_aw_payload_addr[31:0] ), //o
    .io_output_aw_payload_id     (writeOnly_io_output_aw_payload_id[3:0]    ), //o
    .io_output_aw_payload_region (writeOnly_io_output_aw_payload_region[3:0]), //o
    .io_output_aw_payload_len    (writeOnly_io_output_aw_payload_len[7:0]   ), //o
    .io_output_aw_payload_size   (writeOnly_io_output_aw_payload_size[2:0]  ), //o
    .io_output_aw_payload_burst  (writeOnly_io_output_aw_payload_burst[1:0] ), //o
    .io_output_aw_payload_lock   (writeOnly_io_output_aw_payload_lock       ), //o
    .io_output_aw_payload_cache  (writeOnly_io_output_aw_payload_cache[3:0] ), //o
    .io_output_aw_payload_qos    (writeOnly_io_output_aw_payload_qos[3:0]   ), //o
    .io_output_aw_payload_prot   (writeOnly_io_output_aw_payload_prot[2:0]  ), //o
    .io_output_w_valid           (writeOnly_io_output_w_valid               ), //o
    .io_output_w_ready           (io_output_w_ready                         ), //i
    .io_output_w_payload_data    (writeOnly_io_output_w_payload_data[127:0] ), //o
    .io_output_w_payload_strb    (writeOnly_io_output_w_payload_strb[15:0]  ), //o
    .io_output_w_payload_last    (writeOnly_io_output_w_payload_last        ), //o
    .io_output_b_valid           (io_output_b_valid                         ), //i
    .io_output_b_ready           (writeOnly_io_output_b_ready               ), //o
    .io_output_b_payload_id      (io_output_b_payload_id[3:0]               ), //i
    .io_output_b_payload_resp    (io_output_b_payload_resp[1:0]             ), //i
    .io_memoryClk                (io_memoryClk                              ), //i
    .ddrCd_logic_outputReset     (ddrCd_logic_outputReset                   )  //i
  );
  assign io_input_ar_ready = readOnly_io_input_ar_ready;
  assign io_input_r_valid = readOnly_io_input_r_valid;
  assign io_input_r_payload_data = readOnly_io_input_r_payload_data;
  assign io_input_r_payload_id = readOnly_io_input_r_payload_id;
  assign io_input_r_payload_resp = readOnly_io_input_r_payload_resp;
  assign io_input_r_payload_last = readOnly_io_input_r_payload_last;
  assign io_input_aw_ready = writeOnly_io_input_aw_ready;
  assign io_input_w_ready = writeOnly_io_input_w_ready;
  assign io_input_b_valid = writeOnly_io_input_b_valid;
  assign io_input_b_payload_id = writeOnly_io_input_b_payload_id;
  assign io_input_b_payload_resp = writeOnly_io_input_b_payload_resp;
  assign io_output_ar_valid = readOnly_io_output_ar_valid;
  assign io_output_ar_payload_addr = readOnly_io_output_ar_payload_addr;
  assign io_output_ar_payload_id = readOnly_io_output_ar_payload_id;
  assign io_output_ar_payload_region = readOnly_io_output_ar_payload_region;
  assign io_output_ar_payload_len = readOnly_io_output_ar_payload_len;
  assign io_output_ar_payload_size = readOnly_io_output_ar_payload_size;
  assign io_output_ar_payload_burst = readOnly_io_output_ar_payload_burst;
  assign io_output_ar_payload_lock = readOnly_io_output_ar_payload_lock;
  assign io_output_ar_payload_cache = readOnly_io_output_ar_payload_cache;
  assign io_output_ar_payload_qos = readOnly_io_output_ar_payload_qos;
  assign io_output_ar_payload_prot = readOnly_io_output_ar_payload_prot;
  assign io_output_r_ready = readOnly_io_output_r_ready;
  assign io_output_aw_valid = writeOnly_io_output_aw_valid;
  assign io_output_aw_payload_addr = writeOnly_io_output_aw_payload_addr;
  assign io_output_aw_payload_id = writeOnly_io_output_aw_payload_id;
  assign io_output_aw_payload_region = writeOnly_io_output_aw_payload_region;
  assign io_output_aw_payload_len = writeOnly_io_output_aw_payload_len;
  assign io_output_aw_payload_size = writeOnly_io_output_aw_payload_size;
  assign io_output_aw_payload_burst = writeOnly_io_output_aw_payload_burst;
  assign io_output_aw_payload_lock = writeOnly_io_output_aw_payload_lock;
  assign io_output_aw_payload_cache = writeOnly_io_output_aw_payload_cache;
  assign io_output_aw_payload_qos = writeOnly_io_output_aw_payload_qos;
  assign io_output_aw_payload_prot = writeOnly_io_output_aw_payload_prot;
  assign io_output_w_valid = writeOnly_io_output_w_valid;
  assign io_output_w_payload_data = writeOnly_io_output_w_payload_data;
  assign io_output_w_payload_strb = writeOnly_io_output_w_payload_strb;
  assign io_output_w_payload_last = writeOnly_io_output_w_payload_last;
  assign io_output_b_ready = writeOnly_io_output_b_ready;

endmodule

module Axi4CC (
  input  wire          io_input_aw_valid,
  output wire          io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [3:0]    io_input_aw_payload_region,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire [0:0]    io_input_aw_payload_lock,
  input  wire [3:0]    io_input_aw_payload_cache,
  input  wire [3:0]    io_input_aw_payload_qos,
  input  wire [2:0]    io_input_aw_payload_prot,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [31:0]   io_input_w_payload_data,
  input  wire [3:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output wire [3:0]    io_input_b_payload_id,
  output wire [1:0]    io_input_b_payload_resp,
  input  wire          io_input_ar_valid,
  output wire          io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [3:0]    io_input_ar_payload_region,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  input  wire [0:0]    io_input_ar_payload_lock,
  input  wire [3:0]    io_input_ar_payload_cache,
  input  wire [3:0]    io_input_ar_payload_qos,
  input  wire [2:0]    io_input_ar_payload_prot,
  output wire          io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [31:0]   io_input_r_payload_data,
  output wire [3:0]    io_input_r_payload_id,
  output wire [1:0]    io_input_r_payload_resp,
  output wire          io_input_r_payload_last,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [3:0]    io_output_aw_payload_id,
  output wire [3:0]    io_output_aw_payload_region,
  output wire [7:0]    io_output_aw_payload_len,
  output wire [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire [0:0]    io_output_aw_payload_lock,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [3:0]    io_output_aw_payload_qos,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [31:0]   io_output_w_payload_data,
  output wire [3:0]    io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [3:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [3:0]    io_output_ar_payload_id,
  output wire [3:0]    io_output_ar_payload_region,
  output wire [7:0]    io_output_ar_payload_len,
  output wire [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  output wire [0:0]    io_output_ar_payload_lock,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [3:0]    io_output_ar_payload_qos,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [31:0]   io_output_r_payload_data,
  input  wire [3:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_ddrMasters_1_clk,
  input  wire          io_ddrMasters_1_reset,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                io_input_ar_queue_io_push_ready;
  wire                io_input_ar_queue_io_pop_valid;
  wire       [31:0]   io_input_ar_queue_io_pop_payload_addr;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_id;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_region;
  wire       [7:0]    io_input_ar_queue_io_pop_payload_len;
  wire       [2:0]    io_input_ar_queue_io_pop_payload_size;
  wire       [1:0]    io_input_ar_queue_io_pop_payload_burst;
  wire       [0:0]    io_input_ar_queue_io_pop_payload_lock;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_cache;
  wire       [3:0]    io_input_ar_queue_io_pop_payload_qos;
  wire       [2:0]    io_input_ar_queue_io_pop_payload_prot;
  wire       [4:0]    io_input_ar_queue_io_pushOccupancy;
  wire       [4:0]    io_input_ar_queue_io_popOccupancy;
  wire                io_input_ar_queue_system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1;
  wire                io_output_r_queue_io_push_ready;
  wire                io_output_r_queue_io_pop_valid;
  wire       [31:0]   io_output_r_queue_io_pop_payload_data;
  wire       [3:0]    io_output_r_queue_io_pop_payload_id;
  wire       [1:0]    io_output_r_queue_io_pop_payload_resp;
  wire                io_output_r_queue_io_pop_payload_last;
  wire       [4:0]    io_output_r_queue_io_pushOccupancy;
  wire       [4:0]    io_output_r_queue_io_popOccupancy;
  wire                io_output_r_queue_system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1;
  wire                io_input_aw_queue_io_push_ready;
  wire                io_input_aw_queue_io_pop_valid;
  wire       [31:0]   io_input_aw_queue_io_pop_payload_addr;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_id;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_region;
  wire       [7:0]    io_input_aw_queue_io_pop_payload_len;
  wire       [2:0]    io_input_aw_queue_io_pop_payload_size;
  wire       [1:0]    io_input_aw_queue_io_pop_payload_burst;
  wire       [0:0]    io_input_aw_queue_io_pop_payload_lock;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_cache;
  wire       [3:0]    io_input_aw_queue_io_pop_payload_qos;
  wire       [2:0]    io_input_aw_queue_io_pop_payload_prot;
  wire       [4:0]    io_input_aw_queue_io_pushOccupancy;
  wire       [4:0]    io_input_aw_queue_io_popOccupancy;
  wire                io_input_w_queue_io_push_ready;
  wire                io_input_w_queue_io_pop_valid;
  wire       [31:0]   io_input_w_queue_io_pop_payload_data;
  wire       [3:0]    io_input_w_queue_io_pop_payload_strb;
  wire                io_input_w_queue_io_pop_payload_last;
  wire       [4:0]    io_input_w_queue_io_pushOccupancy;
  wire       [4:0]    io_input_w_queue_io_popOccupancy;
  wire                io_output_b_queue_io_push_ready;
  wire                io_output_b_queue_io_pop_valid;
  wire       [3:0]    io_output_b_queue_io_pop_payload_id;
  wire       [1:0]    io_output_b_queue_io_pop_payload_resp;
  wire       [4:0]    io_output_b_queue_io_pushOccupancy;
  wire       [4:0]    io_output_b_queue_io_popOccupancy;

  StreamFifoCC_2 io_input_ar_queue (
    .io_push_valid                                                                           (io_input_ar_valid                                                                                        ), //i
    .io_push_ready                                                                           (io_input_ar_queue_io_push_ready                                                                          ), //o
    .io_push_payload_addr                                                                    (io_input_ar_payload_addr[31:0]                                                                           ), //i
    .io_push_payload_id                                                                      (io_input_ar_payload_id[3:0]                                                                              ), //i
    .io_push_payload_region                                                                  (io_input_ar_payload_region[3:0]                                                                          ), //i
    .io_push_payload_len                                                                     (io_input_ar_payload_len[7:0]                                                                             ), //i
    .io_push_payload_size                                                                    (io_input_ar_payload_size[2:0]                                                                            ), //i
    .io_push_payload_burst                                                                   (io_input_ar_payload_burst[1:0]                                                                           ), //i
    .io_push_payload_lock                                                                    (io_input_ar_payload_lock                                                                                 ), //i
    .io_push_payload_cache                                                                   (io_input_ar_payload_cache[3:0]                                                                           ), //i
    .io_push_payload_qos                                                                     (io_input_ar_payload_qos[3:0]                                                                             ), //i
    .io_push_payload_prot                                                                    (io_input_ar_payload_prot[2:0]                                                                            ), //i
    .io_pop_valid                                                                            (io_input_ar_queue_io_pop_valid                                                                           ), //o
    .io_pop_ready                                                                            (io_output_ar_ready                                                                                       ), //i
    .io_pop_payload_addr                                                                     (io_input_ar_queue_io_pop_payload_addr[31:0]                                                              ), //o
    .io_pop_payload_id                                                                       (io_input_ar_queue_io_pop_payload_id[3:0]                                                                 ), //o
    .io_pop_payload_region                                                                   (io_input_ar_queue_io_pop_payload_region[3:0]                                                             ), //o
    .io_pop_payload_len                                                                      (io_input_ar_queue_io_pop_payload_len[7:0]                                                                ), //o
    .io_pop_payload_size                                                                     (io_input_ar_queue_io_pop_payload_size[2:0]                                                               ), //o
    .io_pop_payload_burst                                                                    (io_input_ar_queue_io_pop_payload_burst[1:0]                                                              ), //o
    .io_pop_payload_lock                                                                     (io_input_ar_queue_io_pop_payload_lock                                                                    ), //o
    .io_pop_payload_cache                                                                    (io_input_ar_queue_io_pop_payload_cache[3:0]                                                              ), //o
    .io_pop_payload_qos                                                                      (io_input_ar_queue_io_pop_payload_qos[3:0]                                                                ), //o
    .io_pop_payload_prot                                                                     (io_input_ar_queue_io_pop_payload_prot[2:0]                                                               ), //o
    .io_pushOccupancy                                                                        (io_input_ar_queue_io_pushOccupancy[4:0]                                                                  ), //o
    .io_popOccupancy                                                                         (io_input_ar_queue_io_popOccupancy[4:0]                                                                   ), //o
    .io_ddrMasters_1_clk                                                                     (io_ddrMasters_1_clk                                                                                      ), //i
    .io_ddrMasters_1_reset                                                                   (io_ddrMasters_1_reset                                                                                    ), //i
    .io_memoryClk                                                                            (io_memoryClk                                                                                             ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1 (io_input_ar_queue_system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1)  //o
  );
  StreamFifoCC_3 io_output_r_queue (
    .io_push_valid                                                                             (io_output_r_valid                                                                                          ), //i
    .io_push_ready                                                                             (io_output_r_queue_io_push_ready                                                                            ), //o
    .io_push_payload_data                                                                      (io_output_r_payload_data[31:0]                                                                             ), //i
    .io_push_payload_id                                                                        (io_output_r_payload_id[3:0]                                                                                ), //i
    .io_push_payload_resp                                                                      (io_output_r_payload_resp[1:0]                                                                              ), //i
    .io_push_payload_last                                                                      (io_output_r_payload_last                                                                                   ), //i
    .io_pop_valid                                                                              (io_output_r_queue_io_pop_valid                                                                             ), //o
    .io_pop_ready                                                                              (io_input_r_ready                                                                                           ), //i
    .io_pop_payload_data                                                                       (io_output_r_queue_io_pop_payload_data[31:0]                                                                ), //o
    .io_pop_payload_id                                                                         (io_output_r_queue_io_pop_payload_id[3:0]                                                                   ), //o
    .io_pop_payload_resp                                                                       (io_output_r_queue_io_pop_payload_resp[1:0]                                                                 ), //o
    .io_pop_payload_last                                                                       (io_output_r_queue_io_pop_payload_last                                                                      ), //o
    .io_pushOccupancy                                                                          (io_output_r_queue_io_pushOccupancy[4:0]                                                                    ), //o
    .io_popOccupancy                                                                           (io_output_r_queue_io_popOccupancy[4:0]                                                                     ), //o
    .io_memoryClk                                                                              (io_memoryClk                                                                                               ), //i
    .ddrCd_logic_outputReset                                                                   (ddrCd_logic_outputReset                                                                                    ), //i
    .io_ddrMasters_1_clk                                                                       (io_ddrMasters_1_clk                                                                                        ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 (io_output_r_queue_system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1)  //o
  );
  StreamFifoCC_4 io_input_aw_queue (
    .io_push_valid                                                                           (io_input_aw_valid                                                                                        ), //i
    .io_push_ready                                                                           (io_input_aw_queue_io_push_ready                                                                          ), //o
    .io_push_payload_addr                                                                    (io_input_aw_payload_addr[31:0]                                                                           ), //i
    .io_push_payload_id                                                                      (io_input_aw_payload_id[3:0]                                                                              ), //i
    .io_push_payload_region                                                                  (io_input_aw_payload_region[3:0]                                                                          ), //i
    .io_push_payload_len                                                                     (io_input_aw_payload_len[7:0]                                                                             ), //i
    .io_push_payload_size                                                                    (io_input_aw_payload_size[2:0]                                                                            ), //i
    .io_push_payload_burst                                                                   (io_input_aw_payload_burst[1:0]                                                                           ), //i
    .io_push_payload_lock                                                                    (io_input_aw_payload_lock                                                                                 ), //i
    .io_push_payload_cache                                                                   (io_input_aw_payload_cache[3:0]                                                                           ), //i
    .io_push_payload_qos                                                                     (io_input_aw_payload_qos[3:0]                                                                             ), //i
    .io_push_payload_prot                                                                    (io_input_aw_payload_prot[2:0]                                                                            ), //i
    .io_pop_valid                                                                            (io_input_aw_queue_io_pop_valid                                                                           ), //o
    .io_pop_ready                                                                            (io_output_aw_ready                                                                                       ), //i
    .io_pop_payload_addr                                                                     (io_input_aw_queue_io_pop_payload_addr[31:0]                                                              ), //o
    .io_pop_payload_id                                                                       (io_input_aw_queue_io_pop_payload_id[3:0]                                                                 ), //o
    .io_pop_payload_region                                                                   (io_input_aw_queue_io_pop_payload_region[3:0]                                                             ), //o
    .io_pop_payload_len                                                                      (io_input_aw_queue_io_pop_payload_len[7:0]                                                                ), //o
    .io_pop_payload_size                                                                     (io_input_aw_queue_io_pop_payload_size[2:0]                                                               ), //o
    .io_pop_payload_burst                                                                    (io_input_aw_queue_io_pop_payload_burst[1:0]                                                              ), //o
    .io_pop_payload_lock                                                                     (io_input_aw_queue_io_pop_payload_lock                                                                    ), //o
    .io_pop_payload_cache                                                                    (io_input_aw_queue_io_pop_payload_cache[3:0]                                                              ), //o
    .io_pop_payload_qos                                                                      (io_input_aw_queue_io_pop_payload_qos[3:0]                                                                ), //o
    .io_pop_payload_prot                                                                     (io_input_aw_queue_io_pop_payload_prot[2:0]                                                               ), //o
    .io_pushOccupancy                                                                        (io_input_aw_queue_io_pushOccupancy[4:0]                                                                  ), //o
    .io_popOccupancy                                                                         (io_input_aw_queue_io_popOccupancy[4:0]                                                                   ), //o
    .io_ddrMasters_1_clk                                                                     (io_ddrMasters_1_clk                                                                                      ), //i
    .io_ddrMasters_1_reset                                                                   (io_ddrMasters_1_reset                                                                                    ), //i
    .io_memoryClk                                                                            (io_memoryClk                                                                                             ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1 (io_input_ar_queue_system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1)  //i
  );
  StreamFifoCC_5 io_input_w_queue (
    .io_push_valid                                                                           (io_input_w_valid                                                                                         ), //i
    .io_push_ready                                                                           (io_input_w_queue_io_push_ready                                                                           ), //o
    .io_push_payload_data                                                                    (io_input_w_payload_data[31:0]                                                                            ), //i
    .io_push_payload_strb                                                                    (io_input_w_payload_strb[3:0]                                                                             ), //i
    .io_push_payload_last                                                                    (io_input_w_payload_last                                                                                  ), //i
    .io_pop_valid                                                                            (io_input_w_queue_io_pop_valid                                                                            ), //o
    .io_pop_ready                                                                            (io_output_w_ready                                                                                        ), //i
    .io_pop_payload_data                                                                     (io_input_w_queue_io_pop_payload_data[31:0]                                                               ), //o
    .io_pop_payload_strb                                                                     (io_input_w_queue_io_pop_payload_strb[3:0]                                                                ), //o
    .io_pop_payload_last                                                                     (io_input_w_queue_io_pop_payload_last                                                                     ), //o
    .io_pushOccupancy                                                                        (io_input_w_queue_io_pushOccupancy[4:0]                                                                   ), //o
    .io_popOccupancy                                                                         (io_input_w_queue_io_popOccupancy[4:0]                                                                    ), //o
    .io_ddrMasters_1_clk                                                                     (io_ddrMasters_1_clk                                                                                      ), //i
    .io_ddrMasters_1_reset                                                                   (io_ddrMasters_1_reset                                                                                    ), //i
    .io_memoryClk                                                                            (io_memoryClk                                                                                             ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1 (io_input_ar_queue_system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1)  //i
  );
  StreamFifoCC_6 io_output_b_queue (
    .io_push_valid                                                                             (io_output_b_valid                                                                                          ), //i
    .io_push_ready                                                                             (io_output_b_queue_io_push_ready                                                                            ), //o
    .io_push_payload_id                                                                        (io_output_b_payload_id[3:0]                                                                                ), //i
    .io_push_payload_resp                                                                      (io_output_b_payload_resp[1:0]                                                                              ), //i
    .io_pop_valid                                                                              (io_output_b_queue_io_pop_valid                                                                             ), //o
    .io_pop_ready                                                                              (io_input_b_ready                                                                                           ), //i
    .io_pop_payload_id                                                                         (io_output_b_queue_io_pop_payload_id[3:0]                                                                   ), //o
    .io_pop_payload_resp                                                                       (io_output_b_queue_io_pop_payload_resp[1:0]                                                                 ), //o
    .io_pushOccupancy                                                                          (io_output_b_queue_io_pushOccupancy[4:0]                                                                    ), //o
    .io_popOccupancy                                                                           (io_output_b_queue_io_popOccupancy[4:0]                                                                     ), //o
    .io_memoryClk                                                                              (io_memoryClk                                                                                               ), //i
    .ddrCd_logic_outputReset                                                                   (ddrCd_logic_outputReset                                                                                    ), //i
    .io_ddrMasters_1_clk                                                                       (io_ddrMasters_1_clk                                                                                        ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 (io_output_r_queue_system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1)  //i
  );
  assign io_input_ar_ready = io_input_ar_queue_io_push_ready;
  assign io_output_ar_valid = io_input_ar_queue_io_pop_valid;
  assign io_output_ar_payload_addr = io_input_ar_queue_io_pop_payload_addr;
  assign io_output_ar_payload_id = io_input_ar_queue_io_pop_payload_id;
  assign io_output_ar_payload_region = io_input_ar_queue_io_pop_payload_region;
  assign io_output_ar_payload_len = io_input_ar_queue_io_pop_payload_len;
  assign io_output_ar_payload_size = io_input_ar_queue_io_pop_payload_size;
  assign io_output_ar_payload_burst = io_input_ar_queue_io_pop_payload_burst;
  assign io_output_ar_payload_lock = io_input_ar_queue_io_pop_payload_lock;
  assign io_output_ar_payload_cache = io_input_ar_queue_io_pop_payload_cache;
  assign io_output_ar_payload_qos = io_input_ar_queue_io_pop_payload_qos;
  assign io_output_ar_payload_prot = io_input_ar_queue_io_pop_payload_prot;
  assign io_output_r_ready = io_output_r_queue_io_push_ready;
  assign io_input_r_valid = io_output_r_queue_io_pop_valid;
  assign io_input_r_payload_data = io_output_r_queue_io_pop_payload_data;
  assign io_input_r_payload_id = io_output_r_queue_io_pop_payload_id;
  assign io_input_r_payload_resp = io_output_r_queue_io_pop_payload_resp;
  assign io_input_r_payload_last = io_output_r_queue_io_pop_payload_last;
  assign io_input_aw_ready = io_input_aw_queue_io_push_ready;
  assign io_output_aw_valid = io_input_aw_queue_io_pop_valid;
  assign io_output_aw_payload_addr = io_input_aw_queue_io_pop_payload_addr;
  assign io_output_aw_payload_id = io_input_aw_queue_io_pop_payload_id;
  assign io_output_aw_payload_region = io_input_aw_queue_io_pop_payload_region;
  assign io_output_aw_payload_len = io_input_aw_queue_io_pop_payload_len;
  assign io_output_aw_payload_size = io_input_aw_queue_io_pop_payload_size;
  assign io_output_aw_payload_burst = io_input_aw_queue_io_pop_payload_burst;
  assign io_output_aw_payload_lock = io_input_aw_queue_io_pop_payload_lock;
  assign io_output_aw_payload_cache = io_input_aw_queue_io_pop_payload_cache;
  assign io_output_aw_payload_qos = io_input_aw_queue_io_pop_payload_qos;
  assign io_output_aw_payload_prot = io_input_aw_queue_io_pop_payload_prot;
  assign io_input_w_ready = io_input_w_queue_io_push_ready;
  assign io_output_w_valid = io_input_w_queue_io_pop_valid;
  assign io_output_w_payload_data = io_input_w_queue_io_pop_payload_data;
  assign io_output_w_payload_strb = io_input_w_queue_io_pop_payload_strb;
  assign io_output_w_payload_last = io_input_w_queue_io_pop_payload_last;
  assign io_output_b_ready = io_output_b_queue_io_push_ready;
  assign io_input_b_valid = io_output_b_queue_io_pop_valid;
  assign io_input_b_payload_id = io_output_b_queue_io_pop_payload_id;
  assign io_input_b_payload_resp = io_output_b_queue_io_pop_payload_resp;

endmodule

module BufferCC_66 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_ddrMasters_1_clk,
  input  wire          io_ddrMasters_1_reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_1_clk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

module Axi4WriteOnlyArbiter (
  input  wire          io_inputs_0_aw_valid,
  output wire          io_inputs_0_aw_ready,
  input  wire [31:0]   io_inputs_0_aw_payload_addr,
  input  wire [5:0]    io_inputs_0_aw_payload_id,
  input  wire [3:0]    io_inputs_0_aw_payload_region,
  input  wire [7:0]    io_inputs_0_aw_payload_len,
  input  wire [2:0]    io_inputs_0_aw_payload_size,
  input  wire [1:0]    io_inputs_0_aw_payload_burst,
  input  wire [0:0]    io_inputs_0_aw_payload_lock,
  input  wire [3:0]    io_inputs_0_aw_payload_cache,
  input  wire [3:0]    io_inputs_0_aw_payload_qos,
  input  wire [2:0]    io_inputs_0_aw_payload_prot,
  input  wire          io_inputs_0_w_valid,
  output wire          io_inputs_0_w_ready,
  input  wire [127:0]  io_inputs_0_w_payload_data,
  input  wire [15:0]   io_inputs_0_w_payload_strb,
  input  wire          io_inputs_0_w_payload_last,
  output wire          io_inputs_0_b_valid,
  input  wire          io_inputs_0_b_ready,
  output wire [5:0]    io_inputs_0_b_payload_id,
  output wire [1:0]    io_inputs_0_b_payload_resp,
  input  wire          io_inputs_1_aw_valid,
  output wire          io_inputs_1_aw_ready,
  input  wire [31:0]   io_inputs_1_aw_payload_addr,
  input  wire [5:0]    io_inputs_1_aw_payload_id,
  input  wire [3:0]    io_inputs_1_aw_payload_region,
  input  wire [7:0]    io_inputs_1_aw_payload_len,
  input  wire [2:0]    io_inputs_1_aw_payload_size,
  input  wire [1:0]    io_inputs_1_aw_payload_burst,
  input  wire [0:0]    io_inputs_1_aw_payload_lock,
  input  wire [3:0]    io_inputs_1_aw_payload_cache,
  input  wire [3:0]    io_inputs_1_aw_payload_qos,
  input  wire [2:0]    io_inputs_1_aw_payload_prot,
  input  wire          io_inputs_1_w_valid,
  output wire          io_inputs_1_w_ready,
  input  wire [127:0]  io_inputs_1_w_payload_data,
  input  wire [15:0]   io_inputs_1_w_payload_strb,
  input  wire          io_inputs_1_w_payload_last,
  output wire          io_inputs_1_b_valid,
  input  wire          io_inputs_1_b_ready,
  output wire [5:0]    io_inputs_1_b_payload_id,
  output wire [1:0]    io_inputs_1_b_payload_resp,
  input  wire          io_inputs_2_aw_valid,
  output wire          io_inputs_2_aw_ready,
  input  wire [31:0]   io_inputs_2_aw_payload_addr,
  input  wire [5:0]    io_inputs_2_aw_payload_id,
  input  wire [3:0]    io_inputs_2_aw_payload_region,
  input  wire [7:0]    io_inputs_2_aw_payload_len,
  input  wire [2:0]    io_inputs_2_aw_payload_size,
  input  wire [1:0]    io_inputs_2_aw_payload_burst,
  input  wire [0:0]    io_inputs_2_aw_payload_lock,
  input  wire [3:0]    io_inputs_2_aw_payload_cache,
  input  wire [3:0]    io_inputs_2_aw_payload_qos,
  input  wire [2:0]    io_inputs_2_aw_payload_prot,
  input  wire          io_inputs_2_w_valid,
  output wire          io_inputs_2_w_ready,
  input  wire [127:0]  io_inputs_2_w_payload_data,
  input  wire [15:0]   io_inputs_2_w_payload_strb,
  input  wire          io_inputs_2_w_payload_last,
  output wire          io_inputs_2_b_valid,
  input  wire          io_inputs_2_b_ready,
  output wire [5:0]    io_inputs_2_b_payload_id,
  output wire [1:0]    io_inputs_2_b_payload_resp,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [7:0]    io_output_aw_payload_id,
  output wire [3:0]    io_output_aw_payload_region,
  output wire [7:0]    io_output_aw_payload_len,
  output wire [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire [0:0]    io_output_aw_payload_lock,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [3:0]    io_output_aw_payload_qos,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [127:0]  io_output_w_payload_data,
  output wire [15:0]   io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [7:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  reg                 cmdArbiter_io_output_ready;
  reg                 cmdRouteFork_translated_fifo_io_pop_ready;
  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_inputs_2_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [31:0]   cmdArbiter_io_output_payload_addr;
  wire       [5:0]    cmdArbiter_io_output_payload_id;
  wire       [3:0]    cmdArbiter_io_output_payload_region;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire       [0:0]    cmdArbiter_io_output_payload_lock;
  wire       [3:0]    cmdArbiter_io_output_payload_cache;
  wire       [3:0]    cmdArbiter_io_output_payload_qos;
  wire       [2:0]    cmdArbiter_io_output_payload_prot;
  wire       [1:0]    cmdArbiter_io_chosen;
  wire       [2:0]    cmdArbiter_io_chosenOH;
  wire                cmdRouteFork_translated_fifo_io_push_ready;
  wire                cmdRouteFork_translated_fifo_io_pop_valid;
  wire       [1:0]    cmdRouteFork_translated_fifo_io_pop_payload;
  wire       [2:0]    cmdRouteFork_translated_fifo_io_occupancy;
  wire       [2:0]    cmdRouteFork_translated_fifo_io_availability;
  reg                 _zz_io_output_w_valid;
  reg        [127:0]  _zz_io_output_w_payload_data;
  reg        [15:0]   _zz_io_output_w_payload_strb;
  reg                 _zz_io_output_w_payload_last;
  reg                 _zz_io_output_b_ready;
  wire                cmdOutputFork_valid;
  wire                cmdOutputFork_ready;
  wire       [31:0]   cmdOutputFork_payload_addr;
  wire       [5:0]    cmdOutputFork_payload_id;
  wire       [3:0]    cmdOutputFork_payload_region;
  wire       [7:0]    cmdOutputFork_payload_len;
  wire       [2:0]    cmdOutputFork_payload_size;
  wire       [1:0]    cmdOutputFork_payload_burst;
  wire       [0:0]    cmdOutputFork_payload_lock;
  wire       [3:0]    cmdOutputFork_payload_cache;
  wire       [3:0]    cmdOutputFork_payload_qos;
  wire       [2:0]    cmdOutputFork_payload_prot;
  wire                cmdRouteFork_valid;
  wire                cmdRouteFork_ready;
  wire       [31:0]   cmdRouteFork_payload_addr;
  wire       [5:0]    cmdRouteFork_payload_id;
  wire       [3:0]    cmdRouteFork_payload_region;
  wire       [7:0]    cmdRouteFork_payload_len;
  wire       [2:0]    cmdRouteFork_payload_size;
  wire       [1:0]    cmdRouteFork_payload_burst;
  wire       [0:0]    cmdRouteFork_payload_lock;
  wire       [3:0]    cmdRouteFork_payload_cache;
  wire       [3:0]    cmdRouteFork_payload_qos;
  wire       [2:0]    cmdRouteFork_payload_prot;
  reg                 cmdArbiter_io_output_fork2_logic_linkEnable_0;
  reg                 cmdArbiter_io_output_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdOutputFork_fire;
  wire                cmdRouteFork_fire;
  wire                cmdRouteFork_translated_valid;
  wire                cmdRouteFork_translated_ready;
  wire       [1:0]    cmdRouteFork_translated_payload;
  wire                cmdRouteFork_translated_fifo_io_pop_m2sPipe_valid;
  wire                cmdRouteFork_translated_fifo_io_pop_m2sPipe_ready;
  wire       [1:0]    cmdRouteFork_translated_fifo_io_pop_m2sPipe_payload;
  reg                 cmdRouteFork_translated_fifo_io_pop_rValid;
  reg        [1:0]    cmdRouteFork_translated_fifo_io_pop_rData;
  wire                when_Stream_l375;
  wire                cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_valid;
  wire                cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_ready;
  wire       [1:0]    cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_payload;
  reg                 cmdRouteFork_translated_fifo_io_pop_m2sPipe_rValidN;
  reg        [1:0]    cmdRouteFork_translated_fifo_io_pop_m2sPipe_rData;
  wire                io_output_w_fire;
  wire       [1:0]    writeRspIndex;
  wire                writeRspSels_0;
  wire                writeRspSels_1;
  wire                writeRspSels_2;

  StreamArbiter_7 cmdArbiter (
    .io_inputs_0_valid          (io_inputs_0_aw_valid                    ), //i
    .io_inputs_0_ready          (cmdArbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_addr   (io_inputs_0_aw_payload_addr[31:0]       ), //i
    .io_inputs_0_payload_id     (io_inputs_0_aw_payload_id[5:0]          ), //i
    .io_inputs_0_payload_region (io_inputs_0_aw_payload_region[3:0]      ), //i
    .io_inputs_0_payload_len    (io_inputs_0_aw_payload_len[7:0]         ), //i
    .io_inputs_0_payload_size   (io_inputs_0_aw_payload_size[2:0]        ), //i
    .io_inputs_0_payload_burst  (io_inputs_0_aw_payload_burst[1:0]       ), //i
    .io_inputs_0_payload_lock   (io_inputs_0_aw_payload_lock             ), //i
    .io_inputs_0_payload_cache  (io_inputs_0_aw_payload_cache[3:0]       ), //i
    .io_inputs_0_payload_qos    (io_inputs_0_aw_payload_qos[3:0]         ), //i
    .io_inputs_0_payload_prot   (io_inputs_0_aw_payload_prot[2:0]        ), //i
    .io_inputs_1_valid          (io_inputs_1_aw_valid                    ), //i
    .io_inputs_1_ready          (cmdArbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_addr   (io_inputs_1_aw_payload_addr[31:0]       ), //i
    .io_inputs_1_payload_id     (io_inputs_1_aw_payload_id[5:0]          ), //i
    .io_inputs_1_payload_region (io_inputs_1_aw_payload_region[3:0]      ), //i
    .io_inputs_1_payload_len    (io_inputs_1_aw_payload_len[7:0]         ), //i
    .io_inputs_1_payload_size   (io_inputs_1_aw_payload_size[2:0]        ), //i
    .io_inputs_1_payload_burst  (io_inputs_1_aw_payload_burst[1:0]       ), //i
    .io_inputs_1_payload_lock   (io_inputs_1_aw_payload_lock             ), //i
    .io_inputs_1_payload_cache  (io_inputs_1_aw_payload_cache[3:0]       ), //i
    .io_inputs_1_payload_qos    (io_inputs_1_aw_payload_qos[3:0]         ), //i
    .io_inputs_1_payload_prot   (io_inputs_1_aw_payload_prot[2:0]        ), //i
    .io_inputs_2_valid          (io_inputs_2_aw_valid                    ), //i
    .io_inputs_2_ready          (cmdArbiter_io_inputs_2_ready            ), //o
    .io_inputs_2_payload_addr   (io_inputs_2_aw_payload_addr[31:0]       ), //i
    .io_inputs_2_payload_id     (io_inputs_2_aw_payload_id[5:0]          ), //i
    .io_inputs_2_payload_region (io_inputs_2_aw_payload_region[3:0]      ), //i
    .io_inputs_2_payload_len    (io_inputs_2_aw_payload_len[7:0]         ), //i
    .io_inputs_2_payload_size   (io_inputs_2_aw_payload_size[2:0]        ), //i
    .io_inputs_2_payload_burst  (io_inputs_2_aw_payload_burst[1:0]       ), //i
    .io_inputs_2_payload_lock   (io_inputs_2_aw_payload_lock             ), //i
    .io_inputs_2_payload_cache  (io_inputs_2_aw_payload_cache[3:0]       ), //i
    .io_inputs_2_payload_qos    (io_inputs_2_aw_payload_qos[3:0]         ), //i
    .io_inputs_2_payload_prot   (io_inputs_2_aw_payload_prot[2:0]        ), //i
    .io_output_valid            (cmdArbiter_io_output_valid              ), //o
    .io_output_ready            (cmdArbiter_io_output_ready              ), //i
    .io_output_payload_addr     (cmdArbiter_io_output_payload_addr[31:0] ), //o
    .io_output_payload_id       (cmdArbiter_io_output_payload_id[5:0]    ), //o
    .io_output_payload_region   (cmdArbiter_io_output_payload_region[3:0]), //o
    .io_output_payload_len      (cmdArbiter_io_output_payload_len[7:0]   ), //o
    .io_output_payload_size     (cmdArbiter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_burst    (cmdArbiter_io_output_payload_burst[1:0] ), //o
    .io_output_payload_lock     (cmdArbiter_io_output_payload_lock       ), //o
    .io_output_payload_cache    (cmdArbiter_io_output_payload_cache[3:0] ), //o
    .io_output_payload_qos      (cmdArbiter_io_output_payload_qos[3:0]   ), //o
    .io_output_payload_prot     (cmdArbiter_io_output_payload_prot[2:0]  ), //o
    .io_chosen                  (cmdArbiter_io_chosen[1:0]               ), //o
    .io_chosenOH                (cmdArbiter_io_chosenOH[2:0]             ), //o
    .io_memoryClk               (io_memoryClk                            ), //i
    .ddrCd_logic_outputReset    (ddrCd_logic_outputReset                 )  //i
  );
  StreamFifoLowLatency cmdRouteFork_translated_fifo (
    .io_push_valid           (cmdRouteFork_translated_valid                    ), //i
    .io_push_ready           (cmdRouteFork_translated_fifo_io_push_ready       ), //o
    .io_push_payload         (cmdRouteFork_translated_payload[1:0]             ), //i
    .io_pop_valid            (cmdRouteFork_translated_fifo_io_pop_valid        ), //o
    .io_pop_ready            (cmdRouteFork_translated_fifo_io_pop_ready        ), //i
    .io_pop_payload          (cmdRouteFork_translated_fifo_io_pop_payload[1:0] ), //o
    .io_flush                (1'b0                                             ), //i
    .io_occupancy            (cmdRouteFork_translated_fifo_io_occupancy[2:0]   ), //o
    .io_availability         (cmdRouteFork_translated_fifo_io_availability[2:0]), //o
    .io_memoryClk            (io_memoryClk                                     ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                          )  //i
  );
  always @(*) begin
    case(cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_payload)
      2'b00 : begin
        _zz_io_output_w_valid = io_inputs_0_w_valid;
        _zz_io_output_w_payload_data = io_inputs_0_w_payload_data;
        _zz_io_output_w_payload_strb = io_inputs_0_w_payload_strb;
        _zz_io_output_w_payload_last = io_inputs_0_w_payload_last;
      end
      2'b01 : begin
        _zz_io_output_w_valid = io_inputs_1_w_valid;
        _zz_io_output_w_payload_data = io_inputs_1_w_payload_data;
        _zz_io_output_w_payload_strb = io_inputs_1_w_payload_strb;
        _zz_io_output_w_payload_last = io_inputs_1_w_payload_last;
      end
      default : begin
        _zz_io_output_w_valid = io_inputs_2_w_valid;
        _zz_io_output_w_payload_data = io_inputs_2_w_payload_data;
        _zz_io_output_w_payload_strb = io_inputs_2_w_payload_strb;
        _zz_io_output_w_payload_last = io_inputs_2_w_payload_last;
      end
    endcase
  end

  always @(*) begin
    case(writeRspIndex)
      2'b00 : _zz_io_output_b_ready = io_inputs_0_b_ready;
      2'b01 : _zz_io_output_b_ready = io_inputs_1_b_ready;
      default : _zz_io_output_b_ready = io_inputs_2_b_ready;
    endcase
  end

  assign io_inputs_0_aw_ready = cmdArbiter_io_inputs_0_ready;
  assign io_inputs_1_aw_ready = cmdArbiter_io_inputs_1_ready;
  assign io_inputs_2_aw_ready = cmdArbiter_io_inputs_2_ready;
  always @(*) begin
    cmdArbiter_io_output_ready = 1'b1;
    if(when_Stream_l1063) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdOutputFork_ready) && cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdRouteFork_ready) && cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdOutputFork_valid = (cmdArbiter_io_output_valid && cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign cmdOutputFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdOutputFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdOutputFork_payload_region = cmdArbiter_io_output_payload_region;
  assign cmdOutputFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdOutputFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdOutputFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdOutputFork_payload_lock = cmdArbiter_io_output_payload_lock;
  assign cmdOutputFork_payload_cache = cmdArbiter_io_output_payload_cache;
  assign cmdOutputFork_payload_qos = cmdArbiter_io_output_payload_qos;
  assign cmdOutputFork_payload_prot = cmdArbiter_io_output_payload_prot;
  assign cmdOutputFork_fire = (cmdOutputFork_valid && cmdOutputFork_ready);
  assign cmdRouteFork_valid = (cmdArbiter_io_output_valid && cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdRouteFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdRouteFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdRouteFork_payload_region = cmdArbiter_io_output_payload_region;
  assign cmdRouteFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdRouteFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdRouteFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdRouteFork_payload_lock = cmdArbiter_io_output_payload_lock;
  assign cmdRouteFork_payload_cache = cmdArbiter_io_output_payload_cache;
  assign cmdRouteFork_payload_qos = cmdArbiter_io_output_payload_qos;
  assign cmdRouteFork_payload_prot = cmdArbiter_io_output_payload_prot;
  assign cmdRouteFork_fire = (cmdRouteFork_valid && cmdRouteFork_ready);
  assign io_output_aw_valid = cmdOutputFork_valid;
  assign cmdOutputFork_ready = io_output_aw_ready;
  assign io_output_aw_payload_addr = cmdOutputFork_payload_addr;
  assign io_output_aw_payload_region = cmdOutputFork_payload_region;
  assign io_output_aw_payload_len = cmdOutputFork_payload_len;
  assign io_output_aw_payload_size = cmdOutputFork_payload_size;
  assign io_output_aw_payload_burst = cmdOutputFork_payload_burst;
  assign io_output_aw_payload_lock = cmdOutputFork_payload_lock;
  assign io_output_aw_payload_cache = cmdOutputFork_payload_cache;
  assign io_output_aw_payload_qos = cmdOutputFork_payload_qos;
  assign io_output_aw_payload_prot = cmdOutputFork_payload_prot;
  assign io_output_aw_payload_id = {cmdArbiter_io_chosen,cmdArbiter_io_output_payload_id};
  assign cmdRouteFork_translated_valid = cmdRouteFork_valid;
  assign cmdRouteFork_ready = cmdRouteFork_translated_ready;
  assign cmdRouteFork_translated_payload = cmdArbiter_io_chosen;
  assign cmdRouteFork_translated_ready = cmdRouteFork_translated_fifo_io_push_ready;
  always @(*) begin
    cmdRouteFork_translated_fifo_io_pop_ready = cmdRouteFork_translated_fifo_io_pop_m2sPipe_ready;
    if(when_Stream_l375) begin
      cmdRouteFork_translated_fifo_io_pop_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! cmdRouteFork_translated_fifo_io_pop_m2sPipe_valid);
  assign cmdRouteFork_translated_fifo_io_pop_m2sPipe_valid = cmdRouteFork_translated_fifo_io_pop_rValid;
  assign cmdRouteFork_translated_fifo_io_pop_m2sPipe_payload = cmdRouteFork_translated_fifo_io_pop_rData;
  assign cmdRouteFork_translated_fifo_io_pop_m2sPipe_ready = cmdRouteFork_translated_fifo_io_pop_m2sPipe_rValidN;
  assign cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_valid = (cmdRouteFork_translated_fifo_io_pop_m2sPipe_valid || (! cmdRouteFork_translated_fifo_io_pop_m2sPipe_rValidN));
  assign cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_payload = (cmdRouteFork_translated_fifo_io_pop_m2sPipe_rValidN ? cmdRouteFork_translated_fifo_io_pop_m2sPipe_payload : cmdRouteFork_translated_fifo_io_pop_m2sPipe_rData);
  assign io_output_w_valid = (cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_valid && _zz_io_output_w_valid);
  assign io_output_w_payload_data = _zz_io_output_w_payload_data;
  assign io_output_w_payload_strb = _zz_io_output_w_payload_strb;
  assign io_output_w_payload_last = _zz_io_output_w_payload_last;
  assign io_inputs_0_w_ready = ((cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_valid && io_output_w_ready) && (cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_payload == 2'b00));
  assign io_inputs_1_w_ready = ((cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_valid && io_output_w_ready) && (cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_payload == 2'b01));
  assign io_inputs_2_w_ready = ((cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_valid && io_output_w_ready) && (cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_payload == 2'b10));
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_ready = (io_output_w_fire && io_output_w_payload_last);
  assign writeRspIndex = io_output_b_payload_id[7 : 6];
  assign writeRspSels_0 = (writeRspIndex == 2'b00);
  assign writeRspSels_1 = (writeRspIndex == 2'b01);
  assign writeRspSels_2 = (writeRspIndex == 2'b10);
  assign io_inputs_0_b_valid = (io_output_b_valid && writeRspSels_0);
  assign io_inputs_0_b_payload_resp = io_output_b_payload_resp;
  assign io_inputs_0_b_payload_id = io_output_b_payload_id[5 : 0];
  assign io_inputs_1_b_valid = (io_output_b_valid && writeRspSels_1);
  assign io_inputs_1_b_payload_resp = io_output_b_payload_resp;
  assign io_inputs_1_b_payload_id = io_output_b_payload_id[5 : 0];
  assign io_inputs_2_b_valid = (io_output_b_valid && writeRspSels_2);
  assign io_inputs_2_b_payload_resp = io_output_b_payload_resp;
  assign io_inputs_2_b_payload_id = io_output_b_payload_id[5 : 0];
  assign io_output_b_ready = _zz_io_output_b_ready;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
      cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
      cmdRouteFork_translated_fifo_io_pop_rValid <= 1'b0;
      cmdRouteFork_translated_fifo_io_pop_m2sPipe_rValidN <= 1'b1;
    end else begin
      if(cmdOutputFork_fire) begin
        cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdRouteFork_fire) begin
        cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(cmdArbiter_io_output_ready) begin
        cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
        cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(cmdRouteFork_translated_fifo_io_pop_ready) begin
        cmdRouteFork_translated_fifo_io_pop_rValid <= cmdRouteFork_translated_fifo_io_pop_valid;
      end
      if(cmdRouteFork_translated_fifo_io_pop_m2sPipe_valid) begin
        cmdRouteFork_translated_fifo_io_pop_m2sPipe_rValidN <= 1'b0;
      end
      if(cmdRouteFork_translated_fifo_io_pop_m2sPipe_s2mPipe_ready) begin
        cmdRouteFork_translated_fifo_io_pop_m2sPipe_rValidN <= 1'b1;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(cmdRouteFork_translated_fifo_io_pop_ready) begin
      cmdRouteFork_translated_fifo_io_pop_rData <= cmdRouteFork_translated_fifo_io_pop_payload;
    end
    if(cmdRouteFork_translated_fifo_io_pop_m2sPipe_ready) begin
      cmdRouteFork_translated_fifo_io_pop_m2sPipe_rData <= cmdRouteFork_translated_fifo_io_pop_m2sPipe_payload;
    end
  end


endmodule

module Axi4ReadOnlyArbiter (
  input  wire          io_inputs_0_ar_valid,
  output wire          io_inputs_0_ar_ready,
  input  wire [31:0]   io_inputs_0_ar_payload_addr,
  input  wire [5:0]    io_inputs_0_ar_payload_id,
  input  wire [3:0]    io_inputs_0_ar_payload_region,
  input  wire [7:0]    io_inputs_0_ar_payload_len,
  input  wire [2:0]    io_inputs_0_ar_payload_size,
  input  wire [1:0]    io_inputs_0_ar_payload_burst,
  input  wire [0:0]    io_inputs_0_ar_payload_lock,
  input  wire [3:0]    io_inputs_0_ar_payload_cache,
  input  wire [3:0]    io_inputs_0_ar_payload_qos,
  input  wire [2:0]    io_inputs_0_ar_payload_prot,
  output wire          io_inputs_0_r_valid,
  input  wire          io_inputs_0_r_ready,
  output wire [127:0]  io_inputs_0_r_payload_data,
  output wire [5:0]    io_inputs_0_r_payload_id,
  output wire [1:0]    io_inputs_0_r_payload_resp,
  output wire          io_inputs_0_r_payload_last,
  input  wire          io_inputs_1_ar_valid,
  output wire          io_inputs_1_ar_ready,
  input  wire [31:0]   io_inputs_1_ar_payload_addr,
  input  wire [5:0]    io_inputs_1_ar_payload_id,
  input  wire [3:0]    io_inputs_1_ar_payload_region,
  input  wire [7:0]    io_inputs_1_ar_payload_len,
  input  wire [2:0]    io_inputs_1_ar_payload_size,
  input  wire [1:0]    io_inputs_1_ar_payload_burst,
  input  wire [0:0]    io_inputs_1_ar_payload_lock,
  input  wire [3:0]    io_inputs_1_ar_payload_cache,
  input  wire [3:0]    io_inputs_1_ar_payload_qos,
  input  wire [2:0]    io_inputs_1_ar_payload_prot,
  output wire          io_inputs_1_r_valid,
  input  wire          io_inputs_1_r_ready,
  output wire [127:0]  io_inputs_1_r_payload_data,
  output wire [5:0]    io_inputs_1_r_payload_id,
  output wire [1:0]    io_inputs_1_r_payload_resp,
  output wire          io_inputs_1_r_payload_last,
  input  wire          io_inputs_2_ar_valid,
  output wire          io_inputs_2_ar_ready,
  input  wire [31:0]   io_inputs_2_ar_payload_addr,
  input  wire [5:0]    io_inputs_2_ar_payload_id,
  input  wire [3:0]    io_inputs_2_ar_payload_region,
  input  wire [7:0]    io_inputs_2_ar_payload_len,
  input  wire [2:0]    io_inputs_2_ar_payload_size,
  input  wire [1:0]    io_inputs_2_ar_payload_burst,
  input  wire [0:0]    io_inputs_2_ar_payload_lock,
  input  wire [3:0]    io_inputs_2_ar_payload_cache,
  input  wire [3:0]    io_inputs_2_ar_payload_qos,
  input  wire [2:0]    io_inputs_2_ar_payload_prot,
  output wire          io_inputs_2_r_valid,
  input  wire          io_inputs_2_r_ready,
  output wire [127:0]  io_inputs_2_r_payload_data,
  output wire [5:0]    io_inputs_2_r_payload_id,
  output wire [1:0]    io_inputs_2_r_payload_resp,
  output wire          io_inputs_2_r_payload_last,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [7:0]    io_output_ar_payload_id,
  output wire [3:0]    io_output_ar_payload_region,
  output wire [7:0]    io_output_ar_payload_len,
  output wire [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  output wire [0:0]    io_output_ar_payload_lock,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [3:0]    io_output_ar_payload_qos,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [127:0]  io_output_r_payload_data,
  input  wire [7:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_inputs_2_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [31:0]   cmdArbiter_io_output_payload_addr;
  wire       [5:0]    cmdArbiter_io_output_payload_id;
  wire       [3:0]    cmdArbiter_io_output_payload_region;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire       [0:0]    cmdArbiter_io_output_payload_lock;
  wire       [3:0]    cmdArbiter_io_output_payload_cache;
  wire       [3:0]    cmdArbiter_io_output_payload_qos;
  wire       [2:0]    cmdArbiter_io_output_payload_prot;
  wire       [1:0]    cmdArbiter_io_chosen;
  wire       [2:0]    cmdArbiter_io_chosenOH;
  reg                 _zz_io_output_r_ready;
  wire       [1:0]    readRspIndex;
  wire                readRspSels_0;
  wire                readRspSels_1;
  wire                readRspSels_2;

  StreamArbiter_7 cmdArbiter (
    .io_inputs_0_valid          (io_inputs_0_ar_valid                    ), //i
    .io_inputs_0_ready          (cmdArbiter_io_inputs_0_ready            ), //o
    .io_inputs_0_payload_addr   (io_inputs_0_ar_payload_addr[31:0]       ), //i
    .io_inputs_0_payload_id     (io_inputs_0_ar_payload_id[5:0]          ), //i
    .io_inputs_0_payload_region (io_inputs_0_ar_payload_region[3:0]      ), //i
    .io_inputs_0_payload_len    (io_inputs_0_ar_payload_len[7:0]         ), //i
    .io_inputs_0_payload_size   (io_inputs_0_ar_payload_size[2:0]        ), //i
    .io_inputs_0_payload_burst  (io_inputs_0_ar_payload_burst[1:0]       ), //i
    .io_inputs_0_payload_lock   (io_inputs_0_ar_payload_lock             ), //i
    .io_inputs_0_payload_cache  (io_inputs_0_ar_payload_cache[3:0]       ), //i
    .io_inputs_0_payload_qos    (io_inputs_0_ar_payload_qos[3:0]         ), //i
    .io_inputs_0_payload_prot   (io_inputs_0_ar_payload_prot[2:0]        ), //i
    .io_inputs_1_valid          (io_inputs_1_ar_valid                    ), //i
    .io_inputs_1_ready          (cmdArbiter_io_inputs_1_ready            ), //o
    .io_inputs_1_payload_addr   (io_inputs_1_ar_payload_addr[31:0]       ), //i
    .io_inputs_1_payload_id     (io_inputs_1_ar_payload_id[5:0]          ), //i
    .io_inputs_1_payload_region (io_inputs_1_ar_payload_region[3:0]      ), //i
    .io_inputs_1_payload_len    (io_inputs_1_ar_payload_len[7:0]         ), //i
    .io_inputs_1_payload_size   (io_inputs_1_ar_payload_size[2:0]        ), //i
    .io_inputs_1_payload_burst  (io_inputs_1_ar_payload_burst[1:0]       ), //i
    .io_inputs_1_payload_lock   (io_inputs_1_ar_payload_lock             ), //i
    .io_inputs_1_payload_cache  (io_inputs_1_ar_payload_cache[3:0]       ), //i
    .io_inputs_1_payload_qos    (io_inputs_1_ar_payload_qos[3:0]         ), //i
    .io_inputs_1_payload_prot   (io_inputs_1_ar_payload_prot[2:0]        ), //i
    .io_inputs_2_valid          (io_inputs_2_ar_valid                    ), //i
    .io_inputs_2_ready          (cmdArbiter_io_inputs_2_ready            ), //o
    .io_inputs_2_payload_addr   (io_inputs_2_ar_payload_addr[31:0]       ), //i
    .io_inputs_2_payload_id     (io_inputs_2_ar_payload_id[5:0]          ), //i
    .io_inputs_2_payload_region (io_inputs_2_ar_payload_region[3:0]      ), //i
    .io_inputs_2_payload_len    (io_inputs_2_ar_payload_len[7:0]         ), //i
    .io_inputs_2_payload_size   (io_inputs_2_ar_payload_size[2:0]        ), //i
    .io_inputs_2_payload_burst  (io_inputs_2_ar_payload_burst[1:0]       ), //i
    .io_inputs_2_payload_lock   (io_inputs_2_ar_payload_lock             ), //i
    .io_inputs_2_payload_cache  (io_inputs_2_ar_payload_cache[3:0]       ), //i
    .io_inputs_2_payload_qos    (io_inputs_2_ar_payload_qos[3:0]         ), //i
    .io_inputs_2_payload_prot   (io_inputs_2_ar_payload_prot[2:0]        ), //i
    .io_output_valid            (cmdArbiter_io_output_valid              ), //o
    .io_output_ready            (io_output_ar_ready                      ), //i
    .io_output_payload_addr     (cmdArbiter_io_output_payload_addr[31:0] ), //o
    .io_output_payload_id       (cmdArbiter_io_output_payload_id[5:0]    ), //o
    .io_output_payload_region   (cmdArbiter_io_output_payload_region[3:0]), //o
    .io_output_payload_len      (cmdArbiter_io_output_payload_len[7:0]   ), //o
    .io_output_payload_size     (cmdArbiter_io_output_payload_size[2:0]  ), //o
    .io_output_payload_burst    (cmdArbiter_io_output_payload_burst[1:0] ), //o
    .io_output_payload_lock     (cmdArbiter_io_output_payload_lock       ), //o
    .io_output_payload_cache    (cmdArbiter_io_output_payload_cache[3:0] ), //o
    .io_output_payload_qos      (cmdArbiter_io_output_payload_qos[3:0]   ), //o
    .io_output_payload_prot     (cmdArbiter_io_output_payload_prot[2:0]  ), //o
    .io_chosen                  (cmdArbiter_io_chosen[1:0]               ), //o
    .io_chosenOH                (cmdArbiter_io_chosenOH[2:0]             ), //o
    .io_memoryClk               (io_memoryClk                            ), //i
    .ddrCd_logic_outputReset    (ddrCd_logic_outputReset                 )  //i
  );
  always @(*) begin
    case(readRspIndex)
      2'b00 : _zz_io_output_r_ready = io_inputs_0_r_ready;
      2'b01 : _zz_io_output_r_ready = io_inputs_1_r_ready;
      default : _zz_io_output_r_ready = io_inputs_2_r_ready;
    endcase
  end

  assign io_inputs_0_ar_ready = cmdArbiter_io_inputs_0_ready;
  assign io_inputs_1_ar_ready = cmdArbiter_io_inputs_1_ready;
  assign io_inputs_2_ar_ready = cmdArbiter_io_inputs_2_ready;
  assign io_output_ar_valid = cmdArbiter_io_output_valid;
  assign io_output_ar_payload_addr = cmdArbiter_io_output_payload_addr;
  assign io_output_ar_payload_region = cmdArbiter_io_output_payload_region;
  assign io_output_ar_payload_len = cmdArbiter_io_output_payload_len;
  assign io_output_ar_payload_size = cmdArbiter_io_output_payload_size;
  assign io_output_ar_payload_burst = cmdArbiter_io_output_payload_burst;
  assign io_output_ar_payload_lock = cmdArbiter_io_output_payload_lock;
  assign io_output_ar_payload_cache = cmdArbiter_io_output_payload_cache;
  assign io_output_ar_payload_qos = cmdArbiter_io_output_payload_qos;
  assign io_output_ar_payload_prot = cmdArbiter_io_output_payload_prot;
  assign io_output_ar_payload_id = {cmdArbiter_io_chosen,cmdArbiter_io_output_payload_id};
  assign readRspIndex = io_output_r_payload_id[7 : 6];
  assign readRspSels_0 = (readRspIndex == 2'b00);
  assign readRspSels_1 = (readRspIndex == 2'b01);
  assign readRspSels_2 = (readRspIndex == 2'b10);
  assign io_inputs_0_r_valid = (io_output_r_valid && readRspSels_0);
  assign io_inputs_0_r_payload_data = io_output_r_payload_data;
  assign io_inputs_0_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_0_r_payload_last = io_output_r_payload_last;
  assign io_inputs_0_r_payload_id = io_output_r_payload_id[5 : 0];
  assign io_inputs_1_r_valid = (io_output_r_valid && readRspSels_1);
  assign io_inputs_1_r_payload_data = io_output_r_payload_data;
  assign io_inputs_1_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_1_r_payload_last = io_output_r_payload_last;
  assign io_inputs_1_r_payload_id = io_output_r_payload_id[5 : 0];
  assign io_inputs_2_r_valid = (io_output_r_valid && readRspSels_2);
  assign io_inputs_2_r_payload_data = io_output_r_payload_data;
  assign io_inputs_2_r_payload_resp = io_output_r_payload_resp;
  assign io_inputs_2_r_payload_last = io_output_r_payload_last;
  assign io_inputs_2_r_payload_id = io_output_r_payload_id[5 : 0];
  assign io_output_r_ready = _zz_io_output_r_ready;

endmodule

module BmbCcFifo (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [127:0]  io_input_cmd_payload_fragment_data,
  input  wire [15:0]   io_input_cmd_payload_fragment_mask,
  input  wire [45:0]   io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [127:0]  io_input_rsp_payload_fragment_data,
  output wire [45:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [1:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output wire [127:0]  io_output_cmd_payload_fragment_data,
  output wire [15:0]   io_output_cmd_payload_fragment_mask,
  output wire [45:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [1:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [127:0]  io_output_rsp_payload_fragment_data,
  input  wire [45:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                io_input_cmd_queue_io_push_ready;
  wire                io_input_cmd_queue_io_pop_valid;
  wire                io_input_cmd_queue_io_pop_payload_last;
  wire       [1:0]    io_input_cmd_queue_io_pop_payload_fragment_source;
  wire       [0:0]    io_input_cmd_queue_io_pop_payload_fragment_opcode;
  wire       [31:0]   io_input_cmd_queue_io_pop_payload_fragment_address;
  wire       [5:0]    io_input_cmd_queue_io_pop_payload_fragment_length;
  wire       [127:0]  io_input_cmd_queue_io_pop_payload_fragment_data;
  wire       [15:0]   io_input_cmd_queue_io_pop_payload_fragment_mask;
  wire       [45:0]   io_input_cmd_queue_io_pop_payload_fragment_context;
  wire       [6:0]    io_input_cmd_queue_io_pushOccupancy;
  wire       [6:0]    io_input_cmd_queue_io_popOccupancy;
  wire                io_output_rsp_queue_io_push_ready;
  wire                io_output_rsp_queue_io_pop_valid;
  wire                io_output_rsp_queue_io_pop_payload_last;
  wire       [1:0]    io_output_rsp_queue_io_pop_payload_fragment_source;
  wire       [0:0]    io_output_rsp_queue_io_pop_payload_fragment_opcode;
  wire       [127:0]  io_output_rsp_queue_io_pop_payload_fragment_data;
  wire       [45:0]   io_output_rsp_queue_io_pop_payload_fragment_context;
  wire       [6:0]    io_output_rsp_queue_io_pushOccupancy;
  wire       [6:0]    io_output_rsp_queue_io_popOccupancy;

  StreamFifoCC io_input_cmd_queue (
    .io_push_valid                    (io_input_cmd_valid                                      ), //i
    .io_push_ready                    (io_input_cmd_queue_io_push_ready                        ), //o
    .io_push_payload_last             (io_input_cmd_payload_last                               ), //i
    .io_push_payload_fragment_source  (io_input_cmd_payload_fragment_source[1:0]               ), //i
    .io_push_payload_fragment_opcode  (io_input_cmd_payload_fragment_opcode                    ), //i
    .io_push_payload_fragment_address (io_input_cmd_payload_fragment_address[31:0]             ), //i
    .io_push_payload_fragment_length  (io_input_cmd_payload_fragment_length[5:0]               ), //i
    .io_push_payload_fragment_data    (io_input_cmd_payload_fragment_data[127:0]               ), //i
    .io_push_payload_fragment_mask    (io_input_cmd_payload_fragment_mask[15:0]                ), //i
    .io_push_payload_fragment_context (io_input_cmd_payload_fragment_context[45:0]             ), //i
    .io_pop_valid                     (io_input_cmd_queue_io_pop_valid                         ), //o
    .io_pop_ready                     (io_output_cmd_ready                                     ), //i
    .io_pop_payload_last              (io_input_cmd_queue_io_pop_payload_last                  ), //o
    .io_pop_payload_fragment_source   (io_input_cmd_queue_io_pop_payload_fragment_source[1:0]  ), //o
    .io_pop_payload_fragment_opcode   (io_input_cmd_queue_io_pop_payload_fragment_opcode       ), //o
    .io_pop_payload_fragment_address  (io_input_cmd_queue_io_pop_payload_fragment_address[31:0]), //o
    .io_pop_payload_fragment_length   (io_input_cmd_queue_io_pop_payload_fragment_length[5:0]  ), //o
    .io_pop_payload_fragment_data     (io_input_cmd_queue_io_pop_payload_fragment_data[127:0]  ), //o
    .io_pop_payload_fragment_mask     (io_input_cmd_queue_io_pop_payload_fragment_mask[15:0]   ), //o
    .io_pop_payload_fragment_context  (io_input_cmd_queue_io_pop_payload_fragment_context[45:0]), //o
    .io_pushOccupancy                 (io_input_cmd_queue_io_pushOccupancy[6:0]                ), //o
    .io_popOccupancy                  (io_input_cmd_queue_io_popOccupancy[6:0]                 ), //o
    .io_systemClk                     (io_systemClk                                            ), //i
    .systemCd_logic_outputReset       (systemCd_logic_outputReset                              ), //i
    .io_memoryClk                     (io_memoryClk                                            )  //i
  );
  StreamFifoCC_1 io_output_rsp_queue (
    .io_push_valid                    (io_output_rsp_valid                                      ), //i
    .io_push_ready                    (io_output_rsp_queue_io_push_ready                        ), //o
    .io_push_payload_last             (io_output_rsp_payload_last                               ), //i
    .io_push_payload_fragment_source  (io_output_rsp_payload_fragment_source[1:0]               ), //i
    .io_push_payload_fragment_opcode  (io_output_rsp_payload_fragment_opcode                    ), //i
    .io_push_payload_fragment_data    (io_output_rsp_payload_fragment_data[127:0]               ), //i
    .io_push_payload_fragment_context (io_output_rsp_payload_fragment_context[45:0]             ), //i
    .io_pop_valid                     (io_output_rsp_queue_io_pop_valid                         ), //o
    .io_pop_ready                     (io_input_rsp_ready                                       ), //i
    .io_pop_payload_last              (io_output_rsp_queue_io_pop_payload_last                  ), //o
    .io_pop_payload_fragment_source   (io_output_rsp_queue_io_pop_payload_fragment_source[1:0]  ), //o
    .io_pop_payload_fragment_opcode   (io_output_rsp_queue_io_pop_payload_fragment_opcode       ), //o
    .io_pop_payload_fragment_data     (io_output_rsp_queue_io_pop_payload_fragment_data[127:0]  ), //o
    .io_pop_payload_fragment_context  (io_output_rsp_queue_io_pop_payload_fragment_context[45:0]), //o
    .io_pushOccupancy                 (io_output_rsp_queue_io_pushOccupancy[6:0]                ), //o
    .io_popOccupancy                  (io_output_rsp_queue_io_popOccupancy[6:0]                 ), //o
    .io_memoryClk                     (io_memoryClk                                             ), //i
    .ddrCd_logic_outputReset          (ddrCd_logic_outputReset                                  ), //i
    .io_systemClk                     (io_systemClk                                             )  //i
  );
  assign io_input_cmd_ready = io_input_cmd_queue_io_push_ready;
  assign io_output_cmd_valid = io_input_cmd_queue_io_pop_valid;
  assign io_output_cmd_payload_last = io_input_cmd_queue_io_pop_payload_last;
  assign io_output_cmd_payload_fragment_source = io_input_cmd_queue_io_pop_payload_fragment_source;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_queue_io_pop_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_queue_io_pop_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_queue_io_pop_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = io_input_cmd_queue_io_pop_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = io_input_cmd_queue_io_pop_payload_fragment_mask;
  assign io_output_cmd_payload_fragment_context = io_input_cmd_queue_io_pop_payload_fragment_context;
  assign io_output_rsp_ready = io_output_rsp_queue_io_push_ready;
  assign io_input_rsp_valid = io_output_rsp_queue_io_pop_valid;
  assign io_input_rsp_payload_last = io_output_rsp_queue_io_pop_payload_last;
  assign io_input_rsp_payload_fragment_source = io_output_rsp_queue_io_pop_payload_fragment_source;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_queue_io_pop_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_queue_io_pop_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = io_output_rsp_queue_io_pop_payload_fragment_context;

endmodule

module BmbToAxi4SharedBridge (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [127:0]  io_input_cmd_payload_fragment_data,
  input  wire [15:0]   io_input_cmd_payload_fragment_mask,
  input  wire [45:0]   io_input_cmd_payload_fragment_context,
  output reg           io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output reg           io_input_rsp_payload_last,
  output reg  [1:0]    io_input_rsp_payload_fragment_source,
  output reg  [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [127:0]  io_input_rsp_payload_fragment_data,
  output reg  [45:0]   io_input_rsp_payload_fragment_context,
  output wire          io_output_arw_valid,
  input  wire          io_output_arw_ready,
  output wire [31:0]   io_output_arw_payload_addr,
  output wire [7:0]    io_output_arw_payload_len,
  output wire [2:0]    io_output_arw_payload_size,
  output wire [3:0]    io_output_arw_payload_cache,
  output wire [2:0]    io_output_arw_payload_prot,
  output wire          io_output_arw_payload_write,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [127:0]  io_output_w_payload_data,
  output wire [15:0]   io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [127:0]  io_output_r_payload_data,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                readCmdInfo_fifo_io_pop_ready;
  wire                writeCmdInfo_fifo_io_push_ready;
  wire                writeCmdInfo_fifo_io_pop_valid;
  wire       [1:0]    writeCmdInfo_fifo_io_pop_payload_source;
  wire       [45:0]   writeCmdInfo_fifo_io_pop_payload_context;
  wire       [6:0]    writeCmdInfo_fifo_io_occupancy;
  wire       [6:0]    writeCmdInfo_fifo_io_availability;
  wire                readCmdInfo_fifo_io_push_ready;
  wire                readCmdInfo_fifo_io_pop_valid;
  wire       [1:0]    readCmdInfo_fifo_io_pop_payload_source;
  wire       [45:0]   readCmdInfo_fifo_io_pop_payload_context;
  wire       [6:0]    readCmdInfo_fifo_io_occupancy;
  wire       [6:0]    readCmdInfo_fifo_io_availability;
  wire       [1:0]    _zz_io_output_arw_payload_len;
  reg                 pendingWrite;
  reg        [5:0]    pendingCounter;
  wire                io_input_cmd_fire;
  wire                when_Utils_l706;
  wire                io_input_rsp_fire;
  wire                when_Utils_l709;
  reg                 states_0_counter_incrementIt;
  reg                 states_0_counter_decrementIt;
  wire       [5:0]    states_0_counter_valueNext;
  reg        [5:0]    states_0_counter_value;
  wire                states_0_counter_mayOverflow;
  wire                states_0_counter_willOverflowIfInc;
  wire                states_0_counter_willOverflow;
  reg        [5:0]    states_0_counter_finalIncrement;
  wire                when_Utils_l735;
  wire                when_Utils_l737;
  wire                when_BmbToAxi4Bridge_l45;
  reg                 states_0_write;
  wire                when_BmbToAxi4Bridge_l47;
  wire                when_Utils_l706_1;
  wire                when_Utils_l709_1;
  reg                 states_1_counter_incrementIt;
  reg                 states_1_counter_decrementIt;
  wire       [5:0]    states_1_counter_valueNext;
  reg        [5:0]    states_1_counter_value;
  wire                states_1_counter_mayOverflow;
  wire                states_1_counter_willOverflowIfInc;
  wire                states_1_counter_willOverflow;
  reg        [5:0]    states_1_counter_finalIncrement;
  wire                when_Utils_l735_1;
  wire                when_Utils_l737_1;
  wire                when_BmbToAxi4Bridge_l45_1;
  reg                 states_1_write;
  wire                when_BmbToAxi4Bridge_l47_1;
  wire                when_Utils_l706_2;
  wire                when_Utils_l709_2;
  reg                 states_2_counter_incrementIt;
  reg                 states_2_counter_decrementIt;
  wire       [5:0]    states_2_counter_valueNext;
  reg        [5:0]    states_2_counter_value;
  wire                states_2_counter_mayOverflow;
  wire                states_2_counter_willOverflowIfInc;
  wire                states_2_counter_willOverflow;
  reg        [5:0]    states_2_counter_finalIncrement;
  wire                when_Utils_l735_2;
  wire                when_Utils_l737_2;
  wire                when_BmbToAxi4Bridge_l45_2;
  reg                 states_2_write;
  wire                when_BmbToAxi4Bridge_l47_2;
  wire                when_Utils_l706_3;
  wire                when_Utils_l709_3;
  reg                 states_3_counter_incrementIt;
  reg                 states_3_counter_decrementIt;
  wire       [5:0]    states_3_counter_valueNext;
  reg        [5:0]    states_3_counter_value;
  wire                states_3_counter_mayOverflow;
  wire                states_3_counter_willOverflowIfInc;
  wire                states_3_counter_willOverflow;
  reg        [5:0]    states_3_counter_finalIncrement;
  wire                when_Utils_l735_3;
  wire                when_Utils_l737_3;
  wire                when_BmbToAxi4Bridge_l45_3;
  reg                 states_3_write;
  wire                when_BmbToAxi4Bridge_l47_3;
  wire                hazard;
  wire                _zz_io_input_cmd_ready;
  wire                _zz_cmdFork_valid;
  reg                 _zz_io_input_cmd_ready_1;
  wire                _zz_cmdFork_payload_last;
  wire       [1:0]    _zz_cmdFork_payload_fragment_source;
  wire       [0:0]    _zz_cmdFork_payload_fragment_opcode;
  wire       [31:0]   _zz_cmdFork_payload_fragment_address;
  wire       [5:0]    _zz_cmdFork_payload_fragment_length;
  wire       [127:0]  _zz_cmdFork_payload_fragment_data;
  wire       [15:0]   _zz_cmdFork_payload_fragment_mask;
  wire       [45:0]   _zz_cmdFork_payload_fragment_context;
  wire                cmdFork_valid;
  reg                 cmdFork_ready;
  wire                cmdFork_payload_last;
  wire       [1:0]    cmdFork_payload_fragment_source;
  wire       [0:0]    cmdFork_payload_fragment_opcode;
  wire       [31:0]   cmdFork_payload_fragment_address;
  wire       [5:0]    cmdFork_payload_fragment_length;
  wire       [127:0]  cmdFork_payload_fragment_data;
  wire       [15:0]   cmdFork_payload_fragment_mask;
  wire       [45:0]   cmdFork_payload_fragment_context;
  wire                dataFork_valid;
  reg                 dataFork_ready;
  wire                dataFork_payload_last;
  wire       [1:0]    dataFork_payload_fragment_source;
  wire       [0:0]    dataFork_payload_fragment_opcode;
  wire       [31:0]   dataFork_payload_fragment_address;
  wire       [5:0]    dataFork_payload_fragment_length;
  wire       [127:0]  dataFork_payload_fragment_data;
  wire       [15:0]   dataFork_payload_fragment_mask;
  wire       [45:0]   dataFork_payload_fragment_context;
  reg                 _zz_cmdFork_valid_1;
  reg                 _zz_dataFork_valid;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdFork_fire;
  wire                dataFork_fire;
  reg                 io_input_cmd_payload_first;
  wire                when_Stream_l445;
  reg                 cmdStage_valid;
  wire                cmdStage_ready;
  wire                cmdStage_payload_last;
  wire       [1:0]    cmdStage_payload_fragment_source;
  wire       [0:0]    cmdStage_payload_fragment_opcode;
  wire       [31:0]   cmdStage_payload_fragment_address;
  wire       [5:0]    cmdStage_payload_fragment_length;
  wire       [127:0]  cmdStage_payload_fragment_data;
  wire       [15:0]   cmdStage_payload_fragment_mask;
  wire       [45:0]   cmdStage_payload_fragment_context;
  wire                when_Stream_l445_1;
  reg                 dataStage_valid;
  wire                dataStage_ready;
  wire                dataStage_payload_last;
  wire       [1:0]    dataStage_payload_fragment_source;
  wire       [0:0]    dataStage_payload_fragment_opcode;
  wire       [31:0]   dataStage_payload_fragment_address;
  wire       [5:0]    dataStage_payload_fragment_length;
  wire       [127:0]  dataStage_payload_fragment_data;
  wire       [15:0]   dataStage_payload_fragment_mask;
  wire       [45:0]   dataStage_payload_fragment_context;
  wire                writeCmdInfo_valid;
  wire                writeCmdInfo_ready;
  wire       [1:0]    writeCmdInfo_payload_source;
  wire       [45:0]   writeCmdInfo_payload_context;
  wire                readCmdInfo_valid;
  wire                readCmdInfo_ready;
  wire       [1:0]    readCmdInfo_payload_source;
  wire       [45:0]   readCmdInfo_payload_context;
  wire                cmdStage_fire;
  wire                writeCmdInfo_fifo_io_pop_s2mPipe_valid;
  reg                 writeCmdInfo_fifo_io_pop_s2mPipe_ready;
  wire       [1:0]    writeCmdInfo_fifo_io_pop_s2mPipe_payload_source;
  wire       [45:0]   writeCmdInfo_fifo_io_pop_s2mPipe_payload_context;
  reg                 writeCmdInfo_fifo_io_pop_rValidN;
  reg        [1:0]    writeCmdInfo_fifo_io_pop_rData_source;
  reg        [45:0]   writeCmdInfo_fifo_io_pop_rData_context;
  wire                writeRspInfo_valid;
  wire                writeRspInfo_ready;
  wire       [1:0]    writeRspInfo_payload_source;
  wire       [45:0]   writeRspInfo_payload_context;
  reg                 writeCmdInfo_fifo_io_pop_s2mPipe_rValid;
  reg        [1:0]    writeCmdInfo_fifo_io_pop_s2mPipe_rData_source;
  reg        [45:0]   writeCmdInfo_fifo_io_pop_s2mPipe_rData_context;
  wire                when_Stream_l375;
  wire                readRspInfo_valid;
  wire                readRspInfo_ready;
  wire       [1:0]    readRspInfo_payload_source;
  wire       [45:0]   readRspInfo_payload_context;
  reg                 readCmdInfo_fifo_io_pop_rValid;
  wire                readRspInfo_fire;
  reg        [1:0]    readCmdInfo_fifo_io_pop_rData_source;
  reg        [45:0]   readCmdInfo_fifo_io_pop_rData_context;
  wire                _zz_io_output_arw_valid;
  reg                 rspSelLock;
  wire                when_BmbToAxi4Bridge_l87;
  wire                io_output_r_fire;
  wire                io_output_b_fire;
  wire                when_BmbToAxi4Bridge_l87_1;
  wire                when_BmbToAxi4Bridge_l88;
  reg                 rspSelReadLast;
  wire                rspSelRead;
  wire                when_BmbToAxi4Bridge_l108;

  assign _zz_io_output_arw_payload_len = io_input_cmd_payload_fragment_length[5 : 4];
  StreamFifo_1 writeCmdInfo_fifo (
    .io_push_valid           (writeCmdInfo_valid                            ), //i
    .io_push_ready           (writeCmdInfo_fifo_io_push_ready               ), //o
    .io_push_payload_source  (writeCmdInfo_payload_source[1:0]              ), //i
    .io_push_payload_context (writeCmdInfo_payload_context[45:0]            ), //i
    .io_pop_valid            (writeCmdInfo_fifo_io_pop_valid                ), //o
    .io_pop_ready            (writeCmdInfo_fifo_io_pop_rValidN              ), //i
    .io_pop_payload_source   (writeCmdInfo_fifo_io_pop_payload_source[1:0]  ), //o
    .io_pop_payload_context  (writeCmdInfo_fifo_io_pop_payload_context[45:0]), //o
    .io_flush                (1'b0                                          ), //i
    .io_occupancy            (writeCmdInfo_fifo_io_occupancy[6:0]           ), //o
    .io_availability         (writeCmdInfo_fifo_io_availability[6:0]        ), //o
    .io_memoryClk            (io_memoryClk                                  ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                       )  //i
  );
  StreamFifo_1 readCmdInfo_fifo (
    .io_push_valid           (readCmdInfo_valid                            ), //i
    .io_push_ready           (readCmdInfo_fifo_io_push_ready               ), //o
    .io_push_payload_source  (readCmdInfo_payload_source[1:0]              ), //i
    .io_push_payload_context (readCmdInfo_payload_context[45:0]            ), //i
    .io_pop_valid            (readCmdInfo_fifo_io_pop_valid                ), //o
    .io_pop_ready            (readCmdInfo_fifo_io_pop_ready                ), //i
    .io_pop_payload_source   (readCmdInfo_fifo_io_pop_payload_source[1:0]  ), //o
    .io_pop_payload_context  (readCmdInfo_fifo_io_pop_payload_context[45:0]), //o
    .io_flush                (1'b0                                         ), //i
    .io_occupancy            (readCmdInfo_fifo_io_occupancy[6:0]           ), //o
    .io_availability         (readCmdInfo_fifo_io_availability[6:0]        ), //o
    .io_memoryClk            (io_memoryClk                                 ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                      )  //i
  );
  always @(*) begin
    pendingWrite = 1'bx;
    if(when_BmbToAxi4Bridge_l47) begin
      pendingWrite = states_0_write;
    end
    if(when_BmbToAxi4Bridge_l47_1) begin
      pendingWrite = states_1_write;
    end
    if(when_BmbToAxi4Bridge_l47_2) begin
      pendingWrite = states_2_write;
    end
    if(when_BmbToAxi4Bridge_l47_3) begin
      pendingWrite = states_3_write;
    end
  end

  always @(*) begin
    pendingCounter = 6'bxxxxxx;
    if(when_BmbToAxi4Bridge_l47) begin
      pendingCounter = states_0_counter_value;
    end
    if(when_BmbToAxi4Bridge_l47_1) begin
      pendingCounter = states_1_counter_value;
    end
    if(when_BmbToAxi4Bridge_l47_2) begin
      pendingCounter = states_2_counter_value;
    end
    if(when_BmbToAxi4Bridge_l47_3) begin
      pendingCounter = states_3_counter_value;
    end
  end

  assign io_input_cmd_fire = (io_input_cmd_valid && io_input_cmd_ready);
  assign when_Utils_l706 = (((io_input_cmd_payload_fragment_source == 2'b00) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign io_input_rsp_fire = (io_input_rsp_valid && io_input_rsp_ready);
  assign when_Utils_l709 = (((io_input_rsp_payload_fragment_source == 2'b00) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_0_counter_incrementIt = 1'b0;
    if(when_Utils_l706) begin
      states_0_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_0_counter_decrementIt = 1'b0;
    if(when_Utils_l709) begin
      states_0_counter_decrementIt = 1'b1;
    end
  end

  assign states_0_counter_mayOverflow = (states_0_counter_value == 6'h3f);
  assign states_0_counter_willOverflowIfInc = (states_0_counter_mayOverflow && (! states_0_counter_decrementIt));
  assign states_0_counter_willOverflow = (states_0_counter_willOverflowIfInc && states_0_counter_incrementIt);
  assign when_Utils_l735 = (states_0_counter_incrementIt && (! states_0_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735) begin
      states_0_counter_finalIncrement = 6'h01;
    end else begin
      if(when_Utils_l737) begin
        states_0_counter_finalIncrement = 6'h3f;
      end else begin
        states_0_counter_finalIncrement = 6'h0;
      end
    end
  end

  assign when_Utils_l737 = ((! states_0_counter_incrementIt) && states_0_counter_decrementIt);
  assign states_0_counter_valueNext = (states_0_counter_value + states_0_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45 = ((io_input_cmd_payload_fragment_source == 2'b00) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47 = (io_input_cmd_payload_fragment_source == 2'b00);
  assign when_Utils_l706_1 = (((io_input_cmd_payload_fragment_source == 2'b10) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign when_Utils_l709_1 = (((io_input_rsp_payload_fragment_source == 2'b10) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_1_counter_incrementIt = 1'b0;
    if(when_Utils_l706_1) begin
      states_1_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_1_counter_decrementIt = 1'b0;
    if(when_Utils_l709_1) begin
      states_1_counter_decrementIt = 1'b1;
    end
  end

  assign states_1_counter_mayOverflow = (states_1_counter_value == 6'h3f);
  assign states_1_counter_willOverflowIfInc = (states_1_counter_mayOverflow && (! states_1_counter_decrementIt));
  assign states_1_counter_willOverflow = (states_1_counter_willOverflowIfInc && states_1_counter_incrementIt);
  assign when_Utils_l735_1 = (states_1_counter_incrementIt && (! states_1_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_1) begin
      states_1_counter_finalIncrement = 6'h01;
    end else begin
      if(when_Utils_l737_1) begin
        states_1_counter_finalIncrement = 6'h3f;
      end else begin
        states_1_counter_finalIncrement = 6'h0;
      end
    end
  end

  assign when_Utils_l737_1 = ((! states_1_counter_incrementIt) && states_1_counter_decrementIt);
  assign states_1_counter_valueNext = (states_1_counter_value + states_1_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45_1 = ((io_input_cmd_payload_fragment_source == 2'b10) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47_1 = (io_input_cmd_payload_fragment_source == 2'b10);
  assign when_Utils_l706_2 = (((io_input_cmd_payload_fragment_source == 2'b01) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign when_Utils_l709_2 = (((io_input_rsp_payload_fragment_source == 2'b01) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_2_counter_incrementIt = 1'b0;
    if(when_Utils_l706_2) begin
      states_2_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_2_counter_decrementIt = 1'b0;
    if(when_Utils_l709_2) begin
      states_2_counter_decrementIt = 1'b1;
    end
  end

  assign states_2_counter_mayOverflow = (states_2_counter_value == 6'h3f);
  assign states_2_counter_willOverflowIfInc = (states_2_counter_mayOverflow && (! states_2_counter_decrementIt));
  assign states_2_counter_willOverflow = (states_2_counter_willOverflowIfInc && states_2_counter_incrementIt);
  assign when_Utils_l735_2 = (states_2_counter_incrementIt && (! states_2_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_2) begin
      states_2_counter_finalIncrement = 6'h01;
    end else begin
      if(when_Utils_l737_2) begin
        states_2_counter_finalIncrement = 6'h3f;
      end else begin
        states_2_counter_finalIncrement = 6'h0;
      end
    end
  end

  assign when_Utils_l737_2 = ((! states_2_counter_incrementIt) && states_2_counter_decrementIt);
  assign states_2_counter_valueNext = (states_2_counter_value + states_2_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45_2 = ((io_input_cmd_payload_fragment_source == 2'b01) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47_2 = (io_input_cmd_payload_fragment_source == 2'b01);
  assign when_Utils_l706_3 = (((io_input_cmd_payload_fragment_source == 2'b11) && io_input_cmd_fire) && io_input_cmd_payload_last);
  assign when_Utils_l709_3 = (((io_input_rsp_payload_fragment_source == 2'b11) && io_input_rsp_fire) && io_input_rsp_payload_last);
  always @(*) begin
    states_3_counter_incrementIt = 1'b0;
    if(when_Utils_l706_3) begin
      states_3_counter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    states_3_counter_decrementIt = 1'b0;
    if(when_Utils_l709_3) begin
      states_3_counter_decrementIt = 1'b1;
    end
  end

  assign states_3_counter_mayOverflow = (states_3_counter_value == 6'h3f);
  assign states_3_counter_willOverflowIfInc = (states_3_counter_mayOverflow && (! states_3_counter_decrementIt));
  assign states_3_counter_willOverflow = (states_3_counter_willOverflowIfInc && states_3_counter_incrementIt);
  assign when_Utils_l735_3 = (states_3_counter_incrementIt && (! states_3_counter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_3) begin
      states_3_counter_finalIncrement = 6'h01;
    end else begin
      if(when_Utils_l737_3) begin
        states_3_counter_finalIncrement = 6'h3f;
      end else begin
        states_3_counter_finalIncrement = 6'h0;
      end
    end
  end

  assign when_Utils_l737_3 = ((! states_3_counter_incrementIt) && states_3_counter_decrementIt);
  assign states_3_counter_valueNext = (states_3_counter_value + states_3_counter_finalIncrement);
  assign when_BmbToAxi4Bridge_l45_3 = ((io_input_cmd_payload_fragment_source == 2'b11) && io_input_cmd_fire);
  assign when_BmbToAxi4Bridge_l47_3 = (io_input_cmd_payload_fragment_source == 2'b11);
  assign hazard = ((((io_input_cmd_payload_fragment_opcode == 1'b1) != pendingWrite) && (pendingCounter != 6'h0)) || (pendingCounter == 6'h3f));
  assign _zz_io_input_cmd_ready = (! hazard);
  assign _zz_cmdFork_valid = (io_input_cmd_valid && _zz_io_input_cmd_ready);
  assign io_input_cmd_ready = (_zz_io_input_cmd_ready_1 && _zz_io_input_cmd_ready);
  assign _zz_cmdFork_payload_last = io_input_cmd_payload_last;
  assign _zz_cmdFork_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign _zz_cmdFork_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign _zz_cmdFork_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign _zz_cmdFork_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign _zz_cmdFork_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign _zz_cmdFork_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign _zz_cmdFork_payload_fragment_context = io_input_cmd_payload_fragment_context;
  always @(*) begin
    _zz_io_input_cmd_ready_1 = 1'b1;
    if(when_Stream_l1063) begin
      _zz_io_input_cmd_ready_1 = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      _zz_io_input_cmd_ready_1 = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdFork_ready) && _zz_cmdFork_valid_1);
  assign when_Stream_l1063_1 = ((! dataFork_ready) && _zz_dataFork_valid);
  assign cmdFork_valid = (_zz_cmdFork_valid && _zz_cmdFork_valid_1);
  assign cmdFork_payload_last = _zz_cmdFork_payload_last;
  assign cmdFork_payload_fragment_source = _zz_cmdFork_payload_fragment_source;
  assign cmdFork_payload_fragment_opcode = _zz_cmdFork_payload_fragment_opcode;
  assign cmdFork_payload_fragment_address = _zz_cmdFork_payload_fragment_address;
  assign cmdFork_payload_fragment_length = _zz_cmdFork_payload_fragment_length;
  assign cmdFork_payload_fragment_data = _zz_cmdFork_payload_fragment_data;
  assign cmdFork_payload_fragment_mask = _zz_cmdFork_payload_fragment_mask;
  assign cmdFork_payload_fragment_context = _zz_cmdFork_payload_fragment_context;
  assign cmdFork_fire = (cmdFork_valid && cmdFork_ready);
  assign dataFork_valid = (_zz_cmdFork_valid && _zz_dataFork_valid);
  assign dataFork_payload_last = _zz_cmdFork_payload_last;
  assign dataFork_payload_fragment_source = _zz_cmdFork_payload_fragment_source;
  assign dataFork_payload_fragment_opcode = _zz_cmdFork_payload_fragment_opcode;
  assign dataFork_payload_fragment_address = _zz_cmdFork_payload_fragment_address;
  assign dataFork_payload_fragment_length = _zz_cmdFork_payload_fragment_length;
  assign dataFork_payload_fragment_data = _zz_cmdFork_payload_fragment_data;
  assign dataFork_payload_fragment_mask = _zz_cmdFork_payload_fragment_mask;
  assign dataFork_payload_fragment_context = _zz_cmdFork_payload_fragment_context;
  assign dataFork_fire = (dataFork_valid && dataFork_ready);
  assign when_Stream_l445 = (! io_input_cmd_payload_first);
  always @(*) begin
    cmdStage_valid = cmdFork_valid;
    if(when_Stream_l445) begin
      cmdStage_valid = 1'b0;
    end
  end

  always @(*) begin
    cmdFork_ready = cmdStage_ready;
    if(when_Stream_l445) begin
      cmdFork_ready = 1'b1;
    end
  end

  assign cmdStage_payload_last = cmdFork_payload_last;
  assign cmdStage_payload_fragment_source = cmdFork_payload_fragment_source;
  assign cmdStage_payload_fragment_opcode = cmdFork_payload_fragment_opcode;
  assign cmdStage_payload_fragment_address = cmdFork_payload_fragment_address;
  assign cmdStage_payload_fragment_length = cmdFork_payload_fragment_length;
  assign cmdStage_payload_fragment_data = cmdFork_payload_fragment_data;
  assign cmdStage_payload_fragment_mask = cmdFork_payload_fragment_mask;
  assign cmdStage_payload_fragment_context = cmdFork_payload_fragment_context;
  assign when_Stream_l445_1 = (! (dataFork_payload_fragment_opcode == 1'b1));
  always @(*) begin
    dataStage_valid = dataFork_valid;
    if(when_Stream_l445_1) begin
      dataStage_valid = 1'b0;
    end
  end

  always @(*) begin
    dataFork_ready = dataStage_ready;
    if(when_Stream_l445_1) begin
      dataFork_ready = 1'b1;
    end
  end

  assign dataStage_payload_last = dataFork_payload_last;
  assign dataStage_payload_fragment_source = dataFork_payload_fragment_source;
  assign dataStage_payload_fragment_opcode = dataFork_payload_fragment_opcode;
  assign dataStage_payload_fragment_address = dataFork_payload_fragment_address;
  assign dataStage_payload_fragment_length = dataFork_payload_fragment_length;
  assign dataStage_payload_fragment_data = dataFork_payload_fragment_data;
  assign dataStage_payload_fragment_mask = dataFork_payload_fragment_mask;
  assign dataStage_payload_fragment_context = dataFork_payload_fragment_context;
  assign cmdStage_fire = (cmdStage_valid && cmdStage_ready);
  assign writeCmdInfo_valid = (cmdStage_fire && (cmdStage_payload_fragment_opcode == 1'b1));
  assign writeCmdInfo_payload_source = cmdStage_payload_fragment_source;
  assign writeCmdInfo_payload_context = cmdStage_payload_fragment_context;
  assign readCmdInfo_valid = (cmdStage_fire && (cmdStage_payload_fragment_opcode == 1'b0));
  assign readCmdInfo_payload_source = cmdStage_payload_fragment_source;
  assign readCmdInfo_payload_context = cmdStage_payload_fragment_context;
  assign writeCmdInfo_ready = writeCmdInfo_fifo_io_push_ready;
  assign writeCmdInfo_fifo_io_pop_s2mPipe_valid = (writeCmdInfo_fifo_io_pop_valid || (! writeCmdInfo_fifo_io_pop_rValidN));
  assign writeCmdInfo_fifo_io_pop_s2mPipe_payload_source = (writeCmdInfo_fifo_io_pop_rValidN ? writeCmdInfo_fifo_io_pop_payload_source : writeCmdInfo_fifo_io_pop_rData_source);
  assign writeCmdInfo_fifo_io_pop_s2mPipe_payload_context = (writeCmdInfo_fifo_io_pop_rValidN ? writeCmdInfo_fifo_io_pop_payload_context : writeCmdInfo_fifo_io_pop_rData_context);
  always @(*) begin
    writeCmdInfo_fifo_io_pop_s2mPipe_ready = writeRspInfo_ready;
    if(when_Stream_l375) begin
      writeCmdInfo_fifo_io_pop_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! writeRspInfo_valid);
  assign writeRspInfo_valid = writeCmdInfo_fifo_io_pop_s2mPipe_rValid;
  assign writeRspInfo_payload_source = writeCmdInfo_fifo_io_pop_s2mPipe_rData_source;
  assign writeRspInfo_payload_context = writeCmdInfo_fifo_io_pop_s2mPipe_rData_context;
  assign readCmdInfo_ready = readCmdInfo_fifo_io_push_ready;
  assign readRspInfo_fire = (readRspInfo_valid && readRspInfo_ready);
  assign readCmdInfo_fifo_io_pop_ready = (! readCmdInfo_fifo_io_pop_rValid);
  assign readRspInfo_valid = readCmdInfo_fifo_io_pop_rValid;
  assign readRspInfo_payload_source = readCmdInfo_fifo_io_pop_rData_source;
  assign readRspInfo_payload_context = readCmdInfo_fifo_io_pop_rData_context;
  assign _zz_io_output_arw_valid = (! ((! writeCmdInfo_ready) || (! readCmdInfo_ready)));
  assign cmdStage_ready = (io_output_arw_ready && _zz_io_output_arw_valid);
  assign io_output_arw_valid = (cmdStage_valid && _zz_io_output_arw_valid);
  assign io_output_arw_payload_write = (io_input_cmd_payload_fragment_opcode == 1'b1);
  assign io_output_arw_payload_addr = io_input_cmd_payload_fragment_address;
  assign io_output_arw_payload_len = {6'd0, _zz_io_output_arw_payload_len};
  assign io_output_arw_payload_size = 3'b100;
  assign io_output_arw_payload_prot = 3'b010;
  assign io_output_arw_payload_cache = 4'b1111;
  assign io_output_w_valid = dataStage_valid;
  assign dataStage_ready = io_output_w_ready;
  assign io_output_w_payload_data = dataStage_payload_fragment_data;
  assign io_output_w_payload_strb = dataStage_payload_fragment_mask;
  assign io_output_w_payload_last = dataStage_payload_last;
  assign when_BmbToAxi4Bridge_l87 = (io_output_r_valid || io_output_b_valid);
  assign io_output_r_fire = (io_output_r_valid && io_output_r_ready);
  assign io_output_b_fire = (io_output_b_valid && io_output_b_ready);
  assign when_BmbToAxi4Bridge_l87_1 = ((io_output_r_fire && io_output_r_payload_last) || io_output_b_fire);
  assign when_BmbToAxi4Bridge_l88 = (! rspSelLock);
  assign rspSelRead = (rspSelLock ? rspSelReadLast : io_output_r_valid);
  assign io_output_b_ready = ((io_input_rsp_ready && (! rspSelRead)) && writeRspInfo_valid);
  assign io_output_r_ready = ((io_input_rsp_ready && rspSelRead) && readRspInfo_valid);
  assign writeRspInfo_ready = ((io_input_rsp_fire && io_input_rsp_payload_last) && (! rspSelRead));
  assign readRspInfo_ready = ((io_input_rsp_fire && io_input_rsp_payload_last) && rspSelRead);
  assign io_input_rsp_payload_fragment_data = io_output_r_payload_data;
  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_valid = (io_output_r_valid && readRspInfo_valid);
    end else begin
      io_input_rsp_valid = (io_output_b_valid && writeRspInfo_valid);
    end
  end

  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_payload_last = io_output_r_payload_last;
    end else begin
      io_input_rsp_payload_last = 1'b1;
    end
  end

  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_payload_fragment_source = readRspInfo_payload_source;
    end else begin
      io_input_rsp_payload_fragment_source = writeRspInfo_payload_source;
    end
  end

  always @(*) begin
    if(rspSelRead) begin
      io_input_rsp_payload_fragment_context = readRspInfo_payload_context;
    end else begin
      io_input_rsp_payload_fragment_context = writeRspInfo_payload_context;
    end
  end

  assign when_BmbToAxi4Bridge_l108 = (rspSelRead ? (io_output_r_payload_resp == 2'b00) : (io_output_b_payload_resp == 2'b00));
  always @(*) begin
    if(when_BmbToAxi4Bridge_l108) begin
      io_input_rsp_payload_fragment_opcode = 1'b0;
    end else begin
      io_input_rsp_payload_fragment_opcode = 1'b1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      states_0_counter_value <= 6'h0;
      states_1_counter_value <= 6'h0;
      states_2_counter_value <= 6'h0;
      states_3_counter_value <= 6'h0;
      _zz_cmdFork_valid_1 <= 1'b1;
      _zz_dataFork_valid <= 1'b1;
      io_input_cmd_payload_first <= 1'b1;
      writeCmdInfo_fifo_io_pop_rValidN <= 1'b1;
      writeCmdInfo_fifo_io_pop_s2mPipe_rValid <= 1'b0;
      readCmdInfo_fifo_io_pop_rValid <= 1'b0;
      rspSelLock <= 1'b0;
    end else begin
      states_0_counter_value <= states_0_counter_valueNext;
      states_1_counter_value <= states_1_counter_valueNext;
      states_2_counter_value <= states_2_counter_valueNext;
      states_3_counter_value <= states_3_counter_valueNext;
      if(cmdFork_fire) begin
        _zz_cmdFork_valid_1 <= 1'b0;
      end
      if(dataFork_fire) begin
        _zz_dataFork_valid <= 1'b0;
      end
      if(_zz_io_input_cmd_ready_1) begin
        _zz_cmdFork_valid_1 <= 1'b1;
        _zz_dataFork_valid <= 1'b1;
      end
      if(io_input_cmd_fire) begin
        io_input_cmd_payload_first <= io_input_cmd_payload_last;
      end
      if(writeCmdInfo_fifo_io_pop_valid) begin
        writeCmdInfo_fifo_io_pop_rValidN <= 1'b0;
      end
      if(writeCmdInfo_fifo_io_pop_s2mPipe_ready) begin
        writeCmdInfo_fifo_io_pop_rValidN <= 1'b1;
      end
      if(writeCmdInfo_fifo_io_pop_s2mPipe_ready) begin
        writeCmdInfo_fifo_io_pop_s2mPipe_rValid <= writeCmdInfo_fifo_io_pop_s2mPipe_valid;
      end
      if(readCmdInfo_fifo_io_pop_valid) begin
        readCmdInfo_fifo_io_pop_rValid <= 1'b1;
      end
      if(readRspInfo_fire) begin
        readCmdInfo_fifo_io_pop_rValid <= 1'b0;
      end
      if(when_BmbToAxi4Bridge_l87) begin
        rspSelLock <= 1'b1;
      end
      if(when_BmbToAxi4Bridge_l87_1) begin
        rspSelLock <= 1'b0;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(when_BmbToAxi4Bridge_l45) begin
      states_0_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(when_BmbToAxi4Bridge_l45_1) begin
      states_1_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(when_BmbToAxi4Bridge_l45_2) begin
      states_2_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(when_BmbToAxi4Bridge_l45_3) begin
      states_3_write <= (io_input_cmd_payload_fragment_opcode == 1'b1);
    end
    if(writeCmdInfo_fifo_io_pop_rValidN) begin
      writeCmdInfo_fifo_io_pop_rData_source <= writeCmdInfo_fifo_io_pop_payload_source;
      writeCmdInfo_fifo_io_pop_rData_context <= writeCmdInfo_fifo_io_pop_payload_context;
    end
    if(writeCmdInfo_fifo_io_pop_s2mPipe_ready) begin
      writeCmdInfo_fifo_io_pop_s2mPipe_rData_source <= writeCmdInfo_fifo_io_pop_s2mPipe_payload_source;
      writeCmdInfo_fifo_io_pop_s2mPipe_rData_context <= writeCmdInfo_fifo_io_pop_s2mPipe_payload_context;
    end
    if(readCmdInfo_fifo_io_pop_ready) begin
      readCmdInfo_fifo_io_pop_rData_source <= readCmdInfo_fifo_io_pop_payload_source;
      readCmdInfo_fifo_io_pop_rData_context <= readCmdInfo_fifo_io_pop_payload_context;
    end
    if(when_BmbToAxi4Bridge_l88) begin
      rspSelReadLast <= io_output_r_valid;
    end
  end


endmodule

module BmbArbiter_2 (
  input  wire          io_inputs_0_cmd_valid,
  output wire          io_inputs_0_cmd_ready,
  input  wire          io_inputs_0_cmd_payload_last,
  input  wire [0:0]    io_inputs_0_cmd_payload_fragment_source,
  input  wire [0:0]    io_inputs_0_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_0_cmd_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_cmd_payload_fragment_length,
  input  wire [63:0]   io_inputs_0_cmd_payload_fragment_data,
  input  wire [7:0]    io_inputs_0_cmd_payload_fragment_mask,
  input  wire [43:0]   io_inputs_0_cmd_payload_fragment_context,
  output wire          io_inputs_0_rsp_valid,
  input  wire          io_inputs_0_rsp_ready,
  output wire          io_inputs_0_rsp_payload_last,
  output wire [0:0]    io_inputs_0_rsp_payload_fragment_source,
  output wire [0:0]    io_inputs_0_rsp_payload_fragment_opcode,
  output wire [63:0]   io_inputs_0_rsp_payload_fragment_data,
  output wire [43:0]   io_inputs_0_rsp_payload_fragment_context,
  input  wire          io_inputs_1_cmd_valid,
  output wire          io_inputs_1_cmd_ready,
  input  wire          io_inputs_1_cmd_payload_last,
  input  wire [0:0]    io_inputs_1_cmd_payload_fragment_source,
  input  wire [0:0]    io_inputs_1_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_1_cmd_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_cmd_payload_fragment_length,
  input  wire [63:0]   io_inputs_1_cmd_payload_fragment_data,
  input  wire [7:0]    io_inputs_1_cmd_payload_fragment_mask,
  output wire          io_inputs_1_rsp_valid,
  input  wire          io_inputs_1_rsp_ready,
  output wire          io_inputs_1_rsp_payload_last,
  output wire [0:0]    io_inputs_1_rsp_payload_fragment_source,
  output wire [0:0]    io_inputs_1_rsp_payload_fragment_opcode,
  output wire [63:0]   io_inputs_1_rsp_payload_fragment_data,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [1:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output wire [63:0]   io_output_cmd_payload_fragment_data,
  output wire [7:0]    io_output_cmd_payload_fragment_mask,
  output wire [43:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [1:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_output_rsp_payload_fragment_data,
  input  wire [43:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [1:0]    memory_arbiter_io_inputs_0_payload_fragment_source;
  wire       [1:0]    memory_arbiter_io_inputs_1_payload_fragment_source;
  wire                memory_arbiter_io_inputs_0_ready;
  wire                memory_arbiter_io_inputs_1_ready;
  wire                memory_arbiter_io_output_valid;
  wire                memory_arbiter_io_output_payload_last;
  wire       [1:0]    memory_arbiter_io_output_payload_fragment_source;
  wire       [0:0]    memory_arbiter_io_output_payload_fragment_opcode;
  wire       [31:0]   memory_arbiter_io_output_payload_fragment_address;
  wire       [5:0]    memory_arbiter_io_output_payload_fragment_length;
  wire       [63:0]   memory_arbiter_io_output_payload_fragment_data;
  wire       [7:0]    memory_arbiter_io_output_payload_fragment_mask;
  wire       [43:0]   memory_arbiter_io_output_payload_fragment_context;
  wire       [0:0]    memory_arbiter_io_chosen;
  wire       [1:0]    memory_arbiter_io_chosenOH;
  wire       [2:0]    _zz_io_output_cmd_payload_fragment_source;
  reg                 _zz_io_output_rsp_ready;
  wire       [0:0]    memory_rspSel;

  assign _zz_io_output_cmd_payload_fragment_source = {memory_arbiter_io_output_payload_fragment_source,memory_arbiter_io_chosen};
  StreamArbiter_6 memory_arbiter (
    .io_inputs_0_valid                    (io_inputs_0_cmd_valid                                  ), //i
    .io_inputs_0_ready                    (memory_arbiter_io_inputs_0_ready                       ), //o
    .io_inputs_0_payload_last             (io_inputs_0_cmd_payload_last                           ), //i
    .io_inputs_0_payload_fragment_source  (memory_arbiter_io_inputs_0_payload_fragment_source[1:0]), //i
    .io_inputs_0_payload_fragment_opcode  (io_inputs_0_cmd_payload_fragment_opcode                ), //i
    .io_inputs_0_payload_fragment_address (io_inputs_0_cmd_payload_fragment_address[31:0]         ), //i
    .io_inputs_0_payload_fragment_length  (io_inputs_0_cmd_payload_fragment_length[5:0]           ), //i
    .io_inputs_0_payload_fragment_data    (io_inputs_0_cmd_payload_fragment_data[63:0]            ), //i
    .io_inputs_0_payload_fragment_mask    (io_inputs_0_cmd_payload_fragment_mask[7:0]             ), //i
    .io_inputs_0_payload_fragment_context (io_inputs_0_cmd_payload_fragment_context[43:0]         ), //i
    .io_inputs_1_valid                    (io_inputs_1_cmd_valid                                  ), //i
    .io_inputs_1_ready                    (memory_arbiter_io_inputs_1_ready                       ), //o
    .io_inputs_1_payload_last             (io_inputs_1_cmd_payload_last                           ), //i
    .io_inputs_1_payload_fragment_source  (memory_arbiter_io_inputs_1_payload_fragment_source[1:0]), //i
    .io_inputs_1_payload_fragment_opcode  (io_inputs_1_cmd_payload_fragment_opcode                ), //i
    .io_inputs_1_payload_fragment_address (io_inputs_1_cmd_payload_fragment_address[31:0]         ), //i
    .io_inputs_1_payload_fragment_length  (io_inputs_1_cmd_payload_fragment_length[5:0]           ), //i
    .io_inputs_1_payload_fragment_data    (io_inputs_1_cmd_payload_fragment_data[63:0]            ), //i
    .io_inputs_1_payload_fragment_mask    (io_inputs_1_cmd_payload_fragment_mask[7:0]             ), //i
    .io_inputs_1_payload_fragment_context (44'h0                                                  ), //i
    .io_output_valid                      (memory_arbiter_io_output_valid                         ), //o
    .io_output_ready                      (io_output_cmd_ready                                    ), //i
    .io_output_payload_last               (memory_arbiter_io_output_payload_last                  ), //o
    .io_output_payload_fragment_source    (memory_arbiter_io_output_payload_fragment_source[1:0]  ), //o
    .io_output_payload_fragment_opcode    (memory_arbiter_io_output_payload_fragment_opcode       ), //o
    .io_output_payload_fragment_address   (memory_arbiter_io_output_payload_fragment_address[31:0]), //o
    .io_output_payload_fragment_length    (memory_arbiter_io_output_payload_fragment_length[5:0]  ), //o
    .io_output_payload_fragment_data      (memory_arbiter_io_output_payload_fragment_data[63:0]   ), //o
    .io_output_payload_fragment_mask      (memory_arbiter_io_output_payload_fragment_mask[7:0]    ), //o
    .io_output_payload_fragment_context   (memory_arbiter_io_output_payload_fragment_context[43:0]), //o
    .io_chosen                            (memory_arbiter_io_chosen                               ), //o
    .io_chosenOH                          (memory_arbiter_io_chosenOH[1:0]                        ), //o
    .io_systemClk                         (io_systemClk                                           ), //i
    .systemCd_logic_outputReset           (systemCd_logic_outputReset                             )  //i
  );
  always @(*) begin
    case(memory_rspSel)
      1'b0 : _zz_io_output_rsp_ready = io_inputs_0_rsp_ready;
      default : _zz_io_output_rsp_ready = io_inputs_1_rsp_ready;
    endcase
  end

  assign io_inputs_0_cmd_ready = memory_arbiter_io_inputs_0_ready;
  assign memory_arbiter_io_inputs_0_payload_fragment_source = {1'd0, io_inputs_0_cmd_payload_fragment_source};
  assign io_inputs_1_cmd_ready = memory_arbiter_io_inputs_1_ready;
  assign memory_arbiter_io_inputs_1_payload_fragment_source = {1'd0, io_inputs_1_cmd_payload_fragment_source};
  assign io_output_cmd_valid = memory_arbiter_io_output_valid;
  assign io_output_cmd_payload_last = memory_arbiter_io_output_payload_last;
  assign io_output_cmd_payload_fragment_opcode = memory_arbiter_io_output_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = memory_arbiter_io_output_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = memory_arbiter_io_output_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = memory_arbiter_io_output_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = memory_arbiter_io_output_payload_fragment_mask;
  assign io_output_cmd_payload_fragment_context = memory_arbiter_io_output_payload_fragment_context;
  assign io_output_cmd_payload_fragment_source = _zz_io_output_cmd_payload_fragment_source[1:0];
  assign memory_rspSel = io_output_rsp_payload_fragment_source[0 : 0];
  assign io_inputs_0_rsp_valid = (io_output_rsp_valid && (memory_rspSel == 1'b0));
  assign io_inputs_0_rsp_payload_last = io_output_rsp_payload_last;
  assign io_inputs_0_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_inputs_0_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_inputs_0_rsp_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign io_inputs_0_rsp_payload_fragment_source = (io_output_rsp_payload_fragment_source >>> 1'd1);
  assign io_inputs_1_rsp_valid = (io_output_rsp_valid && (memory_rspSel == 1'b1));
  assign io_inputs_1_rsp_payload_last = io_output_rsp_payload_last;
  assign io_inputs_1_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_inputs_1_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_inputs_1_rsp_payload_fragment_source = (io_output_rsp_payload_fragment_source >>> 1'd1);
  assign io_output_rsp_ready = _zz_io_output_rsp_ready;

endmodule

module BmbDecoder (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire          io_outputs_0_cmd_valid,
  input  wire          io_outputs_0_cmd_ready,
  output wire          io_outputs_0_cmd_payload_last,
  output wire [0:0]    io_outputs_0_cmd_payload_fragment_source,
  output wire [0:0]    io_outputs_0_cmd_payload_fragment_opcode,
  output wire [31:0]   io_outputs_0_cmd_payload_fragment_address,
  output wire [5:0]    io_outputs_0_cmd_payload_fragment_length,
  input  wire          io_outputs_0_rsp_valid,
  output wire          io_outputs_0_rsp_ready,
  input  wire          io_outputs_0_rsp_payload_last,
  input  wire [0:0]    io_outputs_0_rsp_payload_fragment_source,
  input  wire [0:0]    io_outputs_0_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_outputs_0_rsp_payload_fragment_data
);


  assign io_outputs_0_cmd_valid = io_input_cmd_valid;
  assign io_input_cmd_ready = io_outputs_0_cmd_ready;
  assign io_input_rsp_valid = io_outputs_0_rsp_valid;
  assign io_outputs_0_rsp_ready = io_input_rsp_ready;
  assign io_outputs_0_cmd_payload_last = io_input_cmd_payload_last;
  assign io_input_rsp_payload_last = io_outputs_0_rsp_payload_last;
  assign io_outputs_0_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_outputs_0_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_outputs_0_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_outputs_0_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_input_rsp_payload_fragment_source = io_outputs_0_rsp_payload_fragment_source;
  assign io_input_rsp_payload_fragment_opcode = io_outputs_0_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_outputs_0_rsp_payload_fragment_data;

endmodule

module BmbArbiter_1 (
  input  wire          io_inputs_0_cmd_valid,
  output wire          io_inputs_0_cmd_ready,
  input  wire          io_inputs_0_cmd_payload_last,
  input  wire [0:0]    io_inputs_0_cmd_payload_fragment_opcode,
  input  wire          io_inputs_0_cmd_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_0_cmd_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_cmd_payload_fragment_length,
  input  wire [63:0]   io_inputs_0_cmd_payload_fragment_data,
  input  wire [7:0]    io_inputs_0_cmd_payload_fragment_mask,
  input  wire [3:0]    io_inputs_0_cmd_payload_fragment_context,
  output wire          io_inputs_0_rsp_valid,
  input  wire          io_inputs_0_rsp_ready,
  output wire          io_inputs_0_rsp_payload_last,
  output wire [0:0]    io_inputs_0_rsp_payload_fragment_opcode,
  output wire          io_inputs_0_rsp_payload_fragment_exclusive,
  output wire [63:0]   io_inputs_0_rsp_payload_fragment_data,
  output wire [3:0]    io_inputs_0_rsp_payload_fragment_context,
  output wire          io_inputs_0_inv_valid,
  input  wire          io_inputs_0_inv_ready,
  output wire          io_inputs_0_inv_payload_all,
  output wire [31:0]   io_inputs_0_inv_payload_address,
  output wire [5:0]    io_inputs_0_inv_payload_length,
  input  wire          io_inputs_0_ack_valid,
  output wire          io_inputs_0_ack_ready,
  output wire          io_inputs_0_sync_valid,
  input  wire          io_inputs_0_sync_ready,
  input  wire          io_inputs_1_cmd_valid,
  output wire          io_inputs_1_cmd_ready,
  input  wire          io_inputs_1_cmd_payload_last,
  input  wire [0:0]    io_inputs_1_cmd_payload_fragment_opcode,
  input  wire          io_inputs_1_cmd_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_1_cmd_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_cmd_payload_fragment_length,
  input  wire [63:0]   io_inputs_1_cmd_payload_fragment_data,
  input  wire [7:0]    io_inputs_1_cmd_payload_fragment_mask,
  input  wire [3:0]    io_inputs_1_cmd_payload_fragment_context,
  output wire          io_inputs_1_rsp_valid,
  input  wire          io_inputs_1_rsp_ready,
  output wire          io_inputs_1_rsp_payload_last,
  output wire [0:0]    io_inputs_1_rsp_payload_fragment_opcode,
  output wire          io_inputs_1_rsp_payload_fragment_exclusive,
  output wire [63:0]   io_inputs_1_rsp_payload_fragment_data,
  output wire [3:0]    io_inputs_1_rsp_payload_fragment_context,
  output wire          io_inputs_1_inv_valid,
  input  wire          io_inputs_1_inv_ready,
  output wire          io_inputs_1_inv_payload_all,
  output wire [31:0]   io_inputs_1_inv_payload_address,
  output wire [5:0]    io_inputs_1_inv_payload_length,
  input  wire          io_inputs_1_ack_valid,
  output wire          io_inputs_1_ack_ready,
  output wire          io_inputs_1_sync_valid,
  input  wire          io_inputs_1_sync_ready,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire          io_output_cmd_payload_fragment_exclusive,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output wire [63:0]   io_output_cmd_payload_fragment_data,
  output wire [7:0]    io_output_cmd_payload_fragment_mask,
  output wire [3:0]    io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire          io_output_rsp_payload_fragment_exclusive,
  input  wire [63:0]   io_output_rsp_payload_fragment_data,
  input  wire [3:0]    io_output_rsp_payload_fragment_context,
  input  wire          io_output_inv_valid,
  output wire          io_output_inv_ready,
  input  wire          io_output_inv_payload_all,
  input  wire [31:0]   io_output_inv_payload_address,
  input  wire [5:0]    io_output_inv_payload_length,
  input  wire [0:0]    io_output_inv_payload_source,
  output wire          io_output_ack_valid,
  input  wire          io_output_ack_ready,
  input  wire          io_output_sync_valid,
  output wire          io_output_sync_ready,
  input  wire [0:0]    io_output_sync_payload_source,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire                streamFork_3_io_input_valid;
  wire                memory_arbiter_io_inputs_0_ready;
  wire                memory_arbiter_io_inputs_1_ready;
  wire                memory_arbiter_io_output_valid;
  wire                memory_arbiter_io_output_payload_last;
  wire       [0:0]    memory_arbiter_io_output_payload_fragment_source;
  wire       [0:0]    memory_arbiter_io_output_payload_fragment_opcode;
  wire                memory_arbiter_io_output_payload_fragment_exclusive;
  wire       [31:0]   memory_arbiter_io_output_payload_fragment_address;
  wire       [5:0]    memory_arbiter_io_output_payload_fragment_length;
  wire       [63:0]   memory_arbiter_io_output_payload_fragment_data;
  wire       [7:0]    memory_arbiter_io_output_payload_fragment_mask;
  wire       [3:0]    memory_arbiter_io_output_payload_fragment_context;
  wire       [0:0]    memory_arbiter_io_chosen;
  wire       [1:0]    memory_arbiter_io_chosenOH;
  wire                streamFork_3_io_input_ready;
  wire                streamFork_3_io_outputs_0_valid;
  wire                streamFork_3_io_outputs_0_payload_all;
  wire       [31:0]   streamFork_3_io_outputs_0_payload_address;
  wire       [5:0]    streamFork_3_io_outputs_0_payload_length;
  wire       [0:0]    streamFork_3_io_outputs_0_payload_source;
  wire                streamFork_3_io_outputs_1_valid;
  wire                streamFork_3_io_outputs_1_payload_all;
  wire       [31:0]   streamFork_3_io_outputs_1_payload_address;
  wire       [5:0]    streamFork_3_io_outputs_1_payload_length;
  wire       [0:0]    streamFork_3_io_outputs_1_payload_source;
  wire       [1:0]    _zz_io_output_cmd_payload_fragment_source;
  reg                 _zz_io_output_rsp_ready;
  reg                 _zz_io_output_sync_ready;
  wire       [0:0]    memory_rspSel;
  wire                io_output_inv_fire;
  wire                io_output_ack_fire;
  reg                 invalidate_invCounter_incrementIt;
  reg                 invalidate_invCounter_decrementIt;
  wire       [4:0]    invalidate_invCounter_valueNext;
  reg        [4:0]    invalidate_invCounter_value;
  wire                invalidate_invCounter_mayOverflow;
  wire                invalidate_invCounter_willOverflowIfInc;
  wire                invalidate_invCounter_willOverflow;
  reg        [4:0]    invalidate_invCounter_finalIncrement;
  wire                when_Utils_l735;
  wire                when_Utils_l737;
  wire                invalidate_haltInv;
  wire                _zz_io_output_inv_ready;
  wire                io_inputs_0_ack_fire;
  reg                 invalidate_logics_0_ackCounter_incrementIt;
  reg                 invalidate_logics_0_ackCounter_decrementIt;
  wire       [4:0]    invalidate_logics_0_ackCounter_valueNext;
  reg        [4:0]    invalidate_logics_0_ackCounter_value;
  wire                invalidate_logics_0_ackCounter_mayOverflow;
  wire                invalidate_logics_0_ackCounter_willOverflowIfInc;
  wire                invalidate_logics_0_ackCounter_willOverflow;
  reg        [4:0]    invalidate_logics_0_ackCounter_finalIncrement;
  wire                when_Utils_l735_1;
  wire                when_Utils_l737_1;
  wire                io_inputs_1_ack_fire;
  reg                 invalidate_logics_1_ackCounter_incrementIt;
  reg                 invalidate_logics_1_ackCounter_decrementIt;
  wire       [4:0]    invalidate_logics_1_ackCounter_valueNext;
  reg        [4:0]    invalidate_logics_1_ackCounter_value;
  wire                invalidate_logics_1_ackCounter_mayOverflow;
  wire                invalidate_logics_1_ackCounter_willOverflowIfInc;
  wire                invalidate_logics_1_ackCounter_willOverflow;
  reg        [4:0]    invalidate_logics_1_ackCounter_finalIncrement;
  wire                when_Utils_l735_2;
  wire                when_Utils_l737_2;
  wire       [0:0]    sync_syncSel;

  assign _zz_io_output_cmd_payload_fragment_source = {memory_arbiter_io_output_payload_fragment_source,memory_arbiter_io_chosen};
  StreamArbiter_5 memory_arbiter (
    .io_inputs_0_valid                      (io_inputs_0_cmd_valid                                  ), //i
    .io_inputs_0_ready                      (memory_arbiter_io_inputs_0_ready                       ), //o
    .io_inputs_0_payload_last               (io_inputs_0_cmd_payload_last                           ), //i
    .io_inputs_0_payload_fragment_source    (1'b0                                                   ), //i
    .io_inputs_0_payload_fragment_opcode    (io_inputs_0_cmd_payload_fragment_opcode                ), //i
    .io_inputs_0_payload_fragment_exclusive (io_inputs_0_cmd_payload_fragment_exclusive             ), //i
    .io_inputs_0_payload_fragment_address   (io_inputs_0_cmd_payload_fragment_address[31:0]         ), //i
    .io_inputs_0_payload_fragment_length    (io_inputs_0_cmd_payload_fragment_length[5:0]           ), //i
    .io_inputs_0_payload_fragment_data      (io_inputs_0_cmd_payload_fragment_data[63:0]            ), //i
    .io_inputs_0_payload_fragment_mask      (io_inputs_0_cmd_payload_fragment_mask[7:0]             ), //i
    .io_inputs_0_payload_fragment_context   (io_inputs_0_cmd_payload_fragment_context[3:0]          ), //i
    .io_inputs_1_valid                      (io_inputs_1_cmd_valid                                  ), //i
    .io_inputs_1_ready                      (memory_arbiter_io_inputs_1_ready                       ), //o
    .io_inputs_1_payload_last               (io_inputs_1_cmd_payload_last                           ), //i
    .io_inputs_1_payload_fragment_source    (1'b0                                                   ), //i
    .io_inputs_1_payload_fragment_opcode    (io_inputs_1_cmd_payload_fragment_opcode                ), //i
    .io_inputs_1_payload_fragment_exclusive (io_inputs_1_cmd_payload_fragment_exclusive             ), //i
    .io_inputs_1_payload_fragment_address   (io_inputs_1_cmd_payload_fragment_address[31:0]         ), //i
    .io_inputs_1_payload_fragment_length    (io_inputs_1_cmd_payload_fragment_length[5:0]           ), //i
    .io_inputs_1_payload_fragment_data      (io_inputs_1_cmd_payload_fragment_data[63:0]            ), //i
    .io_inputs_1_payload_fragment_mask      (io_inputs_1_cmd_payload_fragment_mask[7:0]             ), //i
    .io_inputs_1_payload_fragment_context   (io_inputs_1_cmd_payload_fragment_context[3:0]          ), //i
    .io_output_valid                        (memory_arbiter_io_output_valid                         ), //o
    .io_output_ready                        (io_output_cmd_ready                                    ), //i
    .io_output_payload_last                 (memory_arbiter_io_output_payload_last                  ), //o
    .io_output_payload_fragment_source      (memory_arbiter_io_output_payload_fragment_source       ), //o
    .io_output_payload_fragment_opcode      (memory_arbiter_io_output_payload_fragment_opcode       ), //o
    .io_output_payload_fragment_exclusive   (memory_arbiter_io_output_payload_fragment_exclusive    ), //o
    .io_output_payload_fragment_address     (memory_arbiter_io_output_payload_fragment_address[31:0]), //o
    .io_output_payload_fragment_length      (memory_arbiter_io_output_payload_fragment_length[5:0]  ), //o
    .io_output_payload_fragment_data        (memory_arbiter_io_output_payload_fragment_data[63:0]   ), //o
    .io_output_payload_fragment_mask        (memory_arbiter_io_output_payload_fragment_mask[7:0]    ), //o
    .io_output_payload_fragment_context     (memory_arbiter_io_output_payload_fragment_context[3:0] ), //o
    .io_chosen                              (memory_arbiter_io_chosen                               ), //o
    .io_chosenOH                            (memory_arbiter_io_chosenOH[1:0]                        ), //o
    .io_systemClk                           (io_systemClk                                           ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                             )  //i
  );
  StreamFork_2 streamFork_3 (
    .io_input_valid               (streamFork_3_io_input_valid                    ), //i
    .io_input_ready               (streamFork_3_io_input_ready                    ), //o
    .io_input_payload_all         (io_output_inv_payload_all                      ), //i
    .io_input_payload_address     (io_output_inv_payload_address[31:0]            ), //i
    .io_input_payload_length      (io_output_inv_payload_length[5:0]              ), //i
    .io_input_payload_source      (io_output_inv_payload_source                   ), //i
    .io_outputs_0_valid           (streamFork_3_io_outputs_0_valid                ), //o
    .io_outputs_0_ready           (io_inputs_0_inv_ready                          ), //i
    .io_outputs_0_payload_all     (streamFork_3_io_outputs_0_payload_all          ), //o
    .io_outputs_0_payload_address (streamFork_3_io_outputs_0_payload_address[31:0]), //o
    .io_outputs_0_payload_length  (streamFork_3_io_outputs_0_payload_length[5:0]  ), //o
    .io_outputs_0_payload_source  (streamFork_3_io_outputs_0_payload_source       ), //o
    .io_outputs_1_valid           (streamFork_3_io_outputs_1_valid                ), //o
    .io_outputs_1_ready           (io_inputs_1_inv_ready                          ), //i
    .io_outputs_1_payload_all     (streamFork_3_io_outputs_1_payload_all          ), //o
    .io_outputs_1_payload_address (streamFork_3_io_outputs_1_payload_address[31:0]), //o
    .io_outputs_1_payload_length  (streamFork_3_io_outputs_1_payload_length[5:0]  ), //o
    .io_outputs_1_payload_source  (streamFork_3_io_outputs_1_payload_source       ), //o
    .io_systemClk                 (io_systemClk                                   ), //i
    .systemCd_logic_outputReset   (systemCd_logic_outputReset                     )  //i
  );
  always @(*) begin
    case(memory_rspSel)
      1'b0 : _zz_io_output_rsp_ready = io_inputs_0_rsp_ready;
      default : _zz_io_output_rsp_ready = io_inputs_1_rsp_ready;
    endcase
  end

  always @(*) begin
    case(sync_syncSel)
      1'b0 : _zz_io_output_sync_ready = io_inputs_0_sync_ready;
      default : _zz_io_output_sync_ready = io_inputs_1_sync_ready;
    endcase
  end

  assign io_inputs_0_cmd_ready = memory_arbiter_io_inputs_0_ready;
  assign io_inputs_1_cmd_ready = memory_arbiter_io_inputs_1_ready;
  assign io_output_cmd_valid = memory_arbiter_io_output_valid;
  assign io_output_cmd_payload_last = memory_arbiter_io_output_payload_last;
  assign io_output_cmd_payload_fragment_opcode = memory_arbiter_io_output_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_exclusive = memory_arbiter_io_output_payload_fragment_exclusive;
  assign io_output_cmd_payload_fragment_address = memory_arbiter_io_output_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = memory_arbiter_io_output_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = memory_arbiter_io_output_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = memory_arbiter_io_output_payload_fragment_mask;
  assign io_output_cmd_payload_fragment_context = memory_arbiter_io_output_payload_fragment_context;
  assign io_output_cmd_payload_fragment_source = _zz_io_output_cmd_payload_fragment_source[0:0];
  assign memory_rspSel = io_output_rsp_payload_fragment_source[0 : 0];
  assign io_inputs_0_rsp_valid = (io_output_rsp_valid && (memory_rspSel == 1'b0));
  assign io_inputs_0_rsp_payload_last = io_output_rsp_payload_last;
  assign io_inputs_0_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_inputs_0_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_inputs_0_rsp_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign io_inputs_0_rsp_payload_fragment_exclusive = io_output_rsp_payload_fragment_exclusive;
  assign io_inputs_1_rsp_valid = (io_output_rsp_valid && (memory_rspSel == 1'b1));
  assign io_inputs_1_rsp_payload_last = io_output_rsp_payload_last;
  assign io_inputs_1_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_inputs_1_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_inputs_1_rsp_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign io_inputs_1_rsp_payload_fragment_exclusive = io_output_rsp_payload_fragment_exclusive;
  assign io_output_rsp_ready = _zz_io_output_rsp_ready;
  assign io_output_inv_fire = (io_output_inv_valid && io_output_inv_ready);
  assign io_output_ack_fire = (io_output_ack_valid && io_output_ack_ready);
  always @(*) begin
    invalidate_invCounter_incrementIt = 1'b0;
    if(io_output_inv_fire) begin
      invalidate_invCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    invalidate_invCounter_decrementIt = 1'b0;
    if(io_output_ack_fire) begin
      invalidate_invCounter_decrementIt = 1'b1;
    end
  end

  assign invalidate_invCounter_mayOverflow = (invalidate_invCounter_value == 5'h1f);
  assign invalidate_invCounter_willOverflowIfInc = (invalidate_invCounter_mayOverflow && (! invalidate_invCounter_decrementIt));
  assign invalidate_invCounter_willOverflow = (invalidate_invCounter_willOverflowIfInc && invalidate_invCounter_incrementIt);
  assign when_Utils_l735 = (invalidate_invCounter_incrementIt && (! invalidate_invCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l735) begin
      invalidate_invCounter_finalIncrement = 5'h01;
    end else begin
      if(when_Utils_l737) begin
        invalidate_invCounter_finalIncrement = 5'h1f;
      end else begin
        invalidate_invCounter_finalIncrement = 5'h0;
      end
    end
  end

  assign when_Utils_l737 = ((! invalidate_invCounter_incrementIt) && invalidate_invCounter_decrementIt);
  assign invalidate_invCounter_valueNext = (invalidate_invCounter_value + invalidate_invCounter_finalIncrement);
  assign invalidate_haltInv = invalidate_invCounter_value[4];
  assign _zz_io_output_inv_ready = (! invalidate_haltInv);
  assign io_output_inv_ready = (streamFork_3_io_input_ready && _zz_io_output_inv_ready);
  assign streamFork_3_io_input_valid = (io_output_inv_valid && _zz_io_output_inv_ready);
  assign io_inputs_0_ack_fire = (io_inputs_0_ack_valid && io_inputs_0_ack_ready);
  always @(*) begin
    invalidate_logics_0_ackCounter_incrementIt = 1'b0;
    if(io_inputs_0_ack_fire) begin
      invalidate_logics_0_ackCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    invalidate_logics_0_ackCounter_decrementIt = 1'b0;
    if(io_output_ack_fire) begin
      invalidate_logics_0_ackCounter_decrementIt = 1'b1;
    end
  end

  assign invalidate_logics_0_ackCounter_mayOverflow = (invalidate_logics_0_ackCounter_value == 5'h1f);
  assign invalidate_logics_0_ackCounter_willOverflowIfInc = (invalidate_logics_0_ackCounter_mayOverflow && (! invalidate_logics_0_ackCounter_decrementIt));
  assign invalidate_logics_0_ackCounter_willOverflow = (invalidate_logics_0_ackCounter_willOverflowIfInc && invalidate_logics_0_ackCounter_incrementIt);
  assign when_Utils_l735_1 = (invalidate_logics_0_ackCounter_incrementIt && (! invalidate_logics_0_ackCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_1) begin
      invalidate_logics_0_ackCounter_finalIncrement = 5'h01;
    end else begin
      if(when_Utils_l737_1) begin
        invalidate_logics_0_ackCounter_finalIncrement = 5'h1f;
      end else begin
        invalidate_logics_0_ackCounter_finalIncrement = 5'h0;
      end
    end
  end

  assign when_Utils_l737_1 = ((! invalidate_logics_0_ackCounter_incrementIt) && invalidate_logics_0_ackCounter_decrementIt);
  assign invalidate_logics_0_ackCounter_valueNext = (invalidate_logics_0_ackCounter_value + invalidate_logics_0_ackCounter_finalIncrement);
  assign io_inputs_0_inv_valid = streamFork_3_io_outputs_0_valid;
  assign io_inputs_0_inv_payload_address = streamFork_3_io_outputs_0_payload_address;
  assign io_inputs_0_inv_payload_length = streamFork_3_io_outputs_0_payload_length;
  assign io_inputs_0_inv_payload_all = (io_output_inv_payload_all || (io_output_inv_payload_source[0 : 0] != 1'b0));
  assign io_inputs_0_ack_ready = 1'b1;
  assign io_inputs_1_ack_fire = (io_inputs_1_ack_valid && io_inputs_1_ack_ready);
  always @(*) begin
    invalidate_logics_1_ackCounter_incrementIt = 1'b0;
    if(io_inputs_1_ack_fire) begin
      invalidate_logics_1_ackCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    invalidate_logics_1_ackCounter_decrementIt = 1'b0;
    if(io_output_ack_fire) begin
      invalidate_logics_1_ackCounter_decrementIt = 1'b1;
    end
  end

  assign invalidate_logics_1_ackCounter_mayOverflow = (invalidate_logics_1_ackCounter_value == 5'h1f);
  assign invalidate_logics_1_ackCounter_willOverflowIfInc = (invalidate_logics_1_ackCounter_mayOverflow && (! invalidate_logics_1_ackCounter_decrementIt));
  assign invalidate_logics_1_ackCounter_willOverflow = (invalidate_logics_1_ackCounter_willOverflowIfInc && invalidate_logics_1_ackCounter_incrementIt);
  assign when_Utils_l735_2 = (invalidate_logics_1_ackCounter_incrementIt && (! invalidate_logics_1_ackCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_2) begin
      invalidate_logics_1_ackCounter_finalIncrement = 5'h01;
    end else begin
      if(when_Utils_l737_2) begin
        invalidate_logics_1_ackCounter_finalIncrement = 5'h1f;
      end else begin
        invalidate_logics_1_ackCounter_finalIncrement = 5'h0;
      end
    end
  end

  assign when_Utils_l737_2 = ((! invalidate_logics_1_ackCounter_incrementIt) && invalidate_logics_1_ackCounter_decrementIt);
  assign invalidate_logics_1_ackCounter_valueNext = (invalidate_logics_1_ackCounter_value + invalidate_logics_1_ackCounter_finalIncrement);
  assign io_inputs_1_inv_valid = streamFork_3_io_outputs_1_valid;
  assign io_inputs_1_inv_payload_address = streamFork_3_io_outputs_1_payload_address;
  assign io_inputs_1_inv_payload_length = streamFork_3_io_outputs_1_payload_length;
  assign io_inputs_1_inv_payload_all = (io_output_inv_payload_all || (io_output_inv_payload_source[0 : 0] != 1'b1));
  assign io_inputs_1_ack_ready = 1'b1;
  assign io_output_ack_valid = (&{(invalidate_logics_1_ackCounter_value != 5'h0),(invalidate_logics_0_ackCounter_value != 5'h0)});
  assign sync_syncSel = io_output_sync_payload_source[0 : 0];
  assign io_inputs_0_sync_valid = (io_output_sync_valid && (sync_syncSel == 1'b0));
  assign io_inputs_1_sync_valid = (io_output_sync_valid && (sync_syncSel == 1'b1));
  assign io_output_sync_ready = _zz_io_output_sync_ready;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      invalidate_invCounter_value <= 5'h0;
      invalidate_logics_0_ackCounter_value <= 5'h0;
      invalidate_logics_1_ackCounter_value <= 5'h0;
    end else begin
      invalidate_invCounter_value <= invalidate_invCounter_valueNext;
      invalidate_logics_0_ackCounter_value <= invalidate_logics_0_ackCounter_valueNext;
      invalidate_logics_1_ackCounter_value <= invalidate_logics_1_ackCounter_valueNext;
    end
  end


endmodule

module BmbExclusiveMonitor (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire          io_input_cmd_payload_fragment_exclusive,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [63:0]   io_input_cmd_payload_fragment_data,
  input  wire [7:0]    io_input_cmd_payload_fragment_mask,
  input  wire [3:0]    io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire          io_input_rsp_payload_fragment_exclusive,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire [3:0]    io_input_rsp_payload_fragment_context,
  output wire          io_input_inv_valid,
  input  wire          io_input_inv_ready,
  output wire          io_input_inv_payload_all,
  output wire [31:0]   io_input_inv_payload_address,
  output wire [5:0]    io_input_inv_payload_length,
  output wire [0:0]    io_input_inv_payload_source,
  input  wire          io_input_ack_valid,
  output wire          io_input_ack_ready,
  output wire          io_input_sync_valid,
  input  wire          io_input_sync_ready,
  output wire [0:0]    io_input_sync_payload_source,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output wire [63:0]   io_output_cmd_payload_fragment_data,
  output reg  [7:0]    io_output_cmd_payload_fragment_mask,
  output wire [4:0]    io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_output_rsp_payload_fragment_data,
  input  wire [4:0]    io_output_rsp_payload_fragment_context,
  input  wire          io_output_inv_valid,
  output wire          io_output_inv_ready,
  input  wire          io_output_inv_payload_all,
  input  wire [31:0]   io_output_inv_payload_address,
  input  wire [5:0]    io_output_inv_payload_length,
  input  wire [0:0]    io_output_inv_payload_source,
  output wire          io_output_ack_valid,
  input  wire          io_output_ack_ready,
  input  wire          io_output_sync_valid,
  output wire          io_output_sync_ready,
  input  wire [0:0]    io_output_sync_payload_source,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);
  localparam BmbExclusiveMonitorState_IDLE = 2'd0;
  localparam BmbExclusiveMonitorState_FENCE_START = 2'd1;
  localparam BmbExclusiveMonitorState_FENCE_BUSY = 2'd2;
  localparam BmbExclusiveMonitorState_EMIT = 2'd3;

  wire                logic_cmdArbiter_io_output_ready;
  wire                logic_exclusiveReadArbiter_io_inputs_0_ready;
  wire                logic_exclusiveReadArbiter_io_inputs_1_ready;
  wire                logic_exclusiveReadArbiter_io_output_valid;
  wire                logic_exclusiveReadArbiter_io_output_payload_last;
  wire       [0:0]    logic_exclusiveReadArbiter_io_output_payload_fragment_source;
  wire       [0:0]    logic_exclusiveReadArbiter_io_output_payload_fragment_opcode;
  wire                logic_exclusiveReadArbiter_io_output_payload_fragment_exclusive;
  wire       [31:0]   logic_exclusiveReadArbiter_io_output_payload_fragment_address;
  wire       [5:0]    logic_exclusiveReadArbiter_io_output_payload_fragment_length;
  wire       [3:0]    logic_exclusiveReadArbiter_io_output_payload_fragment_context;
  wire       [0:0]    logic_exclusiveReadArbiter_io_chosen;
  wire       [1:0]    logic_exclusiveReadArbiter_io_chosenOH;
  wire                logic_cmdArbiter_io_inputs_0_ready;
  wire                logic_cmdArbiter_io_inputs_1_ready;
  wire                logic_cmdArbiter_io_output_valid;
  wire                logic_cmdArbiter_io_output_payload_last;
  wire       [0:0]    logic_cmdArbiter_io_output_payload_fragment_source;
  wire       [0:0]    logic_cmdArbiter_io_output_payload_fragment_opcode;
  wire                logic_cmdArbiter_io_output_payload_fragment_exclusive;
  wire       [31:0]   logic_cmdArbiter_io_output_payload_fragment_address;
  wire       [5:0]    logic_cmdArbiter_io_output_payload_fragment_length;
  wire       [3:0]    logic_cmdArbiter_io_output_payload_fragment_context;
  wire       [0:0]    logic_cmdArbiter_io_chosen;
  wire       [1:0]    logic_cmdArbiter_io_chosenOH;
  wire       [11:0]   _zz_logic_inputAddressLowEnd;
  wire       [19:0]   _zz_logic_sources_0_addressHitHigh;
  wire       [19:0]   _zz_logic_sources_0_addressHitHigh_1;
  wire       [19:0]   _zz_logic_sources_1_addressHitHigh;
  wire       [19:0]   _zz_logic_sources_1_addressHitHigh_1;
  reg                 logic_fence_start;
  reg                 logic_fence_done;
  reg                 logic_fence_busy;
  reg                 logic_exclusiveWriteCancel;
  wire       [11:0]   logic_inputAddressLow;
  wire       [11:0]   logic_inputAddressLowEnd;
  reg                 logic_sources_0_valid;
  reg                 logic_sources_0_exclusiveWritePending;
  reg        [1:0]    logic_sources_0_state;
  reg        [31:0]   logic_sources_0_address;
  reg        [5:0]    logic_sources_0_length;
  reg        [3:0]    logic_sources_0_context;
  wire       [11:0]   logic_sources_0_addressLow;
  reg        [11:0]   logic_sources_0_addressLowEnd;
  wire                logic_sources_0_addressHitHigh;
  wire                logic_sources_0_addressHitLow;
  wire                logic_sources_0_addressHit;
  wire                logic_sources_0_inputSourceHit;
  wire                logic_sources_0_haltSource;
  wire                io_output_rsp_fire;
  wire                when_BmbExclusiveMonitor_l65;
  wire                when_BmbExclusiveMonitor_l69;
  wire                when_BmbExclusiveMonitor_l70;
  wire                io_input_cmd_fire;
  wire                when_BmbExclusiveMonitor_l79;
  wire                when_BmbExclusiveMonitor_l80;
  reg                 logic_sources_0_exclusiveReadCmd_valid;
  wire                logic_sources_0_exclusiveReadCmd_ready;
  wire                logic_sources_0_exclusiveReadCmd_payload_last;
  wire       [0:0]    logic_sources_0_exclusiveReadCmd_payload_fragment_source;
  wire       [0:0]    logic_sources_0_exclusiveReadCmd_payload_fragment_opcode;
  wire                logic_sources_0_exclusiveReadCmd_payload_fragment_exclusive;
  wire       [31:0]   logic_sources_0_exclusiveReadCmd_payload_fragment_address;
  wire       [5:0]    logic_sources_0_exclusiveReadCmd_payload_fragment_length;
  wire       [3:0]    logic_sources_0_exclusiveReadCmd_payload_fragment_context;
  wire                when_BmbExclusiveMonitor_l101;
  reg                 logic_sources_1_valid;
  reg                 logic_sources_1_exclusiveWritePending;
  reg        [1:0]    logic_sources_1_state;
  reg        [31:0]   logic_sources_1_address;
  reg        [5:0]    logic_sources_1_length;
  reg        [3:0]    logic_sources_1_context;
  wire       [11:0]   logic_sources_1_addressLow;
  reg        [11:0]   logic_sources_1_addressLowEnd;
  wire                logic_sources_1_addressHitHigh;
  wire                logic_sources_1_addressHitLow;
  wire                logic_sources_1_addressHit;
  wire                logic_sources_1_inputSourceHit;
  wire                logic_sources_1_haltSource;
  wire                when_BmbExclusiveMonitor_l65_1;
  wire                when_BmbExclusiveMonitor_l69_1;
  wire                when_BmbExclusiveMonitor_l70_1;
  wire                when_BmbExclusiveMonitor_l79_1;
  wire                when_BmbExclusiveMonitor_l80_1;
  reg                 logic_sources_1_exclusiveReadCmd_valid;
  wire                logic_sources_1_exclusiveReadCmd_ready;
  wire                logic_sources_1_exclusiveReadCmd_payload_last;
  wire       [0:0]    logic_sources_1_exclusiveReadCmd_payload_fragment_source;
  wire       [0:0]    logic_sources_1_exclusiveReadCmd_payload_fragment_opcode;
  wire                logic_sources_1_exclusiveReadCmd_payload_fragment_exclusive;
  wire       [31:0]   logic_sources_1_exclusiveReadCmd_payload_fragment_address;
  wire       [5:0]    logic_sources_1_exclusiveReadCmd_payload_fragment_length;
  wire       [3:0]    logic_sources_1_exclusiveReadCmd_payload_fragment_context;
  wire                when_BmbExclusiveMonitor_l101_1;
  reg        [6:0]    logic_trackers_0_cmdCounter;
  reg        [6:0]    logic_trackers_0_rspCounter;
  wire                logic_trackers_0_full;
  wire                io_output_cmd_fire;
  reg                 io_output_cmd_payload_first;
  wire                when_BmbExclusiveMonitor_l123;
  reg                 io_output_rsp_payload_first;
  wire                when_BmbExclusiveMonitor_l126;
  reg        [6:0]    logic_trackers_0_target;
  wire                logic_trackers_0_hit;
  reg                 logic_trackers_0_done;
  wire                when_BmbExclusiveMonitor_l141;
  reg        [6:0]    logic_trackers_1_cmdCounter;
  reg        [6:0]    logic_trackers_1_rspCounter;
  wire                logic_trackers_1_full;
  wire                when_BmbExclusiveMonitor_l123_1;
  wire                when_BmbExclusiveMonitor_l126_1;
  reg        [6:0]    logic_trackers_1_target;
  wire                logic_trackers_1_hit;
  reg                 logic_trackers_1_done;
  wire                when_BmbExclusiveMonitor_l141_1;
  wire                _zz_io_input_cmd_ready;
  reg                 _zz_io_input_cmd_ready_1;
  wire                when_Stream_l445;
  reg                 logic_inputCmdHalted_valid;
  wire                logic_inputCmdHalted_ready;
  wire                logic_inputCmdHalted_payload_last;
  wire       [0:0]    logic_inputCmdHalted_payload_fragment_source;
  wire       [0:0]    logic_inputCmdHalted_payload_fragment_opcode;
  wire                logic_inputCmdHalted_payload_fragment_exclusive;
  wire       [31:0]   logic_inputCmdHalted_payload_fragment_address;
  wire       [5:0]    logic_inputCmdHalted_payload_fragment_length;
  wire       [63:0]   logic_inputCmdHalted_payload_fragment_data;
  wire       [7:0]    logic_inputCmdHalted_payload_fragment_mask;
  wire       [3:0]    logic_inputCmdHalted_payload_fragment_context;
  wire                logic_exclusiveSuccess;
  wire                _zz_io_output_cmd_valid;
  wire                when_BmbExclusiveMonitor_l163;
  `ifndef SYNTHESIS
  reg [87:0] logic_sources_0_state_string;
  reg [87:0] logic_sources_1_state_string;
  `endif


  assign _zz_logic_inputAddressLowEnd = {6'd0, io_input_cmd_payload_fragment_length};
  assign _zz_logic_sources_0_addressHitHigh = (logic_sources_0_address >>> 4'd12);
  assign _zz_logic_sources_0_addressHitHigh_1 = (io_input_cmd_payload_fragment_address >>> 4'd12);
  assign _zz_logic_sources_1_addressHitHigh = (logic_sources_1_address >>> 4'd12);
  assign _zz_logic_sources_1_addressHitHigh_1 = (io_input_cmd_payload_fragment_address >>> 4'd12);
  StreamArbiter_3 logic_exclusiveReadArbiter (
    .io_inputs_0_valid                      (logic_sources_0_exclusiveReadCmd_valid                             ), //i
    .io_inputs_0_ready                      (logic_exclusiveReadArbiter_io_inputs_0_ready                       ), //o
    .io_inputs_0_payload_last               (logic_sources_0_exclusiveReadCmd_payload_last                      ), //i
    .io_inputs_0_payload_fragment_source    (logic_sources_0_exclusiveReadCmd_payload_fragment_source           ), //i
    .io_inputs_0_payload_fragment_opcode    (logic_sources_0_exclusiveReadCmd_payload_fragment_opcode           ), //i
    .io_inputs_0_payload_fragment_exclusive (logic_sources_0_exclusiveReadCmd_payload_fragment_exclusive        ), //i
    .io_inputs_0_payload_fragment_address   (logic_sources_0_exclusiveReadCmd_payload_fragment_address[31:0]    ), //i
    .io_inputs_0_payload_fragment_length    (logic_sources_0_exclusiveReadCmd_payload_fragment_length[5:0]      ), //i
    .io_inputs_0_payload_fragment_context   (logic_sources_0_exclusiveReadCmd_payload_fragment_context[3:0]     ), //i
    .io_inputs_1_valid                      (logic_sources_1_exclusiveReadCmd_valid                             ), //i
    .io_inputs_1_ready                      (logic_exclusiveReadArbiter_io_inputs_1_ready                       ), //o
    .io_inputs_1_payload_last               (logic_sources_1_exclusiveReadCmd_payload_last                      ), //i
    .io_inputs_1_payload_fragment_source    (logic_sources_1_exclusiveReadCmd_payload_fragment_source           ), //i
    .io_inputs_1_payload_fragment_opcode    (logic_sources_1_exclusiveReadCmd_payload_fragment_opcode           ), //i
    .io_inputs_1_payload_fragment_exclusive (logic_sources_1_exclusiveReadCmd_payload_fragment_exclusive        ), //i
    .io_inputs_1_payload_fragment_address   (logic_sources_1_exclusiveReadCmd_payload_fragment_address[31:0]    ), //i
    .io_inputs_1_payload_fragment_length    (logic_sources_1_exclusiveReadCmd_payload_fragment_length[5:0]      ), //i
    .io_inputs_1_payload_fragment_context   (logic_sources_1_exclusiveReadCmd_payload_fragment_context[3:0]     ), //i
    .io_output_valid                        (logic_exclusiveReadArbiter_io_output_valid                         ), //o
    .io_output_ready                        (logic_cmdArbiter_io_inputs_0_ready                                 ), //i
    .io_output_payload_last                 (logic_exclusiveReadArbiter_io_output_payload_last                  ), //o
    .io_output_payload_fragment_source      (logic_exclusiveReadArbiter_io_output_payload_fragment_source       ), //o
    .io_output_payload_fragment_opcode      (logic_exclusiveReadArbiter_io_output_payload_fragment_opcode       ), //o
    .io_output_payload_fragment_exclusive   (logic_exclusiveReadArbiter_io_output_payload_fragment_exclusive    ), //o
    .io_output_payload_fragment_address     (logic_exclusiveReadArbiter_io_output_payload_fragment_address[31:0]), //o
    .io_output_payload_fragment_length      (logic_exclusiveReadArbiter_io_output_payload_fragment_length[5:0]  ), //o
    .io_output_payload_fragment_context     (logic_exclusiveReadArbiter_io_output_payload_fragment_context[3:0] ), //o
    .io_chosen                              (logic_exclusiveReadArbiter_io_chosen                               ), //o
    .io_chosenOH                            (logic_exclusiveReadArbiter_io_chosenOH[1:0]                        ), //o
    .io_systemClk                           (io_systemClk                                                       ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                         )  //i
  );
  StreamArbiter_4 logic_cmdArbiter (
    .io_inputs_0_valid                      (logic_exclusiveReadArbiter_io_output_valid                         ), //i
    .io_inputs_0_ready                      (logic_cmdArbiter_io_inputs_0_ready                                 ), //o
    .io_inputs_0_payload_last               (logic_exclusiveReadArbiter_io_output_payload_last                  ), //i
    .io_inputs_0_payload_fragment_source    (logic_exclusiveReadArbiter_io_output_payload_fragment_source       ), //i
    .io_inputs_0_payload_fragment_opcode    (logic_exclusiveReadArbiter_io_output_payload_fragment_opcode       ), //i
    .io_inputs_0_payload_fragment_exclusive (logic_exclusiveReadArbiter_io_output_payload_fragment_exclusive    ), //i
    .io_inputs_0_payload_fragment_address   (logic_exclusiveReadArbiter_io_output_payload_fragment_address[31:0]), //i
    .io_inputs_0_payload_fragment_length    (logic_exclusiveReadArbiter_io_output_payload_fragment_length[5:0]  ), //i
    .io_inputs_0_payload_fragment_context   (logic_exclusiveReadArbiter_io_output_payload_fragment_context[3:0] ), //i
    .io_inputs_1_valid                      (logic_inputCmdHalted_valid                                         ), //i
    .io_inputs_1_ready                      (logic_cmdArbiter_io_inputs_1_ready                                 ), //o
    .io_inputs_1_payload_last               (logic_inputCmdHalted_payload_last                                  ), //i
    .io_inputs_1_payload_fragment_source    (logic_inputCmdHalted_payload_fragment_source                       ), //i
    .io_inputs_1_payload_fragment_opcode    (logic_inputCmdHalted_payload_fragment_opcode                       ), //i
    .io_inputs_1_payload_fragment_exclusive (logic_inputCmdHalted_payload_fragment_exclusive                    ), //i
    .io_inputs_1_payload_fragment_address   (logic_inputCmdHalted_payload_fragment_address[31:0]                ), //i
    .io_inputs_1_payload_fragment_length    (logic_inputCmdHalted_payload_fragment_length[5:0]                  ), //i
    .io_inputs_1_payload_fragment_context   (logic_inputCmdHalted_payload_fragment_context[3:0]                 ), //i
    .io_output_valid                        (logic_cmdArbiter_io_output_valid                                   ), //o
    .io_output_ready                        (logic_cmdArbiter_io_output_ready                                   ), //i
    .io_output_payload_last                 (logic_cmdArbiter_io_output_payload_last                            ), //o
    .io_output_payload_fragment_source      (logic_cmdArbiter_io_output_payload_fragment_source                 ), //o
    .io_output_payload_fragment_opcode      (logic_cmdArbiter_io_output_payload_fragment_opcode                 ), //o
    .io_output_payload_fragment_exclusive   (logic_cmdArbiter_io_output_payload_fragment_exclusive              ), //o
    .io_output_payload_fragment_address     (logic_cmdArbiter_io_output_payload_fragment_address[31:0]          ), //o
    .io_output_payload_fragment_length      (logic_cmdArbiter_io_output_payload_fragment_length[5:0]            ), //o
    .io_output_payload_fragment_context     (logic_cmdArbiter_io_output_payload_fragment_context[3:0]           ), //o
    .io_chosen                              (logic_cmdArbiter_io_chosen                                         ), //o
    .io_chosenOH                            (logic_cmdArbiter_io_chosenOH[1:0]                                  ), //o
    .io_systemClk                           (io_systemClk                                                       ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                                         )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(logic_sources_0_state)
      BmbExclusiveMonitorState_IDLE : logic_sources_0_state_string = "IDLE       ";
      BmbExclusiveMonitorState_FENCE_START : logic_sources_0_state_string = "FENCE_START";
      BmbExclusiveMonitorState_FENCE_BUSY : logic_sources_0_state_string = "FENCE_BUSY ";
      BmbExclusiveMonitorState_EMIT : logic_sources_0_state_string = "EMIT       ";
      default : logic_sources_0_state_string = "???????????";
    endcase
  end
  always @(*) begin
    case(logic_sources_1_state)
      BmbExclusiveMonitorState_IDLE : logic_sources_1_state_string = "IDLE       ";
      BmbExclusiveMonitorState_FENCE_START : logic_sources_1_state_string = "FENCE_START";
      BmbExclusiveMonitorState_FENCE_BUSY : logic_sources_1_state_string = "FENCE_BUSY ";
      BmbExclusiveMonitorState_EMIT : logic_sources_1_state_string = "EMIT       ";
      default : logic_sources_1_state_string = "???????????";
    endcase
  end
  `endif

  always @(*) begin
    logic_fence_start = 1'b0;
    case(logic_sources_0_state)
      BmbExclusiveMonitorState_FENCE_START : begin
        if(when_BmbExclusiveMonitor_l101) begin
          logic_fence_start = 1'b1;
        end
      end
      default : begin
      end
    endcase
    case(logic_sources_1_state)
      BmbExclusiveMonitorState_FENCE_START : begin
        if(when_BmbExclusiveMonitor_l101_1) begin
          logic_fence_start = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    logic_fence_done = 1'b1;
    if(when_BmbExclusiveMonitor_l141) begin
      logic_fence_done = 1'b0;
    end
    if(when_BmbExclusiveMonitor_l141_1) begin
      logic_fence_done = 1'b0;
    end
  end

  always @(*) begin
    logic_exclusiveWriteCancel = 1'b0;
    if(when_BmbExclusiveMonitor_l163) begin
      logic_exclusiveWriteCancel = 1'b1;
    end
  end

  assign logic_inputAddressLow = io_input_cmd_payload_fragment_address[11 : 0];
  assign logic_inputAddressLowEnd = (logic_inputAddressLow + _zz_logic_inputAddressLowEnd);
  assign logic_sources_0_addressLow = logic_sources_0_address[11 : 0];
  assign logic_sources_0_addressHitHigh = (_zz_logic_sources_0_addressHitHigh == _zz_logic_sources_0_addressHitHigh_1);
  assign logic_sources_0_addressHitLow = ((logic_sources_0_addressLow <= logic_inputAddressLowEnd) && (logic_inputAddressLow <= logic_sources_0_addressLowEnd));
  assign logic_sources_0_addressHit = (logic_sources_0_addressHitLow && logic_sources_0_addressHitHigh);
  assign logic_sources_0_inputSourceHit = (io_input_cmd_payload_fragment_source == 1'b0);
  assign logic_sources_0_haltSource = (logic_sources_0_state != BmbExclusiveMonitorState_IDLE);
  assign io_output_rsp_fire = (io_output_rsp_valid && io_output_rsp_ready);
  assign when_BmbExclusiveMonitor_l65 = ((io_output_rsp_fire && (io_output_rsp_payload_fragment_source == 1'b0)) && io_output_rsp_payload_fragment_context[4]);
  assign when_BmbExclusiveMonitor_l69 = ((io_input_cmd_valid && (io_input_cmd_payload_fragment_opcode == 1'b0)) && io_input_cmd_payload_fragment_exclusive);
  assign when_BmbExclusiveMonitor_l70 = (logic_sources_0_inputSourceHit && (! logic_sources_0_haltSource));
  assign io_input_cmd_fire = (io_input_cmd_valid && io_input_cmd_ready);
  assign when_BmbExclusiveMonitor_l79 = ((logic_sources_0_addressHit && (io_input_cmd_fire && io_input_cmd_payload_last)) && (io_input_cmd_payload_fragment_opcode == 1'b1));
  assign when_BmbExclusiveMonitor_l80 = (! logic_exclusiveWriteCancel);
  always @(*) begin
    logic_sources_0_exclusiveReadCmd_valid = 1'b0;
    case(logic_sources_0_state)
      BmbExclusiveMonitorState_EMIT : begin
        logic_sources_0_exclusiveReadCmd_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign logic_sources_0_exclusiveReadCmd_payload_fragment_opcode = 1'b0;
  assign logic_sources_0_exclusiveReadCmd_payload_fragment_exclusive = 1'b1;
  assign logic_sources_0_exclusiveReadCmd_payload_fragment_address = logic_sources_0_address;
  assign logic_sources_0_exclusiveReadCmd_payload_fragment_length = logic_sources_0_length;
  assign logic_sources_0_exclusiveReadCmd_payload_fragment_context = logic_sources_0_context;
  assign logic_sources_0_exclusiveReadCmd_payload_fragment_source = 1'b0;
  assign logic_sources_0_exclusiveReadCmd_payload_last = 1'b1;
  assign when_BmbExclusiveMonitor_l101 = (! logic_fence_busy);
  assign logic_sources_1_addressLow = logic_sources_1_address[11 : 0];
  assign logic_sources_1_addressHitHigh = (_zz_logic_sources_1_addressHitHigh == _zz_logic_sources_1_addressHitHigh_1);
  assign logic_sources_1_addressHitLow = ((logic_sources_1_addressLow <= logic_inputAddressLowEnd) && (logic_inputAddressLow <= logic_sources_1_addressLowEnd));
  assign logic_sources_1_addressHit = (logic_sources_1_addressHitLow && logic_sources_1_addressHitHigh);
  assign logic_sources_1_inputSourceHit = (io_input_cmd_payload_fragment_source == 1'b1);
  assign logic_sources_1_haltSource = (logic_sources_1_state != BmbExclusiveMonitorState_IDLE);
  assign when_BmbExclusiveMonitor_l65_1 = ((io_output_rsp_fire && (io_output_rsp_payload_fragment_source == 1'b1)) && io_output_rsp_payload_fragment_context[4]);
  assign when_BmbExclusiveMonitor_l69_1 = ((io_input_cmd_valid && (io_input_cmd_payload_fragment_opcode == 1'b0)) && io_input_cmd_payload_fragment_exclusive);
  assign when_BmbExclusiveMonitor_l70_1 = (logic_sources_1_inputSourceHit && (! logic_sources_1_haltSource));
  assign when_BmbExclusiveMonitor_l79_1 = ((logic_sources_1_addressHit && (io_input_cmd_fire && io_input_cmd_payload_last)) && (io_input_cmd_payload_fragment_opcode == 1'b1));
  assign when_BmbExclusiveMonitor_l80_1 = (! logic_exclusiveWriteCancel);
  always @(*) begin
    logic_sources_1_exclusiveReadCmd_valid = 1'b0;
    case(logic_sources_1_state)
      BmbExclusiveMonitorState_EMIT : begin
        logic_sources_1_exclusiveReadCmd_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign logic_sources_1_exclusiveReadCmd_payload_fragment_opcode = 1'b0;
  assign logic_sources_1_exclusiveReadCmd_payload_fragment_exclusive = 1'b1;
  assign logic_sources_1_exclusiveReadCmd_payload_fragment_address = logic_sources_1_address;
  assign logic_sources_1_exclusiveReadCmd_payload_fragment_length = logic_sources_1_length;
  assign logic_sources_1_exclusiveReadCmd_payload_fragment_context = logic_sources_1_context;
  assign logic_sources_1_exclusiveReadCmd_payload_fragment_source = 1'b1;
  assign logic_sources_1_exclusiveReadCmd_payload_last = 1'b1;
  assign when_BmbExclusiveMonitor_l101_1 = (! logic_fence_busy);
  assign logic_trackers_0_full = ((logic_trackers_0_cmdCounter[6] != logic_trackers_0_rspCounter[6]) && (logic_trackers_0_cmdCounter[5 : 0] == logic_trackers_0_rspCounter[5 : 0]));
  assign io_output_cmd_fire = (io_output_cmd_valid && io_output_cmd_ready);
  assign when_BmbExclusiveMonitor_l123 = ((io_output_cmd_fire && io_output_cmd_payload_first) && (io_output_cmd_payload_fragment_source == 1'b0));
  assign when_BmbExclusiveMonitor_l126 = ((io_output_rsp_fire && io_output_rsp_payload_first) && (io_output_rsp_payload_fragment_source == 1'b0));
  assign logic_trackers_0_hit = (logic_trackers_0_target == logic_trackers_0_rspCounter);
  assign when_BmbExclusiveMonitor_l141 = (! logic_trackers_0_done);
  assign logic_trackers_1_full = ((logic_trackers_1_cmdCounter[6] != logic_trackers_1_rspCounter[6]) && (logic_trackers_1_cmdCounter[5 : 0] == logic_trackers_1_rspCounter[5 : 0]));
  assign when_BmbExclusiveMonitor_l123_1 = ((io_output_cmd_fire && io_output_cmd_payload_first) && (io_output_cmd_payload_fragment_source == 1'b1));
  assign when_BmbExclusiveMonitor_l126_1 = ((io_output_rsp_fire && io_output_rsp_payload_first) && (io_output_rsp_payload_fragment_source == 1'b1));
  assign logic_trackers_1_hit = (logic_trackers_1_target == logic_trackers_1_rspCounter);
  assign when_BmbExclusiveMonitor_l141_1 = (! logic_trackers_1_done);
  assign logic_sources_0_exclusiveReadCmd_ready = logic_exclusiveReadArbiter_io_inputs_0_ready;
  assign logic_sources_1_exclusiveReadCmd_ready = logic_exclusiveReadArbiter_io_inputs_1_ready;
  assign _zz_io_input_cmd_ready = (! (|{(logic_sources_1_inputSourceHit && logic_sources_1_haltSource),(logic_sources_0_inputSourceHit && logic_sources_0_haltSource)}));
  assign io_input_cmd_ready = (_zz_io_input_cmd_ready_1 && _zz_io_input_cmd_ready);
  assign when_Stream_l445 = ((io_input_cmd_valid && (io_input_cmd_payload_fragment_opcode == 1'b0)) && io_input_cmd_payload_fragment_exclusive);
  always @(*) begin
    logic_inputCmdHalted_valid = (io_input_cmd_valid && _zz_io_input_cmd_ready);
    if(when_Stream_l445) begin
      logic_inputCmdHalted_valid = 1'b0;
    end
  end

  always @(*) begin
    _zz_io_input_cmd_ready_1 = logic_inputCmdHalted_ready;
    if(when_Stream_l445) begin
      _zz_io_input_cmd_ready_1 = 1'b1;
    end
  end

  assign logic_inputCmdHalted_payload_last = io_input_cmd_payload_last;
  assign logic_inputCmdHalted_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign logic_inputCmdHalted_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign logic_inputCmdHalted_payload_fragment_exclusive = io_input_cmd_payload_fragment_exclusive;
  assign logic_inputCmdHalted_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign logic_inputCmdHalted_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign logic_inputCmdHalted_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign logic_inputCmdHalted_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign logic_inputCmdHalted_payload_fragment_context = io_input_cmd_payload_fragment_context;
  assign logic_inputCmdHalted_ready = logic_cmdArbiter_io_inputs_1_ready;
  assign logic_exclusiveSuccess = (|{((logic_sources_1_valid && logic_sources_1_addressHit) && logic_sources_1_inputSourceHit),((logic_sources_0_valid && logic_sources_0_addressHit) && logic_sources_0_inputSourceHit)});
  assign _zz_io_output_cmd_valid = (! (|{logic_trackers_1_full,logic_trackers_0_full}));
  assign logic_cmdArbiter_io_output_ready = (io_output_cmd_ready && _zz_io_output_cmd_valid);
  assign io_output_cmd_valid = (logic_cmdArbiter_io_output_valid && _zz_io_output_cmd_valid);
  assign io_output_cmd_payload_last = logic_cmdArbiter_io_output_payload_last;
  assign io_output_cmd_payload_fragment_source = logic_cmdArbiter_io_output_payload_fragment_source;
  assign io_output_cmd_payload_fragment_opcode = logic_cmdArbiter_io_output_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = logic_cmdArbiter_io_output_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = logic_cmdArbiter_io_output_payload_fragment_length;
  assign io_output_cmd_payload_fragment_context = {(io_input_cmd_payload_fragment_exclusive && logic_exclusiveSuccess),logic_cmdArbiter_io_output_payload_fragment_context};
  assign io_output_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  always @(*) begin
    io_output_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
    if(when_BmbExclusiveMonitor_l163) begin
      io_output_cmd_payload_fragment_mask = 8'h0;
    end
  end

  assign when_BmbExclusiveMonitor_l163 = (io_input_cmd_payload_fragment_exclusive && (! logic_exclusiveSuccess));
  assign io_input_rsp_valid = io_output_rsp_valid;
  assign io_output_rsp_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = io_output_rsp_payload_last;
  assign io_input_rsp_payload_fragment_source = io_output_rsp_payload_fragment_source;
  assign io_input_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = io_output_rsp_payload_fragment_context[3:0];
  assign io_input_rsp_payload_fragment_exclusive = io_output_rsp_payload_fragment_context[4];
  assign io_input_inv_valid = io_output_inv_valid;
  assign io_output_inv_ready = io_input_inv_ready;
  assign io_input_inv_payload_all = io_output_inv_payload_all;
  assign io_input_inv_payload_address = io_output_inv_payload_address;
  assign io_input_inv_payload_length = io_output_inv_payload_length;
  assign io_input_inv_payload_source = io_output_inv_payload_source;
  assign io_output_ack_valid = io_input_ack_valid;
  assign io_input_ack_ready = io_output_ack_ready;
  assign io_input_sync_valid = io_output_sync_valid;
  assign io_output_sync_ready = io_input_sync_ready;
  assign io_input_sync_payload_source = io_output_sync_payload_source;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      logic_fence_busy <= 1'b0;
      logic_sources_0_valid <= 1'b0;
      logic_sources_0_exclusiveWritePending <= 1'b0;
      logic_sources_0_state <= BmbExclusiveMonitorState_IDLE;
      logic_sources_1_valid <= 1'b0;
      logic_sources_1_exclusiveWritePending <= 1'b0;
      logic_sources_1_state <= BmbExclusiveMonitorState_IDLE;
      logic_trackers_0_cmdCounter <= 7'h0;
      logic_trackers_0_rspCounter <= 7'h0;
      io_output_cmd_payload_first <= 1'b1;
      io_output_rsp_payload_first <= 1'b1;
      logic_trackers_1_cmdCounter <= 7'h0;
      logic_trackers_1_rspCounter <= 7'h0;
    end else begin
      if(logic_fence_done) begin
        logic_fence_busy <= 1'b0;
      end
      if(logic_fence_start) begin
        logic_fence_busy <= 1'b1;
      end
      if(when_BmbExclusiveMonitor_l65) begin
        logic_sources_0_exclusiveWritePending <= 1'b0;
      end
      if(when_BmbExclusiveMonitor_l69) begin
        if(when_BmbExclusiveMonitor_l70) begin
          logic_sources_0_valid <= 1'b1;
          logic_sources_0_state <= BmbExclusiveMonitorState_FENCE_START;
        end
      end
      if(when_BmbExclusiveMonitor_l79) begin
        if(when_BmbExclusiveMonitor_l80) begin
          logic_sources_0_valid <= 1'b0;
        end
        if(logic_sources_0_inputSourceHit) begin
          logic_sources_0_exclusiveWritePending <= 1'b1;
        end
      end
      case(logic_sources_0_state)
        BmbExclusiveMonitorState_FENCE_START : begin
          if(when_BmbExclusiveMonitor_l101) begin
            logic_sources_0_state <= BmbExclusiveMonitorState_FENCE_BUSY;
          end
        end
        BmbExclusiveMonitorState_FENCE_BUSY : begin
          if(logic_fence_done) begin
            logic_sources_0_state <= BmbExclusiveMonitorState_EMIT;
          end
        end
        BmbExclusiveMonitorState_EMIT : begin
          if(logic_sources_0_exclusiveReadCmd_ready) begin
            logic_sources_0_state <= BmbExclusiveMonitorState_IDLE;
          end
        end
        default : begin
        end
      endcase
      if(when_BmbExclusiveMonitor_l65_1) begin
        logic_sources_1_exclusiveWritePending <= 1'b0;
      end
      if(when_BmbExclusiveMonitor_l69_1) begin
        if(when_BmbExclusiveMonitor_l70_1) begin
          logic_sources_1_valid <= 1'b1;
          logic_sources_1_state <= BmbExclusiveMonitorState_FENCE_START;
        end
      end
      if(when_BmbExclusiveMonitor_l79_1) begin
        if(when_BmbExclusiveMonitor_l80_1) begin
          logic_sources_1_valid <= 1'b0;
        end
        if(logic_sources_1_inputSourceHit) begin
          logic_sources_1_exclusiveWritePending <= 1'b1;
        end
      end
      case(logic_sources_1_state)
        BmbExclusiveMonitorState_FENCE_START : begin
          if(when_BmbExclusiveMonitor_l101_1) begin
            logic_sources_1_state <= BmbExclusiveMonitorState_FENCE_BUSY;
          end
        end
        BmbExclusiveMonitorState_FENCE_BUSY : begin
          if(logic_fence_done) begin
            logic_sources_1_state <= BmbExclusiveMonitorState_EMIT;
          end
        end
        BmbExclusiveMonitorState_EMIT : begin
          if(logic_sources_1_exclusiveReadCmd_ready) begin
            logic_sources_1_state <= BmbExclusiveMonitorState_IDLE;
          end
        end
        default : begin
        end
      endcase
      if(io_output_cmd_fire) begin
        io_output_cmd_payload_first <= io_output_cmd_payload_last;
      end
      if(when_BmbExclusiveMonitor_l123) begin
        logic_trackers_0_cmdCounter <= (logic_trackers_0_cmdCounter + 7'h01);
      end
      if(io_output_rsp_fire) begin
        io_output_rsp_payload_first <= io_output_rsp_payload_last;
      end
      if(when_BmbExclusiveMonitor_l126) begin
        logic_trackers_0_rspCounter <= (logic_trackers_0_rspCounter + 7'h01);
      end
      if(when_BmbExclusiveMonitor_l123_1) begin
        logic_trackers_1_cmdCounter <= (logic_trackers_1_cmdCounter + 7'h01);
      end
      if(when_BmbExclusiveMonitor_l126_1) begin
        logic_trackers_1_rspCounter <= (logic_trackers_1_rspCounter + 7'h01);
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(when_BmbExclusiveMonitor_l69) begin
      if(when_BmbExclusiveMonitor_l70) begin
        logic_sources_0_address <= io_input_cmd_payload_fragment_address;
        logic_sources_0_length <= io_input_cmd_payload_fragment_length;
        logic_sources_0_addressLowEnd <= logic_inputAddressLowEnd;
        logic_sources_0_context <= io_input_cmd_payload_fragment_context;
      end
    end
    if(when_BmbExclusiveMonitor_l69_1) begin
      if(when_BmbExclusiveMonitor_l70_1) begin
        logic_sources_1_address <= io_input_cmd_payload_fragment_address;
        logic_sources_1_length <= io_input_cmd_payload_fragment_length;
        logic_sources_1_addressLowEnd <= logic_inputAddressLowEnd;
        logic_sources_1_context <= io_input_cmd_payload_fragment_context;
      end
    end
    if(logic_trackers_0_hit) begin
      logic_trackers_0_done <= 1'b1;
    end
    if(logic_fence_start) begin
      logic_trackers_0_target <= logic_trackers_0_cmdCounter;
      logic_trackers_0_done <= 1'b0;
    end
    if(logic_trackers_1_hit) begin
      logic_trackers_1_done <= 1'b1;
    end
    if(logic_fence_start) begin
      logic_trackers_1_target <= logic_trackers_1_cmdCounter;
      logic_trackers_1_done <= 1'b0;
    end
  end


endmodule

module BmbInvalidateMonitor (
  input  wire          io_input_cmd_valid,
  output wire          io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [0:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [63:0]   io_input_cmd_payload_fragment_data,
  input  wire [7:0]    io_input_cmd_payload_fragment_mask,
  input  wire [4:0]    io_input_cmd_payload_fragment_context,
  output wire          io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [0:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire [4:0]    io_input_rsp_payload_fragment_context,
  output wire          io_input_inv_valid,
  input  wire          io_input_inv_ready,
  output wire          io_input_inv_payload_all,
  output wire [31:0]   io_input_inv_payload_address,
  output wire [5:0]    io_input_inv_payload_length,
  output wire [0:0]    io_input_inv_payload_source,
  input  wire          io_input_ack_valid,
  output wire          io_input_ack_ready,
  output wire          io_input_sync_valid,
  input  wire          io_input_sync_ready,
  output wire [0:0]    io_input_sync_payload_source,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  output wire [63:0]   io_output_cmd_payload_fragment_data,
  output wire [7:0]    io_output_cmd_payload_fragment_mask,
  output wire [43:0]   io_output_cmd_payload_fragment_context,
  input  wire          io_output_rsp_valid,
  output reg           io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_output_rsp_payload_fragment_data,
  input  wire [43:0]   io_output_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire                rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_push_ready;
  wire                rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_pop_valid;
  wire       [0:0]    rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_pop_payload;
  wire       [4:0]    rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_occupancy;
  wire       [4:0]    rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_availability;
  wire       [4:0]    cmdLogic_cmdContext_context;
  wire       [31:0]   cmdLogic_cmdContext_address;
  wire       [5:0]    cmdLogic_cmdContext_length;
  wire                cmdLogic_cmdContext_write;
  wire       [4:0]    rspLogic_rspContext_context;
  wire       [31:0]   rspLogic_rspContext_address;
  wire       [5:0]    rspLogic_rspContext_length;
  wire                rspLogic_rspContext_write;
  wire       [43:0]   _zz_rspLogic_rspContext_context;
  wire                rspLogic_rspToRsp_valid;
  wire                rspLogic_rspToRsp_ready;
  wire                rspLogic_rspToRsp_payload_last;
  wire       [0:0]    rspLogic_rspToRsp_payload_fragment_source;
  wire       [0:0]    rspLogic_rspToRsp_payload_fragment_opcode;
  wire       [63:0]   rspLogic_rspToRsp_payload_fragment_data;
  wire       [43:0]   rspLogic_rspToRsp_payload_fragment_context;
  wire                rspLogic_rspToInv_valid;
  reg                 rspLogic_rspToInv_ready;
  wire                rspLogic_rspToInv_payload_last;
  wire       [0:0]    rspLogic_rspToInv_payload_fragment_source;
  wire       [0:0]    rspLogic_rspToInv_payload_fragment_opcode;
  wire       [63:0]   rspLogic_rspToInv_payload_fragment_data;
  wire       [43:0]   rspLogic_rspToInv_payload_fragment_context;
  wire                rspLogic_rspToSync_valid;
  wire                rspLogic_rspToSync_ready;
  wire                rspLogic_rspToSync_payload_last;
  wire       [0:0]    rspLogic_rspToSync_payload_fragment_source;
  wire       [0:0]    rspLogic_rspToSync_payload_fragment_opcode;
  wire       [63:0]   rspLogic_rspToSync_payload_fragment_data;
  wire       [43:0]   rspLogic_rspToSync_payload_fragment_context;
  reg                 io_output_rsp_fork3_logic_linkEnable_0;
  reg                 io_output_rsp_fork3_logic_linkEnable_1;
  reg                 io_output_rsp_fork3_logic_linkEnable_2;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                when_Stream_l1063_2;
  wire                rspLogic_rspToRsp_fire;
  wire                rspLogic_rspToInv_fire;
  wire                rspLogic_rspToSync_fire;
  wire                when_Stream_l445;
  reg                 rspLogic_rspToInvFiltred_valid;
  wire                rspLogic_rspToInvFiltred_ready;
  wire                rspLogic_rspToInvFiltred_payload_last;
  wire       [0:0]    rspLogic_rspToInvFiltred_payload_fragment_source;
  wire       [0:0]    rspLogic_rspToInvFiltred_payload_fragment_opcode;
  wire       [63:0]   rspLogic_rspToInvFiltred_payload_fragment_data;
  wire       [43:0]   rspLogic_rspToInvFiltred_payload_fragment_context;
  wire                rspLogic_rspToSync_translated_valid;
  reg                 rspLogic_rspToSync_translated_ready;
  wire       [0:0]    rspLogic_rspToSync_translated_payload;
  wire                when_Stream_l445_1;
  reg                 rspLogic_rspToSyncFiltred_valid;
  wire                rspLogic_rspToSyncFiltred_ready;
  wire       [0:0]    rspLogic_rspToSyncFiltred_payload;
  wire                rspLogic_rspToSyncFiltred_s2mPipe_valid;
  wire                rspLogic_rspToSyncFiltred_s2mPipe_ready;
  wire       [0:0]    rspLogic_rspToSyncFiltred_s2mPipe_payload;
  reg                 rspLogic_rspToSyncFiltred_rValidN;
  reg        [0:0]    rspLogic_rspToSyncFiltred_rData;
  wire                io_input_ack_fire;

  StreamFifo rspLogic_rspToSyncFiltred_s2mPipe_fifo (
    .io_push_valid              (rspLogic_rspToSyncFiltred_s2mPipe_valid                    ), //i
    .io_push_ready              (rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_push_ready       ), //o
    .io_push_payload            (rspLogic_rspToSyncFiltred_s2mPipe_payload                  ), //i
    .io_pop_valid               (rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_pop_valid        ), //o
    .io_pop_ready               (io_input_ack_fire                                          ), //i
    .io_pop_payload             (rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_pop_payload      ), //o
    .io_flush                   (1'b0                                                       ), //i
    .io_occupancy               (rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_occupancy[4:0]   ), //o
    .io_availability            (rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_availability[4:0]), //o
    .io_systemClk               (io_systemClk                                               ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                                 )  //i
  );
  assign cmdLogic_cmdContext_context = io_input_cmd_payload_fragment_context;
  assign cmdLogic_cmdContext_write = (io_input_cmd_payload_fragment_opcode == 1'b1);
  assign cmdLogic_cmdContext_address = io_input_cmd_payload_fragment_address;
  assign cmdLogic_cmdContext_length = io_input_cmd_payload_fragment_length;
  assign io_output_cmd_valid = io_input_cmd_valid;
  assign io_input_cmd_ready = io_output_cmd_ready;
  assign io_output_cmd_payload_last = io_input_cmd_payload_last;
  assign io_output_cmd_payload_fragment_source = io_input_cmd_payload_fragment_source;
  assign io_output_cmd_payload_fragment_opcode = io_input_cmd_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = io_input_cmd_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = io_input_cmd_payload_fragment_length;
  assign io_output_cmd_payload_fragment_data = io_input_cmd_payload_fragment_data;
  assign io_output_cmd_payload_fragment_mask = io_input_cmd_payload_fragment_mask;
  assign io_output_cmd_payload_fragment_context = {cmdLogic_cmdContext_write,{cmdLogic_cmdContext_length,{cmdLogic_cmdContext_address,cmdLogic_cmdContext_context}}};
  assign _zz_rspLogic_rspContext_context = io_output_rsp_payload_fragment_context;
  assign rspLogic_rspContext_context = _zz_rspLogic_rspContext_context[4 : 0];
  assign rspLogic_rspContext_address = _zz_rspLogic_rspContext_context[36 : 5];
  assign rspLogic_rspContext_length = _zz_rspLogic_rspContext_context[42 : 37];
  assign rspLogic_rspContext_write = _zz_rspLogic_rspContext_context[43];
  always @(*) begin
    io_output_rsp_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_output_rsp_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_output_rsp_ready = 1'b0;
    end
    if(when_Stream_l1063_2) begin
      io_output_rsp_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! rspLogic_rspToRsp_ready) && io_output_rsp_fork3_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! rspLogic_rspToInv_ready) && io_output_rsp_fork3_logic_linkEnable_1);
  assign when_Stream_l1063_2 = ((! rspLogic_rspToSync_ready) && io_output_rsp_fork3_logic_linkEnable_2);
  assign rspLogic_rspToRsp_valid = (io_output_rsp_valid && io_output_rsp_fork3_logic_linkEnable_0);
  assign rspLogic_rspToRsp_payload_last = io_output_rsp_payload_last;
  assign rspLogic_rspToRsp_payload_fragment_source = io_output_rsp_payload_fragment_source;
  assign rspLogic_rspToRsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign rspLogic_rspToRsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign rspLogic_rspToRsp_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign rspLogic_rspToRsp_fire = (rspLogic_rspToRsp_valid && rspLogic_rspToRsp_ready);
  assign rspLogic_rspToInv_valid = (io_output_rsp_valid && io_output_rsp_fork3_logic_linkEnable_1);
  assign rspLogic_rspToInv_payload_last = io_output_rsp_payload_last;
  assign rspLogic_rspToInv_payload_fragment_source = io_output_rsp_payload_fragment_source;
  assign rspLogic_rspToInv_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign rspLogic_rspToInv_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign rspLogic_rspToInv_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign rspLogic_rspToInv_fire = (rspLogic_rspToInv_valid && rspLogic_rspToInv_ready);
  assign rspLogic_rspToSync_valid = (io_output_rsp_valid && io_output_rsp_fork3_logic_linkEnable_2);
  assign rspLogic_rspToSync_payload_last = io_output_rsp_payload_last;
  assign rspLogic_rspToSync_payload_fragment_source = io_output_rsp_payload_fragment_source;
  assign rspLogic_rspToSync_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign rspLogic_rspToSync_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign rspLogic_rspToSync_payload_fragment_context = io_output_rsp_payload_fragment_context;
  assign rspLogic_rspToSync_fire = (rspLogic_rspToSync_valid && rspLogic_rspToSync_ready);
  assign io_input_rsp_valid = rspLogic_rspToRsp_valid;
  assign rspLogic_rspToRsp_ready = io_input_rsp_ready;
  assign io_input_rsp_payload_last = rspLogic_rspToRsp_payload_last;
  assign io_input_rsp_payload_fragment_source = rspLogic_rspToRsp_payload_fragment_source;
  assign io_input_rsp_payload_fragment_opcode = rspLogic_rspToRsp_payload_fragment_opcode;
  assign io_input_rsp_payload_fragment_data = rspLogic_rspToRsp_payload_fragment_data;
  assign io_input_rsp_payload_fragment_context = rspLogic_rspContext_context;
  assign when_Stream_l445 = (! rspLogic_rspContext_write);
  always @(*) begin
    rspLogic_rspToInvFiltred_valid = rspLogic_rspToInv_valid;
    if(when_Stream_l445) begin
      rspLogic_rspToInvFiltred_valid = 1'b0;
    end
  end

  always @(*) begin
    rspLogic_rspToInv_ready = rspLogic_rspToInvFiltred_ready;
    if(when_Stream_l445) begin
      rspLogic_rspToInv_ready = 1'b1;
    end
  end

  assign rspLogic_rspToInvFiltred_payload_last = rspLogic_rspToInv_payload_last;
  assign rspLogic_rspToInvFiltred_payload_fragment_source = rspLogic_rspToInv_payload_fragment_source;
  assign rspLogic_rspToInvFiltred_payload_fragment_opcode = rspLogic_rspToInv_payload_fragment_opcode;
  assign rspLogic_rspToInvFiltred_payload_fragment_data = rspLogic_rspToInv_payload_fragment_data;
  assign rspLogic_rspToInvFiltred_payload_fragment_context = rspLogic_rspToInv_payload_fragment_context;
  assign io_input_inv_valid = rspLogic_rspToInvFiltred_valid;
  assign rspLogic_rspToInvFiltred_ready = io_input_inv_ready;
  assign io_input_inv_payload_address = rspLogic_rspContext_address;
  assign io_input_inv_payload_length = rspLogic_rspContext_length;
  assign io_input_inv_payload_source = rspLogic_rspToInvFiltred_payload_fragment_source;
  assign io_input_inv_payload_all = 1'b0;
  assign rspLogic_rspToSync_translated_valid = rspLogic_rspToSync_valid;
  assign rspLogic_rspToSync_ready = rspLogic_rspToSync_translated_ready;
  assign rspLogic_rspToSync_translated_payload = rspLogic_rspToInv_payload_fragment_source;
  assign when_Stream_l445_1 = (! rspLogic_rspContext_write);
  always @(*) begin
    rspLogic_rspToSyncFiltred_valid = rspLogic_rspToSync_translated_valid;
    if(when_Stream_l445_1) begin
      rspLogic_rspToSyncFiltred_valid = 1'b0;
    end
  end

  always @(*) begin
    rspLogic_rspToSync_translated_ready = rspLogic_rspToSyncFiltred_ready;
    if(when_Stream_l445_1) begin
      rspLogic_rspToSync_translated_ready = 1'b1;
    end
  end

  assign rspLogic_rspToSyncFiltred_payload = rspLogic_rspToSync_translated_payload;
  assign rspLogic_rspToSyncFiltred_ready = rspLogic_rspToSyncFiltred_rValidN;
  assign rspLogic_rspToSyncFiltred_s2mPipe_valid = (rspLogic_rspToSyncFiltred_valid || (! rspLogic_rspToSyncFiltred_rValidN));
  assign rspLogic_rspToSyncFiltred_s2mPipe_payload = (rspLogic_rspToSyncFiltred_rValidN ? rspLogic_rspToSyncFiltred_payload : rspLogic_rspToSyncFiltred_rData);
  assign rspLogic_rspToSyncFiltred_s2mPipe_ready = rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_push_ready;
  assign io_input_ack_fire = (io_input_ack_valid && io_input_ack_ready);
  assign io_input_sync_valid = io_input_ack_valid;
  assign io_input_ack_ready = io_input_sync_ready;
  assign io_input_sync_payload_source = rspLogic_rspToSyncFiltred_s2mPipe_fifo_io_pop_payload;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      io_output_rsp_fork3_logic_linkEnable_0 <= 1'b1;
      io_output_rsp_fork3_logic_linkEnable_1 <= 1'b1;
      io_output_rsp_fork3_logic_linkEnable_2 <= 1'b1;
      rspLogic_rspToSyncFiltred_rValidN <= 1'b1;
    end else begin
      if(rspLogic_rspToRsp_fire) begin
        io_output_rsp_fork3_logic_linkEnable_0 <= 1'b0;
      end
      if(rspLogic_rspToInv_fire) begin
        io_output_rsp_fork3_logic_linkEnable_1 <= 1'b0;
      end
      if(rspLogic_rspToSync_fire) begin
        io_output_rsp_fork3_logic_linkEnable_2 <= 1'b0;
      end
      if(io_output_rsp_ready) begin
        io_output_rsp_fork3_logic_linkEnable_0 <= 1'b1;
        io_output_rsp_fork3_logic_linkEnable_1 <= 1'b1;
        io_output_rsp_fork3_logic_linkEnable_2 <= 1'b1;
      end
      if(rspLogic_rspToSyncFiltred_valid) begin
        rspLogic_rspToSyncFiltred_rValidN <= 1'b0;
      end
      if(rspLogic_rspToSyncFiltred_s2mPipe_ready) begin
        rspLogic_rspToSyncFiltred_rValidN <= 1'b1;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(rspLogic_rspToSyncFiltred_ready) begin
      rspLogic_rspToSyncFiltred_rData <= rspLogic_rspToSyncFiltred_payload;
    end
  end


endmodule

module BmbArbiter (
  input  wire          io_inputs_0_cmd_valid,
  output wire          io_inputs_0_cmd_ready,
  input  wire          io_inputs_0_cmd_payload_last,
  input  wire [0:0]    io_inputs_0_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_0_cmd_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_cmd_payload_fragment_length,
  output wire          io_inputs_0_rsp_valid,
  input  wire          io_inputs_0_rsp_ready,
  output wire          io_inputs_0_rsp_payload_last,
  output wire [0:0]    io_inputs_0_rsp_payload_fragment_opcode,
  output wire [63:0]   io_inputs_0_rsp_payload_fragment_data,
  input  wire          io_inputs_1_cmd_valid,
  output wire          io_inputs_1_cmd_ready,
  input  wire          io_inputs_1_cmd_payload_last,
  input  wire [0:0]    io_inputs_1_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_1_cmd_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_cmd_payload_fragment_length,
  output wire          io_inputs_1_rsp_valid,
  input  wire          io_inputs_1_rsp_ready,
  output wire          io_inputs_1_rsp_payload_last,
  output wire [0:0]    io_inputs_1_rsp_payload_fragment_opcode,
  output wire [63:0]   io_inputs_1_rsp_payload_fragment_data,
  output wire          io_output_cmd_valid,
  input  wire          io_output_cmd_ready,
  output wire          io_output_cmd_payload_last,
  output wire [0:0]    io_output_cmd_payload_fragment_source,
  output wire [0:0]    io_output_cmd_payload_fragment_opcode,
  output wire [31:0]   io_output_cmd_payload_fragment_address,
  output wire [5:0]    io_output_cmd_payload_fragment_length,
  input  wire          io_output_rsp_valid,
  output wire          io_output_rsp_ready,
  input  wire          io_output_rsp_payload_last,
  input  wire [0:0]    io_output_rsp_payload_fragment_source,
  input  wire [0:0]    io_output_rsp_payload_fragment_opcode,
  input  wire [63:0]   io_output_rsp_payload_fragment_data,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire                memory_arbiter_io_inputs_0_ready;
  wire                memory_arbiter_io_inputs_1_ready;
  wire                memory_arbiter_io_output_valid;
  wire                memory_arbiter_io_output_payload_last;
  wire       [0:0]    memory_arbiter_io_output_payload_fragment_source;
  wire       [0:0]    memory_arbiter_io_output_payload_fragment_opcode;
  wire       [31:0]   memory_arbiter_io_output_payload_fragment_address;
  wire       [5:0]    memory_arbiter_io_output_payload_fragment_length;
  wire       [0:0]    memory_arbiter_io_chosen;
  wire       [1:0]    memory_arbiter_io_chosenOH;
  wire       [1:0]    _zz_io_output_cmd_payload_fragment_source;
  reg                 _zz_io_output_rsp_ready;
  wire       [0:0]    memory_rspSel;

  assign _zz_io_output_cmd_payload_fragment_source = {memory_arbiter_io_output_payload_fragment_source,memory_arbiter_io_chosen};
  StreamArbiter_2 memory_arbiter (
    .io_inputs_0_valid                    (io_inputs_0_cmd_valid                                  ), //i
    .io_inputs_0_ready                    (memory_arbiter_io_inputs_0_ready                       ), //o
    .io_inputs_0_payload_last             (io_inputs_0_cmd_payload_last                           ), //i
    .io_inputs_0_payload_fragment_source  (1'b0                                                   ), //i
    .io_inputs_0_payload_fragment_opcode  (io_inputs_0_cmd_payload_fragment_opcode                ), //i
    .io_inputs_0_payload_fragment_address (io_inputs_0_cmd_payload_fragment_address[31:0]         ), //i
    .io_inputs_0_payload_fragment_length  (io_inputs_0_cmd_payload_fragment_length[5:0]           ), //i
    .io_inputs_1_valid                    (io_inputs_1_cmd_valid                                  ), //i
    .io_inputs_1_ready                    (memory_arbiter_io_inputs_1_ready                       ), //o
    .io_inputs_1_payload_last             (io_inputs_1_cmd_payload_last                           ), //i
    .io_inputs_1_payload_fragment_source  (1'b0                                                   ), //i
    .io_inputs_1_payload_fragment_opcode  (io_inputs_1_cmd_payload_fragment_opcode                ), //i
    .io_inputs_1_payload_fragment_address (io_inputs_1_cmd_payload_fragment_address[31:0]         ), //i
    .io_inputs_1_payload_fragment_length  (io_inputs_1_cmd_payload_fragment_length[5:0]           ), //i
    .io_output_valid                      (memory_arbiter_io_output_valid                         ), //o
    .io_output_ready                      (io_output_cmd_ready                                    ), //i
    .io_output_payload_last               (memory_arbiter_io_output_payload_last                  ), //o
    .io_output_payload_fragment_source    (memory_arbiter_io_output_payload_fragment_source       ), //o
    .io_output_payload_fragment_opcode    (memory_arbiter_io_output_payload_fragment_opcode       ), //o
    .io_output_payload_fragment_address   (memory_arbiter_io_output_payload_fragment_address[31:0]), //o
    .io_output_payload_fragment_length    (memory_arbiter_io_output_payload_fragment_length[5:0]  ), //o
    .io_chosen                            (memory_arbiter_io_chosen                               ), //o
    .io_chosenOH                          (memory_arbiter_io_chosenOH[1:0]                        ), //o
    .io_systemClk                         (io_systemClk                                           ), //i
    .systemCd_logic_outputReset           (systemCd_logic_outputReset                             )  //i
  );
  always @(*) begin
    case(memory_rspSel)
      1'b0 : _zz_io_output_rsp_ready = io_inputs_0_rsp_ready;
      default : _zz_io_output_rsp_ready = io_inputs_1_rsp_ready;
    endcase
  end

  assign io_inputs_0_cmd_ready = memory_arbiter_io_inputs_0_ready;
  assign io_inputs_1_cmd_ready = memory_arbiter_io_inputs_1_ready;
  assign io_output_cmd_valid = memory_arbiter_io_output_valid;
  assign io_output_cmd_payload_last = memory_arbiter_io_output_payload_last;
  assign io_output_cmd_payload_fragment_opcode = memory_arbiter_io_output_payload_fragment_opcode;
  assign io_output_cmd_payload_fragment_address = memory_arbiter_io_output_payload_fragment_address;
  assign io_output_cmd_payload_fragment_length = memory_arbiter_io_output_payload_fragment_length;
  assign io_output_cmd_payload_fragment_source = _zz_io_output_cmd_payload_fragment_source[0:0];
  assign memory_rspSel = io_output_rsp_payload_fragment_source[0 : 0];
  assign io_inputs_0_rsp_valid = (io_output_rsp_valid && (memory_rspSel == 1'b0));
  assign io_inputs_0_rsp_payload_last = io_output_rsp_payload_last;
  assign io_inputs_0_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_inputs_0_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_inputs_1_rsp_valid = (io_output_rsp_valid && (memory_rspSel == 1'b1));
  assign io_inputs_1_rsp_payload_last = io_output_rsp_payload_last;
  assign io_inputs_1_rsp_payload_fragment_opcode = io_output_rsp_payload_fragment_opcode;
  assign io_inputs_1_rsp_payload_fragment_data = io_output_rsp_payload_fragment_data;
  assign io_output_rsp_ready = _zz_io_output_rsp_ready;

endmodule

module DebugTransportModuleTunneled (
  input  wire          io_instruction_tdi,
  input  wire          io_instruction_enable,
  input  wire          io_instruction_capture,
  input  wire          io_instruction_shift,
  input  wire          io_instruction_update,
  input  wire          io_instruction_reset,
  output wire          io_instruction_tdo,
  output wire          io_bus_cmd_valid,
  input  wire          io_bus_cmd_ready,
  output wire          io_bus_cmd_payload_write,
  output wire [31:0]   io_bus_cmd_payload_data,
  output wire [6:0]    io_bus_cmd_payload_address,
  input  wire          io_bus_rsp_valid,
  input  wire          io_bus_rsp_payload_error,
  input  wire [31:0]   io_bus_rsp_payload_data,
  input  wire          jtagCtrl_tck,
  input  wire          io_systemClk,
  input  wire          debugCd_logic_outputReset
);
  localparam DebugCaptureOp_SUCCESS = 2'd0;
  localparam DebugCaptureOp_RESERVED = 2'd1;
  localparam DebugCaptureOp_FAILED = 2'd2;
  localparam DebugCaptureOp_OVERRUN = 2'd3;
  localparam DebugUpdateOp_NOP = 2'd0;
  localparam DebugUpdateOp_READ = 2'd1;
  localparam DebugUpdateOp_WRITE = 2'd2;
  localparam DebugUpdateOp_RESERVED = 2'd3;

  wire                logic_jtagLogic_dmiCmd_ccToggle_io_output_valid;
  wire                logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_write;
  wire       [31:0]   logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_data;
  wire       [6:0]    logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_address;
  wire                logic_systemLogic_bus_rsp_ccToggle_io_output_valid;
  wire                logic_systemLogic_bus_rsp_ccToggle_io_output_payload_error;
  wire       [31:0]   logic_systemLogic_bus_rsp_ccToggle_io_output_payload_data;
  reg        [1:0]    logic_jtagLogic_dmiStat_value_aheadValue;
  reg        [13:0]   tap_shiftBuffer;
  reg        [5:0]    tap_instruction;
  reg                 tap_sendCapture;
  reg                 tap_sendShift;
  reg                 tap_sendUpdate;
  wire                when_JtagTunnel_l30;
  reg                 io_instruction_tdi_delay_1;
  reg                 io_instruction_tdi_delay_2;
  reg                 io_instruction_tdi_delay_3;
  reg                 io_instruction_tdi_delay_4;
  reg                 io_instruction_tdi_delay_5;
  reg                 io_instruction_tdi_delay_6;
  reg                 io_instruction_tdi_delay_7;
  reg                 io_instruction_tdi_delay_8;
  reg                 tap_tdiBuffer;
  reg                 tap_tdoBuffer;
  reg                 tap_tdoBuffer_delay_1;
  reg                 tap_tdoBuffer_delay_2;
  reg                 tap_tdoBuffer_delay_3;
  reg                 tap_tdoShifter;
  wire                logic_jtagLogic_dmiCmd_valid;
  wire                logic_jtagLogic_dmiCmd_payload_write;
  wire       [31:0]   logic_jtagLogic_dmiCmd_payload_data;
  wire       [6:0]    logic_jtagLogic_dmiCmd_payload_address;
  wire                logic_jtagLogic_dmiRsp_valid;
  wire                logic_jtagLogic_dmiRsp_payload_error;
  wire       [31:0]   logic_jtagLogic_dmiRsp_payload_data;
  wire       [31:0]   logic_jtagLogic_dtmcs_captureData;
  wire       [31:0]   logic_jtagLogic_dtmcs_updateData;
  wire                logic_jtagLogic_dtmcs_captureValid;
  wire                logic_jtagLogic_dtmcs_updateValid;
  wire                logic_jtagLogic_dtmcs_logic_ctrl_tdi;
  wire                logic_jtagLogic_dtmcs_logic_ctrl_enable;
  wire                logic_jtagLogic_dtmcs_logic_ctrl_capture;
  wire                logic_jtagLogic_dtmcs_logic_ctrl_shift;
  wire                logic_jtagLogic_dtmcs_logic_ctrl_update;
  wire                logic_jtagLogic_dtmcs_logic_ctrl_reset;
  wire                logic_jtagLogic_dtmcs_logic_ctrl_tdo;
  reg        [31:0]   logic_jtagLogic_dtmcs_logic_store;
  wire                when_JtagTunnel_l53;
  wire       [1:0]    logic_jtagLogic_dmi_captureData_op;
  wire       [31:0]   logic_jtagLogic_dmi_captureData_data;
  wire       [6:0]    logic_jtagLogic_dmi_captureData_padding;
  wire       [1:0]    logic_jtagLogic_dmi_updateData_op;
  wire       [31:0]   logic_jtagLogic_dmi_updateData_data;
  wire       [6:0]    logic_jtagLogic_dmi_updateData_address;
  wire                logic_jtagLogic_dmi_captureValid;
  wire                logic_jtagLogic_dmi_updateValid;
  wire                logic_jtagLogic_dmi_logic_ctrl_tdi;
  wire                logic_jtagLogic_dmi_logic_ctrl_enable;
  wire                logic_jtagLogic_dmi_logic_ctrl_capture;
  wire                logic_jtagLogic_dmi_logic_ctrl_shift;
  wire                logic_jtagLogic_dmi_logic_ctrl_update;
  wire                logic_jtagLogic_dmi_logic_ctrl_reset;
  wire                logic_jtagLogic_dmi_logic_ctrl_tdo;
  reg        [40:0]   logic_jtagLogic_dmi_logic_store;
  wire       [1:0]    _zz_logic_jtagLogic_dmi_updateData_op;
  wire                when_JtagTunnel_l53_1;
  reg        [1:0]    logic_jtagLogic_dmiStat_value;
  reg                 logic_jtagLogic_dmiStat_failure;
  reg                 logic_jtagLogic_dmiStat_busy;
  reg                 logic_jtagLogic_dmiStat_clear;
  wire                when_DebugTransportModuleJtag_l30;
  reg                 logic_jtagLogic_pending;
  wire                logic_jtagLogic_trigger_dmiHardReset;
  wire                logic_jtagLogic_trigger_dmiReset;
  reg                 logic_jtagLogic_trigger_dmiCmd;
  reg        [31:0]   logic_jtagLogic_rspLogic_buffer;
  wire                when_DebugTransportModuleJtag_l78;
  wire                logic_systemLogic_bus_cmd_valid;
  wire                logic_systemLogic_bus_cmd_ready;
  wire                logic_systemLogic_bus_cmd_payload_write;
  wire       [31:0]   logic_systemLogic_bus_cmd_payload_data;
  wire       [6:0]    logic_systemLogic_bus_cmd_payload_address;
  wire                logic_systemLogic_bus_rsp_valid;
  wire                logic_systemLogic_bus_rsp_payload_error;
  wire       [31:0]   logic_systemLogic_bus_rsp_payload_data;
  wire                logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_valid;
  reg                 logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_ready;
  wire                logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_write;
  wire       [31:0]   logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_data;
  wire       [6:0]    logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_address;
  wire                logic_systemLogic_cmd_valid;
  wire                logic_systemLogic_cmd_ready;
  wire                logic_systemLogic_cmd_payload_write;
  wire       [31:0]   logic_systemLogic_cmd_payload_data;
  wire       [6:0]    logic_systemLogic_cmd_payload_address;
  reg                 logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rValid;
  wire                logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_fire;
  (* async_reg = "true" *) reg                 logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_write;
  (* async_reg = "true" *) reg        [31:0]   logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_data;
  (* async_reg = "true" *) reg        [6:0]    logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_address;
  wire                when_Stream_l375;
  `ifndef SYNTHESIS
  reg [63:0] logic_jtagLogic_dmiStat_value_aheadValue_string;
  reg [63:0] logic_jtagLogic_dmi_captureData_op_string;
  reg [63:0] logic_jtagLogic_dmi_updateData_op_string;
  reg [63:0] _zz_logic_jtagLogic_dmi_updateData_op_string;
  reg [63:0] logic_jtagLogic_dmiStat_value_string;
  `endif


  FlowCCByToggle logic_jtagLogic_dmiCmd_ccToggle (
    .io_input_valid            (logic_jtagLogic_dmiCmd_valid                                  ), //i
    .io_input_payload_write    (logic_jtagLogic_dmiCmd_payload_write                          ), //i
    .io_input_payload_data     (logic_jtagLogic_dmiCmd_payload_data[31:0]                     ), //i
    .io_input_payload_address  (logic_jtagLogic_dmiCmd_payload_address[6:0]                   ), //i
    .io_output_valid           (logic_jtagLogic_dmiCmd_ccToggle_io_output_valid               ), //o
    .io_output_payload_write   (logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_write       ), //o
    .io_output_payload_data    (logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_data[31:0]  ), //o
    .io_output_payload_address (logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_address[6:0]), //o
    .jtagCtrl_tck              (jtagCtrl_tck                                                  ), //i
    .io_systemClk              (io_systemClk                                                  ), //i
    .debugCd_logic_outputReset (debugCd_logic_outputReset                                     )  //i
  );
  FlowCCByToggle_1 logic_systemLogic_bus_rsp_ccToggle (
    .io_input_valid            (logic_systemLogic_bus_rsp_valid                                ), //i
    .io_input_payload_error    (logic_systemLogic_bus_rsp_payload_error                        ), //i
    .io_input_payload_data     (logic_systemLogic_bus_rsp_payload_data[31:0]                   ), //i
    .io_output_valid           (logic_systemLogic_bus_rsp_ccToggle_io_output_valid             ), //o
    .io_output_payload_error   (logic_systemLogic_bus_rsp_ccToggle_io_output_payload_error     ), //o
    .io_output_payload_data    (logic_systemLogic_bus_rsp_ccToggle_io_output_payload_data[31:0]), //o
    .io_systemClk              (io_systemClk                                                   ), //i
    .debugCd_logic_outputReset (debugCd_logic_outputReset                                      ), //i
    .jtagCtrl_tck              (jtagCtrl_tck                                                   )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(logic_jtagLogic_dmiStat_value_aheadValue)
      DebugCaptureOp_SUCCESS : logic_jtagLogic_dmiStat_value_aheadValue_string = "SUCCESS ";
      DebugCaptureOp_RESERVED : logic_jtagLogic_dmiStat_value_aheadValue_string = "RESERVED";
      DebugCaptureOp_FAILED : logic_jtagLogic_dmiStat_value_aheadValue_string = "FAILED  ";
      DebugCaptureOp_OVERRUN : logic_jtagLogic_dmiStat_value_aheadValue_string = "OVERRUN ";
      default : logic_jtagLogic_dmiStat_value_aheadValue_string = "????????";
    endcase
  end
  always @(*) begin
    case(logic_jtagLogic_dmi_captureData_op)
      DebugCaptureOp_SUCCESS : logic_jtagLogic_dmi_captureData_op_string = "SUCCESS ";
      DebugCaptureOp_RESERVED : logic_jtagLogic_dmi_captureData_op_string = "RESERVED";
      DebugCaptureOp_FAILED : logic_jtagLogic_dmi_captureData_op_string = "FAILED  ";
      DebugCaptureOp_OVERRUN : logic_jtagLogic_dmi_captureData_op_string = "OVERRUN ";
      default : logic_jtagLogic_dmi_captureData_op_string = "????????";
    endcase
  end
  always @(*) begin
    case(logic_jtagLogic_dmi_updateData_op)
      DebugUpdateOp_NOP : logic_jtagLogic_dmi_updateData_op_string = "NOP     ";
      DebugUpdateOp_READ : logic_jtagLogic_dmi_updateData_op_string = "READ    ";
      DebugUpdateOp_WRITE : logic_jtagLogic_dmi_updateData_op_string = "WRITE   ";
      DebugUpdateOp_RESERVED : logic_jtagLogic_dmi_updateData_op_string = "RESERVED";
      default : logic_jtagLogic_dmi_updateData_op_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_logic_jtagLogic_dmi_updateData_op)
      DebugUpdateOp_NOP : _zz_logic_jtagLogic_dmi_updateData_op_string = "NOP     ";
      DebugUpdateOp_READ : _zz_logic_jtagLogic_dmi_updateData_op_string = "READ    ";
      DebugUpdateOp_WRITE : _zz_logic_jtagLogic_dmi_updateData_op_string = "WRITE   ";
      DebugUpdateOp_RESERVED : _zz_logic_jtagLogic_dmi_updateData_op_string = "RESERVED";
      default : _zz_logic_jtagLogic_dmi_updateData_op_string = "????????";
    endcase
  end
  always @(*) begin
    case(logic_jtagLogic_dmiStat_value)
      DebugCaptureOp_SUCCESS : logic_jtagLogic_dmiStat_value_string = "SUCCESS ";
      DebugCaptureOp_RESERVED : logic_jtagLogic_dmiStat_value_string = "RESERVED";
      DebugCaptureOp_FAILED : logic_jtagLogic_dmiStat_value_string = "FAILED  ";
      DebugCaptureOp_OVERRUN : logic_jtagLogic_dmiStat_value_string = "OVERRUN ";
      default : logic_jtagLogic_dmiStat_value_string = "????????";
    endcase
  end
  `endif

  always @(*) begin
    logic_jtagLogic_dmiStat_value_aheadValue = logic_jtagLogic_dmiStat_value;
    if(when_DebugTransportModuleJtag_l30) begin
      if(logic_jtagLogic_dmiStat_failure) begin
        logic_jtagLogic_dmiStat_value_aheadValue = DebugCaptureOp_FAILED;
      end
      if(logic_jtagLogic_dmiStat_busy) begin
        logic_jtagLogic_dmiStat_value_aheadValue = DebugCaptureOp_OVERRUN;
      end
    end
    if(logic_jtagLogic_dmiStat_clear) begin
      logic_jtagLogic_dmiStat_value_aheadValue = DebugCaptureOp_SUCCESS;
    end
  end

  always @(*) begin
    tap_sendCapture = 1'b0;
    if(io_instruction_enable) begin
      if(io_instruction_capture) begin
        tap_sendCapture = 1'b1;
      end
    end
  end

  always @(*) begin
    tap_sendShift = 1'b0;
    if(io_instruction_enable) begin
      if(io_instruction_shift) begin
        tap_sendShift = 1'b1;
      end
    end
  end

  always @(*) begin
    tap_sendUpdate = 1'b0;
    if(io_instruction_enable) begin
      if(io_instruction_update) begin
        if(!when_JtagTunnel_l30) begin
          tap_sendUpdate = 1'b1;
        end
      end
    end
  end

  assign when_JtagTunnel_l30 = (! tap_shiftBuffer[13]);
  always @(*) begin
    tap_tdoBuffer = 1'b0;
    if(when_JtagTunnel_l53) begin
      tap_tdoBuffer = logic_jtagLogic_dtmcs_logic_ctrl_tdo;
    end
    if(when_JtagTunnel_l53_1) begin
      tap_tdoBuffer = logic_jtagLogic_dmi_logic_ctrl_tdo;
    end
  end

  assign io_instruction_tdo = tap_tdoShifter;
  assign logic_jtagLogic_dtmcs_captureValid = ((tap_instruction == 6'h10) && tap_sendCapture);
  assign logic_jtagLogic_dtmcs_updateValid = ((tap_instruction == 6'h10) && tap_sendUpdate);
  assign logic_jtagLogic_dtmcs_logic_ctrl_tdo = logic_jtagLogic_dtmcs_logic_store[0];
  assign logic_jtagLogic_dtmcs_updateData = logic_jtagLogic_dtmcs_logic_store;
  assign when_JtagTunnel_l53 = (tap_instruction == 6'h10);
  assign logic_jtagLogic_dtmcs_logic_ctrl_tdi = tap_tdiBuffer;
  assign logic_jtagLogic_dtmcs_logic_ctrl_enable = when_JtagTunnel_l53;
  assign logic_jtagLogic_dtmcs_logic_ctrl_capture = (when_JtagTunnel_l53 && tap_sendCapture);
  assign logic_jtagLogic_dtmcs_logic_ctrl_shift = (when_JtagTunnel_l53 && tap_sendShift);
  assign logic_jtagLogic_dtmcs_logic_ctrl_update = (when_JtagTunnel_l53 && tap_sendUpdate);
  assign logic_jtagLogic_dtmcs_logic_ctrl_reset = io_instruction_reset;
  assign logic_jtagLogic_dmi_captureValid = ((tap_instruction == 6'h11) && tap_sendCapture);
  assign logic_jtagLogic_dmi_updateValid = ((tap_instruction == 6'h11) && tap_sendUpdate);
  assign logic_jtagLogic_dmi_logic_ctrl_tdo = logic_jtagLogic_dmi_logic_store[0];
  assign _zz_logic_jtagLogic_dmi_updateData_op = logic_jtagLogic_dmi_logic_store[1 : 0];
  assign logic_jtagLogic_dmi_updateData_op = _zz_logic_jtagLogic_dmi_updateData_op;
  assign logic_jtagLogic_dmi_updateData_data = logic_jtagLogic_dmi_logic_store[33 : 2];
  assign logic_jtagLogic_dmi_updateData_address = logic_jtagLogic_dmi_logic_store[40 : 34];
  assign when_JtagTunnel_l53_1 = (tap_instruction == 6'h11);
  assign logic_jtagLogic_dmi_logic_ctrl_tdi = tap_tdiBuffer;
  assign logic_jtagLogic_dmi_logic_ctrl_enable = when_JtagTunnel_l53_1;
  assign logic_jtagLogic_dmi_logic_ctrl_capture = (when_JtagTunnel_l53_1 && tap_sendCapture);
  assign logic_jtagLogic_dmi_logic_ctrl_shift = (when_JtagTunnel_l53_1 && tap_sendShift);
  assign logic_jtagLogic_dmi_logic_ctrl_update = (when_JtagTunnel_l53_1 && tap_sendUpdate);
  assign logic_jtagLogic_dmi_logic_ctrl_reset = io_instruction_reset;
  always @(*) begin
    logic_jtagLogic_dmiStat_failure = 1'b0;
    if(logic_jtagLogic_dmi_updateValid) begin
      case(logic_jtagLogic_dmi_updateData_op)
        DebugUpdateOp_NOP : begin
        end
        DebugUpdateOp_READ : begin
        end
        DebugUpdateOp_WRITE : begin
        end
        default : begin
          logic_jtagLogic_dmiStat_failure = 1'b1;
        end
      endcase
    end
    if(logic_jtagLogic_dmiRsp_valid) begin
      if(logic_jtagLogic_dmiRsp_payload_error) begin
        logic_jtagLogic_dmiStat_failure = 1'b1;
      end
    end
  end

  always @(*) begin
    logic_jtagLogic_dmiStat_busy = 1'b0;
    if(when_DebugTransportModuleJtag_l78) begin
      logic_jtagLogic_dmiStat_busy = 1'b1;
    end
  end

  always @(*) begin
    logic_jtagLogic_dmiStat_clear = 1'b0;
    if(logic_jtagLogic_trigger_dmiReset) begin
      logic_jtagLogic_dmiStat_clear = 1'b1;
    end
    if(logic_jtagLogic_trigger_dmiHardReset) begin
      logic_jtagLogic_dmiStat_clear = 1'b1;
    end
  end

  assign when_DebugTransportModuleJtag_l30 = (logic_jtagLogic_dmiStat_value == DebugCaptureOp_SUCCESS);
  assign logic_jtagLogic_trigger_dmiHardReset = ((logic_jtagLogic_dtmcs_updateData[17] && logic_jtagLogic_dtmcs_updateValid) || io_instruction_reset);
  assign logic_jtagLogic_trigger_dmiReset = ((logic_jtagLogic_dtmcs_updateData[16] && logic_jtagLogic_dtmcs_updateValid) || io_instruction_reset);
  always @(*) begin
    logic_jtagLogic_trigger_dmiCmd = 1'b0;
    if(logic_jtagLogic_dmi_updateValid) begin
      case(logic_jtagLogic_dmi_updateData_op)
        DebugUpdateOp_NOP : begin
        end
        DebugUpdateOp_READ : begin
          logic_jtagLogic_trigger_dmiCmd = 1'b1;
        end
        DebugUpdateOp_WRITE : begin
          logic_jtagLogic_trigger_dmiCmd = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  assign logic_jtagLogic_dtmcs_captureData = {{{{17'h0,3'b111},logic_jtagLogic_dmiStat_value},6'h07},4'b0001};
  assign logic_jtagLogic_dmiCmd_valid = logic_jtagLogic_trigger_dmiCmd;
  assign logic_jtagLogic_dmiCmd_payload_write = (logic_jtagLogic_dmi_updateData_op == DebugUpdateOp_WRITE);
  assign logic_jtagLogic_dmiCmd_payload_address = logic_jtagLogic_dmi_updateData_address;
  assign logic_jtagLogic_dmiCmd_payload_data = logic_jtagLogic_dmi_updateData_data;
  assign logic_jtagLogic_dmi_captureData_op = logic_jtagLogic_dmiStat_value_aheadValue;
  assign logic_jtagLogic_dmi_captureData_data = logic_jtagLogic_rspLogic_buffer;
  assign logic_jtagLogic_dmi_captureData_padding = 7'h0;
  assign when_DebugTransportModuleJtag_l78 = (logic_jtagLogic_dmi_captureValid && logic_jtagLogic_pending);
  assign logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_valid = logic_jtagLogic_dmiCmd_ccToggle_io_output_valid;
  assign logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_write = logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_write;
  assign logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_data = logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_data;
  assign logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_address = logic_jtagLogic_dmiCmd_ccToggle_io_output_payload_address;
  assign logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_fire = (logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_valid && logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_ready);
  always @(*) begin
    logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_ready = logic_systemLogic_cmd_ready;
    if(when_Stream_l375) begin
      logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_systemLogic_cmd_valid);
  assign logic_systemLogic_cmd_valid = logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rValid;
  assign logic_systemLogic_cmd_payload_write = logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_write;
  assign logic_systemLogic_cmd_payload_data = logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_data;
  assign logic_systemLogic_cmd_payload_address = logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_address;
  assign logic_systemLogic_bus_cmd_valid = logic_systemLogic_cmd_valid;
  assign logic_systemLogic_cmd_ready = logic_systemLogic_bus_cmd_ready;
  assign logic_systemLogic_bus_cmd_payload_write = logic_systemLogic_cmd_payload_write;
  assign logic_systemLogic_bus_cmd_payload_data = logic_systemLogic_cmd_payload_data;
  assign logic_systemLogic_bus_cmd_payload_address = logic_systemLogic_cmd_payload_address;
  assign logic_jtagLogic_dmiRsp_valid = logic_systemLogic_bus_rsp_ccToggle_io_output_valid;
  assign logic_jtagLogic_dmiRsp_payload_error = logic_systemLogic_bus_rsp_ccToggle_io_output_payload_error;
  assign logic_jtagLogic_dmiRsp_payload_data = logic_systemLogic_bus_rsp_ccToggle_io_output_payload_data;
  assign io_bus_cmd_valid = logic_systemLogic_bus_cmd_valid;
  assign logic_systemLogic_bus_cmd_ready = io_bus_cmd_ready;
  assign io_bus_cmd_payload_write = logic_systemLogic_bus_cmd_payload_write;
  assign io_bus_cmd_payload_data = logic_systemLogic_bus_cmd_payload_data;
  assign io_bus_cmd_payload_address = logic_systemLogic_bus_cmd_payload_address;
  assign logic_systemLogic_bus_rsp_valid = io_bus_rsp_valid;
  assign logic_systemLogic_bus_rsp_payload_error = io_bus_rsp_payload_error;
  assign logic_systemLogic_bus_rsp_payload_data = io_bus_rsp_payload_data;
  always @(posedge jtagCtrl_tck) begin
    if(io_instruction_reset) begin
      tap_instruction <= 6'h0;
    end
    if(io_instruction_enable) begin
      if(io_instruction_shift) begin
        tap_shiftBuffer <= ({io_instruction_tdi,tap_shiftBuffer} >>> 1'd1);
      end
      if(io_instruction_update) begin
        if(when_JtagTunnel_l30) begin
          tap_instruction <= tap_shiftBuffer[5:0];
        end
      end
    end
    io_instruction_tdi_delay_1 <= io_instruction_tdi;
    io_instruction_tdi_delay_2 <= io_instruction_tdi_delay_1;
    io_instruction_tdi_delay_3 <= io_instruction_tdi_delay_2;
    io_instruction_tdi_delay_4 <= io_instruction_tdi_delay_3;
    io_instruction_tdi_delay_5 <= io_instruction_tdi_delay_4;
    io_instruction_tdi_delay_6 <= io_instruction_tdi_delay_5;
    io_instruction_tdi_delay_7 <= io_instruction_tdi_delay_6;
    io_instruction_tdi_delay_8 <= io_instruction_tdi_delay_7;
    tap_tdiBuffer <= io_instruction_tdi_delay_8;
    tap_tdoBuffer_delay_1 <= tap_tdoBuffer;
    tap_tdoBuffer_delay_2 <= tap_tdoBuffer_delay_1;
    tap_tdoBuffer_delay_3 <= tap_tdoBuffer_delay_2;
    tap_tdoShifter <= tap_tdoBuffer_delay_3;
    if(logic_jtagLogic_dtmcs_logic_ctrl_enable) begin
      if(logic_jtagLogic_dtmcs_logic_ctrl_capture) begin
        logic_jtagLogic_dtmcs_logic_store <= logic_jtagLogic_dtmcs_captureData;
      end
      if(logic_jtagLogic_dtmcs_logic_ctrl_shift) begin
        logic_jtagLogic_dtmcs_logic_store <= ({logic_jtagLogic_dtmcs_logic_ctrl_tdi,logic_jtagLogic_dtmcs_logic_store} >>> 1'd1);
      end
    end
    if(logic_jtagLogic_dmi_logic_ctrl_enable) begin
      if(logic_jtagLogic_dmi_logic_ctrl_capture) begin
        logic_jtagLogic_dmi_logic_store <= {logic_jtagLogic_dmi_captureData_padding,{logic_jtagLogic_dmi_captureData_data,logic_jtagLogic_dmi_captureData_op}};
      end
      if(logic_jtagLogic_dmi_logic_ctrl_shift) begin
        logic_jtagLogic_dmi_logic_store <= ({logic_jtagLogic_dmi_logic_ctrl_tdi,logic_jtagLogic_dmi_logic_store} >>> 1'd1);
      end
    end
    if(logic_jtagLogic_dmiCmd_valid) begin
      logic_jtagLogic_pending <= 1'b1;
    end
    if(logic_jtagLogic_dmiRsp_valid) begin
      logic_jtagLogic_pending <= 1'b0;
    end
    if(logic_jtagLogic_trigger_dmiHardReset) begin
      logic_jtagLogic_pending <= 1'b0;
    end
    if(logic_jtagLogic_dmiRsp_valid) begin
      logic_jtagLogic_rspLogic_buffer <= logic_jtagLogic_dmiRsp_payload_data;
    end
    logic_jtagLogic_dmiStat_value <= logic_jtagLogic_dmiStat_value_aheadValue;
  end

  always @(posedge io_systemClk) begin
    if(debugCd_logic_outputReset) begin
      logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rValid <= 1'b0;
    end else begin
      if(logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_ready) begin
        logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rValid <= logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_valid;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_fire) begin
      logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_write <= logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_write;
      logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_data <= logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_data;
      logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_rData_address <= logic_jtagLogic_dmiCmd_ccToggle_io_output_toStream_payload_address;
    end
  end


endmodule

module BufferCC_65 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_memoryClk,
  input  wire          system_riscvJtag_debug_systemReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk or posedge system_riscvJtag_debug_systemReset) begin
    if(system_riscvJtag_debug_systemReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_64 replaced by BufferCC_60

//StreamFifo_16 replaced by StreamFifo_15

module StreamFifo_15 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [3:0]    io_push_payload,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [3:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [5:0]    io_occupancy,
  output wire [5:0]    io_availability,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg        [3:0]    logic_ram_spinal_port1;
  wire       [3:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [5:0]    logic_ptr_push;
  reg        [5:0]    logic_ptr_pop;
  wire       [5:0]    logic_ptr_occupancy;
  wire       [5:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [4:0]    logic_push_onRam_write_payload_address;
  wire       [3:0]    logic_push_onRam_write_payload_data;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [4:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [4:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [4:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [4:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [3:0]    logic_pop_sync_readPort_rsp;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [5:0]    logic_pop_sync_popReg;
  reg [3:0] logic_ram [0:31];

  assign _zz_logic_ram_port = logic_push_onRam_write_payload_data;
  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge io_systemClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 6'h20) == 6'h0);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[4:0];
  assign logic_push_onRam_write_payload_data = io_push_payload;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[4:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign logic_pop_sync_readPort_rsp = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload = logic_pop_sync_readPort_rsp;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload = logic_pop_sync_readArbitation_translated_payload;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (6'h20 - logic_ptr_occupancy);
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      logic_ptr_push <= 6'h0;
      logic_ptr_pop <= 6'h0;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 6'h0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 6'h01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 6'h01);
      end
      if(io_flush) begin
        logic_ptr_push <= 6'h0;
        logic_ptr_pop <= 6'h0;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 6'h0;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

//BufferCC_63 replaced by BufferCC_60

//BufferCC_62 replaced by BufferCC_60

//BufferCC_61 replaced by BufferCC_60

module BufferCC_60 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

module BufferCC_59 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          ddrCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk or posedge ddrCd_logic_outputReset) begin
    if(ddrCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_58 replaced by BufferCC_39

module BufferCC_57 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_memoryClk,
  input  wire          debugCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk or posedge debugCd_logic_outputReset) begin
    if(debugCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_56 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_systemClk,
  input  wire          io_asyncReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk or posedge io_asyncReset) begin
    if(io_asyncReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module DebugModule (
  input  wire          io_ctrl_cmd_valid,
  output wire          io_ctrl_cmd_ready,
  input  wire          io_ctrl_cmd_payload_write,
  input  wire [31:0]   io_ctrl_cmd_payload_data,
  input  wire [6:0]    io_ctrl_cmd_payload_address,
  output wire          io_ctrl_rsp_valid,
  output wire          io_ctrl_rsp_payload_error,
  output wire [31:0]   io_ctrl_rsp_payload_data,
  output wire          io_ndmreset,
  input  wire          io_harts_0_halted,
  input  wire          io_harts_0_running,
  input  wire          io_harts_0_unavailable,
  input  wire          io_harts_0_exception,
  input  wire          io_harts_0_commit,
  input  wire          io_harts_0_ebreak,
  input  wire          io_harts_0_redo,
  input  wire          io_harts_0_regSuccess,
  output wire          io_harts_0_ackReset,
  input  wire          io_harts_0_haveReset,
  output reg           io_harts_0_resume_cmd_valid,
  input  wire          io_harts_0_resume_rsp_valid,
  output wire          io_harts_0_haltReq,
  output wire          io_harts_0_dmToHart_valid,
  output wire [1:0]    io_harts_0_dmToHart_payload_op,
  output wire [4:0]    io_harts_0_dmToHart_payload_address,
  output wire [31:0]   io_harts_0_dmToHart_payload_data,
  output wire [2:0]    io_harts_0_dmToHart_payload_size,
  input  wire          io_harts_0_hartToDm_valid,
  input  wire [3:0]    io_harts_0_hartToDm_payload_address,
  input  wire [31:0]   io_harts_0_hartToDm_payload_data,
  input  wire          io_harts_1_halted,
  input  wire          io_harts_1_running,
  input  wire          io_harts_1_unavailable,
  input  wire          io_harts_1_exception,
  input  wire          io_harts_1_commit,
  input  wire          io_harts_1_ebreak,
  input  wire          io_harts_1_redo,
  input  wire          io_harts_1_regSuccess,
  output wire          io_harts_1_ackReset,
  input  wire          io_harts_1_haveReset,
  output reg           io_harts_1_resume_cmd_valid,
  input  wire          io_harts_1_resume_rsp_valid,
  output wire          io_harts_1_haltReq,
  output wire          io_harts_1_dmToHart_valid,
  output wire [1:0]    io_harts_1_dmToHart_payload_op,
  output wire [4:0]    io_harts_1_dmToHart_payload_address,
  output wire [31:0]   io_harts_1_dmToHart_payload_data,
  output wire [2:0]    io_harts_1_dmToHart_payload_size,
  input  wire          io_harts_1_hartToDm_valid,
  input  wire [3:0]    io_harts_1_hartToDm_payload_address,
  input  wire [31:0]   io_harts_1_hartToDm_payload_data,
  input  wire          io_systemClk,
  input  wire          debugCd_logic_outputReset
);
  localparam DebugDmToHartOp_DATA = 2'd0;
  localparam DebugDmToHartOp_EXECUTE = 2'd1;
  localparam DebugDmToHartOp_REG_WRITE = 2'd2;
  localparam DebugDmToHartOp_REG_READ = 2'd3;
  localparam DebugModuleCmdErr_NONE = 3'd0;
  localparam DebugModuleCmdErr_BUSY = 3'd1;
  localparam DebugModuleCmdErr_NOT_SUPPORTED = 3'd2;
  localparam DebugModuleCmdErr_EXCEPTION = 3'd3;
  localparam DebugModuleCmdErr_HALT_RESUME = 3'd4;
  localparam DebugModuleCmdErr_BUS_1 = 3'd5;
  localparam DebugModuleCmdErr_OTHER = 3'd6;
  localparam logic_command_enumDef_BOOT = 4'd0;
  localparam logic_command_enumDef_IDLE = 4'd1;
  localparam logic_command_enumDef_DECODE = 4'd2;
  localparam logic_command_enumDef_READ_INT_REG = 4'd3;
  localparam logic_command_enumDef_WRITE_INT_REG = 4'd4;
  localparam logic_command_enumDef_WAIT_DONE = 4'd5;
  localparam logic_command_enumDef_POST_EXEC = 4'd6;
  localparam logic_command_enumDef_POST_EXEC_WAIT = 4'd7;
  localparam logic_command_enumDef_READ_FPU_REG = 4'd8;
  localparam logic_command_enumDef_WRITE_FPU_REG = 4'd9;

  wire       [31:0]   logic_progbufX_mem_spinal_port1;
  wire       [31:0]   logic_dataX_readMem_spinal_port1;
  wire       [0:0]    _zz_logic_dmcontrol_haltSet;
  wire       [0:0]    _zz_logic_dmcontrol_haltClear;
  wire       [0:0]    _zz_logic_dmcontrol_resumeReq;
  wire       [0:0]    _zz_logic_dmcontrol_ackhavereset;
  reg        [1:0]    _zz_logic_dmcontrol_hartSelAarsizeLimit;
  wire       [0:0]    _zz_logic_dmcontrol_hartSelAarsizeLimit_1;
  reg        [1:0]    _zz_logic_dmcontrol_hartSelAarsizeLimitF;
  wire       [0:0]    _zz_logic_dmcontrol_hartSelAarsizeLimitF_1;
  reg                 _zz_logic_selected_running;
  reg                 _zz_logic_selected_halted;
  reg                 _zz_logic_selected_commit;
  reg                 _zz_logic_selected_regSuccess;
  reg                 _zz_logic_selected_exception;
  reg                 _zz_logic_selected_ebreak;
  reg                 _zz_logic_selected_redo;
  wire       [14:0]   _zz_when_DebugModule_l143;
  wire       [0:0]    _zz_logic_progbufX_mem_port;
  wire       [0:0]    _zz_logic_dataX_readMem_port;
  wire       [6:0]    _zz_logic_dataX_cmdAddress;
  wire       [0:0]    _zz_logic_abstractAuto_trigger;
  wire       [2:0]    _zz_logic_command_access_notSupported;
  wire       [1:0]    _zz_logic_command_access_notSupported_1;
  reg                 _zz_when_DebugModule_l276;
  wire       [0:0]    _zz_when_DebugModule_l276_1;
  wire       [31:0]   _zz_logic_toHarts_payload_data;
  wire       [19:0]   _zz_logic_toHarts_payload_data_1;
  wire       [31:0]   _zz_logic_toHarts_payload_data_2;
  wire       [11:0]   _zz_logic_toHarts_payload_data_3;
  reg                 _zz_1;
  wire                factory_readErrorFlag;
  wire                factory_writeErrorFlag;
  wire                factory_cmdToRsp_valid;
  reg                 factory_cmdToRsp_payload_error;
  reg        [31:0]   factory_cmdToRsp_payload_data;
  reg                 factory_rspBuffer_valid;
  reg                 factory_rspBuffer_payload_error;
  reg        [31:0]   factory_rspBuffer_payload_data;
  wire                factory_askWrite;
  wire                factory_askRead;
  wire                factory_doWrite;
  wire                factory_doRead;
  wire                io_ctrl_cmd_fire;
  reg                 dmactive;
  reg                 logic_dmcontrol_ndmreset;
  wire       [9:0]    logic_dmcontrol_hartSelLoNew;
  wire       [9:0]    logic_dmcontrol_hartSelHiNew;
  wire       [19:0]   logic_dmcontrol_hartSelNew;
  reg        [9:0]    logic_dmcontrol_hartSelLo;
  reg        [9:0]    logic_dmcontrol_hartSelHi;
  wire       [19:0]   logic_dmcontrol_hartSel;
  reg                 logic_dmcontrol_haltSet;
  reg                 when_BusSlaveFactory_l377;
  wire                when_BusSlaveFactory_l379;
  reg                 logic_dmcontrol_haltClear;
  reg                 when_BusSlaveFactory_l391;
  wire                when_BusSlaveFactory_l393;
  reg                 logic_dmcontrol_resumeReq;
  reg                 when_BusSlaveFactory_l377_1;
  wire                when_BusSlaveFactory_l379_1;
  reg                 logic_dmcontrol_ackhavereset;
  reg                 when_BusSlaveFactory_l377_2;
  wire                when_BusSlaveFactory_l379_2;
  wire       [1:0]    logic_dmcontrol_hartSelAarsizeLimit;
  wire       [1:0]    logic_dmcontrol_hartSelAarsizeLimitF;
  reg                 logic_dmcontrol_harts_0_haltReq;
  wire                when_DebugModule_l102;
  reg                 logic_dmcontrol_harts_1_haltReq;
  wire                when_DebugModule_l102_1;
  reg                 logic_toHarts_valid;
  reg        [1:0]    logic_toHarts_payload_op;
  reg        [4:0]    logic_toHarts_payload_address;
  reg        [31:0]   logic_toHarts_payload_data;
  reg        [2:0]    logic_toHarts_payload_size;
  wire                logic_fromHarts_valid;
  wire       [3:0]    logic_fromHarts_payload_address;
  wire       [31:0]   logic_fromHarts_payload_data;
  wire       [35:0]   _zz_logic_fromHarts_payload_address;
  wire                logic_harts_0_sel;
  reg                 _zz_logic_harts_0_resumeReady;
  reg                 _zz_logic_harts_0_resumeReady_1;
  wire                logic_harts_0_resumeReady;
  wire                logic_toHarts_takeWhen_valid;
  wire       [1:0]    logic_toHarts_takeWhen_payload_op;
  wire       [4:0]    logic_toHarts_takeWhen_payload_address;
  wire       [31:0]   logic_toHarts_takeWhen_payload_data;
  wire       [2:0]    logic_toHarts_takeWhen_payload_size;
  reg                 _zz_io_harts_0_ackReset;
  wire                logic_harts_1_sel;
  reg                 _zz_logic_harts_1_resumeReady;
  reg                 _zz_logic_harts_1_resumeReady_1;
  wire                logic_harts_1_resumeReady;
  wire                logic_toHarts_takeWhen_valid_1;
  wire       [1:0]    logic_toHarts_takeWhen_payload_op_1;
  wire       [4:0]    logic_toHarts_takeWhen_payload_address_1;
  wire       [31:0]   logic_toHarts_takeWhen_payload_data_1;
  wire       [2:0]    logic_toHarts_takeWhen_payload_size_1;
  reg                 _zz_io_harts_1_ackReset;
  reg        [0:0]    logic_selected_hart;
  wire                logic_selected_running;
  wire                logic_selected_halted;
  wire                logic_selected_commit;
  wire                logic_selected_regSuccess;
  wire                logic_selected_exception;
  wire                logic_selected_ebreak;
  wire                logic_selected_redo;
  reg        [31:0]   logic_haltsum_value;
  wire                when_DebugModule_l143;
  wire       [3:0]    logic_dmstatus_version;
  wire                logic_dmstatus_authenticated;
  wire                logic_dmstatus_anyHalted;
  wire                logic_dmstatus_allHalted;
  wire                logic_dmstatus_anyRunning;
  wire                logic_dmstatus_allRunning;
  wire                logic_dmstatus_anyUnavail;
  wire                logic_dmstatus_allUnavail;
  wire                logic_dmstatus_anyNonExistent;
  wire                logic_dmstatus_anyResumeAck;
  wire                logic_dmstatus_allResumeAck;
  wire                logic_dmstatus_anyHaveReset;
  wire                logic_dmstatus_allHaveReset;
  wire                logic_dmstatus_impebreak;
  wire       [3:0]    logic_hartInfo_dataaddr;
  wire       [3:0]    logic_hartInfo_datasize;
  wire                logic_hartInfo_dataaccess;
  wire       [3:0]    logic_hartInfo_nscratch;
  wire       [2:0]    logic_sbcs_sbversion;
  wire       [2:0]    logic_sbcs_sbaccess;
  wire                logic_progbufX_trigged;
  reg                 logic_dataX_trigged;
  wire       [0:0]    logic_dataX_cmdAddress;
  wire                when_DebugModule_l205;
  wire       [0:0]    _zz_factory_cmdToRsp_payload_data;
  wire       [3:0]    logic_abstractcs_dataCount;
  reg        [2:0]    logic_abstractcs_cmdErr;
  reg                 when_BusSlaveFactory_l341;
  wire       [2:0]    _zz_logic_abstractcs_cmdErr;
  reg                 logic_abstractcs_busy;
  wire       [4:0]    logic_abstractcs_progBufSize;
  wire                logic_abstractcs_noError;
  reg        [1:0]    logic_abstractAuto_autoexecdata;
  reg        [1:0]    logic_abstractAuto_autoexecProgbuf;
  wire                logic_abstractAuto_trigger;
  wire                logic_command_wantExit;
  reg                 logic_command_wantStart;
  wire                logic_command_wantKill;
  reg        [0:0]    logic_command_executionCounter;
  reg                 logic_command_commandRequest;
  reg        [31:0]   logic_command_data;
  wire       [15:0]   logic_command_access_args_regno;
  wire                logic_command_access_args_write;
  wire                logic_command_access_args_transfer;
  wire                logic_command_access_args_postExec;
  wire                logic_command_access_args_aarpostincrement;
  wire       [2:0]    logic_command_access_args_aarsize;
  wire       [31:0]   _zz_logic_command_access_args_regno;
  wire                logic_command_access_transferFloat;
  wire                logic_command_access_notSupported;
  wire                logic_command_request;
  wire                when_DebugModule_l260;
  wire                when_DebugModule_l263;
  wire                when_DebugModule_l266;
  reg        [3:0]    logic_command_stateReg;
  reg        [3:0]    logic_command_stateNext;
  wire                when_DebugModule_l275;
  wire                when_DebugModule_l276;
  wire       [7:0]    switch_DebugModule_l287;
  wire                when_DebugModule_l296;
  wire                when_DebugModule_l350;
  wire                when_DebugModule_l366;
  wire                when_DebugModule_l370;
  wire                when_StateMachine_l253;
  `ifndef SYNTHESIS
  reg [71:0] io_harts_0_dmToHart_payload_op_string;
  reg [71:0] io_harts_1_dmToHart_payload_op_string;
  reg [71:0] logic_toHarts_payload_op_string;
  reg [71:0] logic_toHarts_takeWhen_payload_op_string;
  reg [71:0] logic_toHarts_takeWhen_payload_op_1_string;
  reg [103:0] logic_abstractcs_cmdErr_string;
  reg [103:0] _zz_logic_abstractcs_cmdErr_string;
  reg [111:0] logic_command_stateReg_string;
  reg [111:0] logic_command_stateNext_string;
  `endif

  (* ram_style = "distributed" *) reg [31:0] logic_progbufX_mem [0:1];
  (* ram_style = "distributed" *) reg [31:0] logic_dataX_readMem [0:1];

  assign _zz_logic_dmcontrol_haltSet = 1'b1;
  assign _zz_logic_dmcontrol_haltClear = 1'b1;
  assign _zz_logic_dmcontrol_resumeReq = 1'b1;
  assign _zz_logic_dmcontrol_ackhavereset = 1'b1;
  assign _zz_logic_dmcontrol_hartSelAarsizeLimit_1 = logic_dmcontrol_hartSel[0:0];
  assign _zz_logic_dmcontrol_hartSelAarsizeLimitF_1 = logic_dmcontrol_hartSel[0:0];
  assign _zz_when_DebugModule_l143 = (logic_dmcontrol_hartSel >>> 3'd5);
  assign _zz_logic_progbufX_mem_port = io_ctrl_cmd_payload_address[0:0];
  assign _zz_logic_dataX_readMem_port = logic_fromHarts_payload_address[0:0];
  assign _zz_logic_dataX_cmdAddress = (io_ctrl_cmd_payload_address - 7'h04);
  assign _zz_logic_abstractAuto_trigger = io_ctrl_cmd_payload_address[0:0];
  assign _zz_logic_command_access_notSupported_1 = (logic_command_access_transferFloat ? logic_dmcontrol_hartSelAarsizeLimitF : logic_dmcontrol_hartSelAarsizeLimit);
  assign _zz_logic_command_access_notSupported = {1'd0, _zz_logic_command_access_notSupported_1};
  assign _zz_when_DebugModule_l276_1 = logic_dmcontrol_hartSel[0:0];
  assign _zz_logic_toHarts_payload_data_1 = ({15'd0,logic_command_access_args_regno[4 : 0]} <<< 4'd15);
  assign _zz_logic_toHarts_payload_data = {12'd0, _zz_logic_toHarts_payload_data_1};
  assign _zz_logic_toHarts_payload_data_3 = ({7'd0,logic_command_access_args_regno[4 : 0]} <<< 3'd7);
  assign _zz_logic_toHarts_payload_data_2 = {20'd0, _zz_logic_toHarts_payload_data_3};
  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      logic_progbufX_mem[_zz_logic_progbufX_mem_port] <= io_ctrl_cmd_payload_data;
    end
  end

  assign logic_progbufX_mem_spinal_port1 = logic_progbufX_mem[logic_command_executionCounter];
  always @(posedge io_systemClk) begin
    if(logic_fromHarts_valid) begin
      logic_dataX_readMem[_zz_logic_dataX_readMem_port] <= logic_fromHarts_payload_data;
    end
  end

  assign logic_dataX_readMem_spinal_port1 = logic_dataX_readMem[_zz_factory_cmdToRsp_payload_data];
  always @(*) begin
    case(_zz_logic_dmcontrol_hartSelAarsizeLimit_1)
      1'b0 : _zz_logic_dmcontrol_hartSelAarsizeLimit = 2'b10;
      default : _zz_logic_dmcontrol_hartSelAarsizeLimit = 2'b10;
    endcase
  end

  always @(*) begin
    case(_zz_logic_dmcontrol_hartSelAarsizeLimitF_1)
      1'b0 : _zz_logic_dmcontrol_hartSelAarsizeLimitF = 2'b11;
      default : _zz_logic_dmcontrol_hartSelAarsizeLimitF = 2'b11;
    endcase
  end

  always @(*) begin
    case(logic_selected_hart)
      1'b0 : begin
        _zz_logic_selected_running = io_harts_0_running;
        _zz_logic_selected_halted = io_harts_0_halted;
        _zz_logic_selected_commit = io_harts_0_commit;
        _zz_logic_selected_regSuccess = io_harts_0_regSuccess;
        _zz_logic_selected_exception = io_harts_0_exception;
        _zz_logic_selected_ebreak = io_harts_0_ebreak;
        _zz_logic_selected_redo = io_harts_0_redo;
      end
      default : begin
        _zz_logic_selected_running = io_harts_1_running;
        _zz_logic_selected_halted = io_harts_1_halted;
        _zz_logic_selected_commit = io_harts_1_commit;
        _zz_logic_selected_regSuccess = io_harts_1_regSuccess;
        _zz_logic_selected_exception = io_harts_1_exception;
        _zz_logic_selected_ebreak = io_harts_1_ebreak;
        _zz_logic_selected_redo = io_harts_1_redo;
      end
    endcase
  end

  always @(*) begin
    case(_zz_when_DebugModule_l276_1)
      1'b0 : _zz_when_DebugModule_l276 = io_harts_0_halted;
      default : _zz_when_DebugModule_l276 = io_harts_1_halted;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_harts_0_dmToHart_payload_op)
      DebugDmToHartOp_DATA : io_harts_0_dmToHart_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : io_harts_0_dmToHart_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : io_harts_0_dmToHart_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : io_harts_0_dmToHart_payload_op_string = "REG_READ ";
      default : io_harts_0_dmToHart_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(io_harts_1_dmToHart_payload_op)
      DebugDmToHartOp_DATA : io_harts_1_dmToHart_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : io_harts_1_dmToHart_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : io_harts_1_dmToHart_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : io_harts_1_dmToHart_payload_op_string = "REG_READ ";
      default : io_harts_1_dmToHart_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(logic_toHarts_payload_op)
      DebugDmToHartOp_DATA : logic_toHarts_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : logic_toHarts_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : logic_toHarts_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : logic_toHarts_payload_op_string = "REG_READ ";
      default : logic_toHarts_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(logic_toHarts_takeWhen_payload_op)
      DebugDmToHartOp_DATA : logic_toHarts_takeWhen_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : logic_toHarts_takeWhen_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : logic_toHarts_takeWhen_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : logic_toHarts_takeWhen_payload_op_string = "REG_READ ";
      default : logic_toHarts_takeWhen_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(logic_toHarts_takeWhen_payload_op_1)
      DebugDmToHartOp_DATA : logic_toHarts_takeWhen_payload_op_1_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : logic_toHarts_takeWhen_payload_op_1_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : logic_toHarts_takeWhen_payload_op_1_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : logic_toHarts_takeWhen_payload_op_1_string = "REG_READ ";
      default : logic_toHarts_takeWhen_payload_op_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(logic_abstractcs_cmdErr)
      DebugModuleCmdErr_NONE : logic_abstractcs_cmdErr_string = "NONE         ";
      DebugModuleCmdErr_BUSY : logic_abstractcs_cmdErr_string = "BUSY         ";
      DebugModuleCmdErr_NOT_SUPPORTED : logic_abstractcs_cmdErr_string = "NOT_SUPPORTED";
      DebugModuleCmdErr_EXCEPTION : logic_abstractcs_cmdErr_string = "EXCEPTION    ";
      DebugModuleCmdErr_HALT_RESUME : logic_abstractcs_cmdErr_string = "HALT_RESUME  ";
      DebugModuleCmdErr_BUS_1 : logic_abstractcs_cmdErr_string = "BUS_1        ";
      DebugModuleCmdErr_OTHER : logic_abstractcs_cmdErr_string = "OTHER        ";
      default : logic_abstractcs_cmdErr_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(_zz_logic_abstractcs_cmdErr)
      DebugModuleCmdErr_NONE : _zz_logic_abstractcs_cmdErr_string = "NONE         ";
      DebugModuleCmdErr_BUSY : _zz_logic_abstractcs_cmdErr_string = "BUSY         ";
      DebugModuleCmdErr_NOT_SUPPORTED : _zz_logic_abstractcs_cmdErr_string = "NOT_SUPPORTED";
      DebugModuleCmdErr_EXCEPTION : _zz_logic_abstractcs_cmdErr_string = "EXCEPTION    ";
      DebugModuleCmdErr_HALT_RESUME : _zz_logic_abstractcs_cmdErr_string = "HALT_RESUME  ";
      DebugModuleCmdErr_BUS_1 : _zz_logic_abstractcs_cmdErr_string = "BUS_1        ";
      DebugModuleCmdErr_OTHER : _zz_logic_abstractcs_cmdErr_string = "OTHER        ";
      default : _zz_logic_abstractcs_cmdErr_string = "?????????????";
    endcase
  end
  always @(*) begin
    case(logic_command_stateReg)
      logic_command_enumDef_BOOT : logic_command_stateReg_string = "BOOT          ";
      logic_command_enumDef_IDLE : logic_command_stateReg_string = "IDLE          ";
      logic_command_enumDef_DECODE : logic_command_stateReg_string = "DECODE        ";
      logic_command_enumDef_READ_INT_REG : logic_command_stateReg_string = "READ_INT_REG  ";
      logic_command_enumDef_WRITE_INT_REG : logic_command_stateReg_string = "WRITE_INT_REG ";
      logic_command_enumDef_WAIT_DONE : logic_command_stateReg_string = "WAIT_DONE     ";
      logic_command_enumDef_POST_EXEC : logic_command_stateReg_string = "POST_EXEC     ";
      logic_command_enumDef_POST_EXEC_WAIT : logic_command_stateReg_string = "POST_EXEC_WAIT";
      logic_command_enumDef_READ_FPU_REG : logic_command_stateReg_string = "READ_FPU_REG  ";
      logic_command_enumDef_WRITE_FPU_REG : logic_command_stateReg_string = "WRITE_FPU_REG ";
      default : logic_command_stateReg_string = "??????????????";
    endcase
  end
  always @(*) begin
    case(logic_command_stateNext)
      logic_command_enumDef_BOOT : logic_command_stateNext_string = "BOOT          ";
      logic_command_enumDef_IDLE : logic_command_stateNext_string = "IDLE          ";
      logic_command_enumDef_DECODE : logic_command_stateNext_string = "DECODE        ";
      logic_command_enumDef_READ_INT_REG : logic_command_stateNext_string = "READ_INT_REG  ";
      logic_command_enumDef_WRITE_INT_REG : logic_command_stateNext_string = "WRITE_INT_REG ";
      logic_command_enumDef_WAIT_DONE : logic_command_stateNext_string = "WAIT_DONE     ";
      logic_command_enumDef_POST_EXEC : logic_command_stateNext_string = "POST_EXEC     ";
      logic_command_enumDef_POST_EXEC_WAIT : logic_command_stateNext_string = "POST_EXEC_WAIT";
      logic_command_enumDef_READ_FPU_REG : logic_command_stateNext_string = "READ_FPU_REG  ";
      logic_command_enumDef_WRITE_FPU_REG : logic_command_stateNext_string = "WRITE_FPU_REG ";
      default : logic_command_stateNext_string = "??????????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_progbufX_trigged) begin
      _zz_1 = 1'b1;
    end
  end

  assign factory_readErrorFlag = 1'b0;
  assign factory_writeErrorFlag = 1'b0;
  assign io_ctrl_cmd_ready = 1'b1;
  assign factory_askWrite = (io_ctrl_cmd_valid && io_ctrl_cmd_payload_write);
  assign factory_askRead = (io_ctrl_cmd_valid && (! io_ctrl_cmd_payload_write));
  assign factory_doWrite = (factory_askWrite && io_ctrl_cmd_ready);
  assign factory_doRead = (factory_askRead && io_ctrl_cmd_ready);
  assign io_ctrl_rsp_valid = factory_rspBuffer_valid;
  assign io_ctrl_rsp_payload_error = factory_rspBuffer_payload_error;
  assign io_ctrl_rsp_payload_data = factory_rspBuffer_payload_data;
  assign io_ctrl_cmd_fire = (io_ctrl_cmd_valid && io_ctrl_cmd_ready);
  assign factory_cmdToRsp_valid = io_ctrl_cmd_fire;
  always @(*) begin
    factory_cmdToRsp_payload_error = 1'b0;
    if(logic_progbufX_trigged) begin
      factory_cmdToRsp_payload_error = 1'b0;
    end
    if(when_DebugModule_l205) begin
      factory_cmdToRsp_payload_error = 1'b0;
    end
    case(io_ctrl_cmd_payload_address)
      7'h10 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      7'h40 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      7'h11 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      7'h12 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      7'h38 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      7'h16 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      7'h18 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      7'h17 : begin
        factory_cmdToRsp_payload_error = 1'b0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    factory_cmdToRsp_payload_data = 32'h0;
    if(when_DebugModule_l205) begin
      factory_cmdToRsp_payload_data = logic_dataX_readMem_spinal_port1;
    end
    case(io_ctrl_cmd_payload_address)
      7'h10 : begin
        factory_cmdToRsp_payload_data[0 : 0] = dmactive;
        factory_cmdToRsp_payload_data[1 : 1] = logic_dmcontrol_ndmreset;
        factory_cmdToRsp_payload_data[25 : 16] = logic_dmcontrol_hartSelLo;
        factory_cmdToRsp_payload_data[15 : 6] = logic_dmcontrol_hartSelHi;
      end
      7'h40 : begin
        factory_cmdToRsp_payload_data[31 : 0] = logic_haltsum_value;
      end
      7'h11 : begin
        factory_cmdToRsp_payload_data[3 : 0] = logic_dmstatus_version;
        factory_cmdToRsp_payload_data[7 : 7] = logic_dmstatus_authenticated;
        factory_cmdToRsp_payload_data[8 : 8] = logic_dmstatus_anyHalted;
        factory_cmdToRsp_payload_data[9 : 9] = logic_dmstatus_allHalted;
        factory_cmdToRsp_payload_data[10 : 10] = logic_dmstatus_anyRunning;
        factory_cmdToRsp_payload_data[11 : 11] = logic_dmstatus_allRunning;
        factory_cmdToRsp_payload_data[12 : 12] = logic_dmstatus_anyUnavail;
        factory_cmdToRsp_payload_data[13 : 13] = logic_dmstatus_allUnavail;
        factory_cmdToRsp_payload_data[14 : 14] = logic_dmstatus_anyNonExistent;
        factory_cmdToRsp_payload_data[15 : 15] = logic_dmstatus_anyNonExistent;
        factory_cmdToRsp_payload_data[16 : 16] = logic_dmstatus_anyResumeAck;
        factory_cmdToRsp_payload_data[17 : 17] = logic_dmstatus_allResumeAck;
        factory_cmdToRsp_payload_data[18 : 18] = logic_dmstatus_anyHaveReset;
        factory_cmdToRsp_payload_data[19 : 19] = logic_dmstatus_allHaveReset;
        factory_cmdToRsp_payload_data[22 : 22] = logic_dmstatus_impebreak;
      end
      7'h12 : begin
        factory_cmdToRsp_payload_data[3 : 0] = logic_hartInfo_dataaddr;
        factory_cmdToRsp_payload_data[15 : 12] = logic_hartInfo_datasize;
        factory_cmdToRsp_payload_data[16 : 16] = logic_hartInfo_dataaccess;
        factory_cmdToRsp_payload_data[23 : 20] = logic_hartInfo_nscratch;
      end
      7'h38 : begin
        factory_cmdToRsp_payload_data[31 : 29] = logic_sbcs_sbversion;
        factory_cmdToRsp_payload_data[19 : 17] = logic_sbcs_sbaccess;
      end
      7'h16 : begin
        factory_cmdToRsp_payload_data[3 : 0] = logic_abstractcs_dataCount;
        factory_cmdToRsp_payload_data[10 : 8] = logic_abstractcs_cmdErr;
        factory_cmdToRsp_payload_data[12 : 12] = logic_abstractcs_busy;
        factory_cmdToRsp_payload_data[28 : 24] = logic_abstractcs_progBufSize;
      end
      7'h18 : begin
        factory_cmdToRsp_payload_data[1 : 0] = logic_abstractAuto_autoexecdata;
        factory_cmdToRsp_payload_data[17 : 16] = logic_abstractAuto_autoexecProgbuf;
      end
      default : begin
      end
    endcase
  end

  assign logic_dmcontrol_hartSelNew = {logic_dmcontrol_hartSelHiNew,logic_dmcontrol_hartSelLoNew};
  assign logic_dmcontrol_hartSel = {logic_dmcontrol_hartSelHi,logic_dmcontrol_hartSelLo};
  always @(*) begin
    logic_dmcontrol_haltSet = 1'b0;
    if(when_BusSlaveFactory_l377) begin
      if(when_BusSlaveFactory_l379) begin
        logic_dmcontrol_haltSet = _zz_logic_dmcontrol_haltSet[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377 = 1'b0;
    case(io_ctrl_cmd_payload_address)
      7'h10 : begin
        if(factory_doWrite) begin
          when_BusSlaveFactory_l377 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379 = io_ctrl_cmd_payload_data[31];
  always @(*) begin
    logic_dmcontrol_haltClear = 1'b0;
    if(when_BusSlaveFactory_l391) begin
      if(when_BusSlaveFactory_l393) begin
        logic_dmcontrol_haltClear = _zz_logic_dmcontrol_haltClear[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l391 = 1'b0;
    case(io_ctrl_cmd_payload_address)
      7'h10 : begin
        if(factory_doWrite) begin
          when_BusSlaveFactory_l391 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l393 = (! io_ctrl_cmd_payload_data[31]);
  always @(*) begin
    logic_dmcontrol_resumeReq = 1'b0;
    if(when_BusSlaveFactory_l377_1) begin
      if(when_BusSlaveFactory_l379_1) begin
        logic_dmcontrol_resumeReq = _zz_logic_dmcontrol_resumeReq[0];
      end
    end
    if(logic_dmcontrol_haltSet) begin
      logic_dmcontrol_resumeReq = 1'b0;
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_1 = 1'b0;
    case(io_ctrl_cmd_payload_address)
      7'h10 : begin
        if(factory_doWrite) begin
          when_BusSlaveFactory_l377_1 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_1 = io_ctrl_cmd_payload_data[30];
  always @(*) begin
    logic_dmcontrol_ackhavereset = 1'b0;
    if(when_BusSlaveFactory_l377_2) begin
      if(when_BusSlaveFactory_l379_2) begin
        logic_dmcontrol_ackhavereset = _zz_logic_dmcontrol_ackhavereset[0];
      end
    end
  end

  always @(*) begin
    when_BusSlaveFactory_l377_2 = 1'b0;
    case(io_ctrl_cmd_payload_address)
      7'h10 : begin
        if(factory_doWrite) begin
          when_BusSlaveFactory_l377_2 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_BusSlaveFactory_l379_2 = io_ctrl_cmd_payload_data[28];
  assign logic_dmcontrol_hartSelAarsizeLimit = _zz_logic_dmcontrol_hartSelAarsizeLimit;
  assign logic_dmcontrol_hartSelAarsizeLimitF = _zz_logic_dmcontrol_hartSelAarsizeLimitF;
  assign io_harts_0_haltReq = logic_dmcontrol_harts_0_haltReq;
  always @(*) begin
    io_harts_0_resume_cmd_valid = 1'b0;
    if(when_DebugModule_l102) begin
      io_harts_0_resume_cmd_valid = logic_dmcontrol_resumeReq;
    end
  end

  assign when_DebugModule_l102 = (logic_dmcontrol_hartSelNew == 20'h0);
  assign io_harts_1_haltReq = logic_dmcontrol_harts_1_haltReq;
  always @(*) begin
    io_harts_1_resume_cmd_valid = 1'b0;
    if(when_DebugModule_l102_1) begin
      io_harts_1_resume_cmd_valid = logic_dmcontrol_resumeReq;
    end
  end

  assign when_DebugModule_l102_1 = (logic_dmcontrol_hartSelNew == 20'h00001);
  assign io_ndmreset = logic_dmcontrol_ndmreset;
  always @(*) begin
    logic_toHarts_valid = 1'b0;
    if(when_DebugModule_l205) begin
      if(io_ctrl_cmd_payload_write) begin
        logic_toHarts_valid = 1'b1;
      end
    end
    if(logic_abstractcs_busy) begin
      logic_toHarts_valid = 1'b0;
    end
    case(logic_command_stateReg)
      logic_command_enumDef_IDLE : begin
      end
      logic_command_enumDef_DECODE : begin
      end
      logic_command_enumDef_READ_INT_REG : begin
        logic_toHarts_valid = 1'b1;
      end
      logic_command_enumDef_WRITE_INT_REG : begin
        logic_toHarts_valid = 1'b1;
      end
      logic_command_enumDef_WAIT_DONE : begin
      end
      logic_command_enumDef_POST_EXEC : begin
        logic_toHarts_valid = 1'b1;
      end
      logic_command_enumDef_POST_EXEC_WAIT : begin
      end
      logic_command_enumDef_READ_FPU_REG : begin
        logic_toHarts_valid = 1'b1;
      end
      logic_command_enumDef_WRITE_FPU_REG : begin
        logic_toHarts_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    logic_toHarts_payload_op = (2'bxx);
    if(when_DebugModule_l205) begin
      logic_toHarts_payload_op = DebugDmToHartOp_DATA;
    end
    case(logic_command_stateReg)
      logic_command_enumDef_IDLE : begin
      end
      logic_command_enumDef_DECODE : begin
      end
      logic_command_enumDef_READ_INT_REG : begin
        logic_toHarts_payload_op = DebugDmToHartOp_EXECUTE;
      end
      logic_command_enumDef_WRITE_INT_REG : begin
        logic_toHarts_payload_op = DebugDmToHartOp_EXECUTE;
      end
      logic_command_enumDef_WAIT_DONE : begin
      end
      logic_command_enumDef_POST_EXEC : begin
        logic_toHarts_payload_op = DebugDmToHartOp_EXECUTE;
      end
      logic_command_enumDef_POST_EXEC_WAIT : begin
      end
      logic_command_enumDef_READ_FPU_REG : begin
        logic_toHarts_payload_op = DebugDmToHartOp_REG_READ;
      end
      logic_command_enumDef_WRITE_FPU_REG : begin
        logic_toHarts_payload_op = DebugDmToHartOp_REG_WRITE;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    logic_toHarts_payload_address = 5'bxxxxx;
    if(when_DebugModule_l205) begin
      logic_toHarts_payload_address = {4'd0, logic_dataX_cmdAddress};
    end
    case(logic_command_stateReg)
      logic_command_enumDef_IDLE : begin
      end
      logic_command_enumDef_DECODE : begin
      end
      logic_command_enumDef_READ_INT_REG : begin
      end
      logic_command_enumDef_WRITE_INT_REG : begin
      end
      logic_command_enumDef_WAIT_DONE : begin
      end
      logic_command_enumDef_POST_EXEC : begin
      end
      logic_command_enumDef_POST_EXEC_WAIT : begin
      end
      logic_command_enumDef_READ_FPU_REG : begin
        logic_toHarts_payload_address = logic_command_access_args_regno[4:0];
      end
      logic_command_enumDef_WRITE_FPU_REG : begin
        logic_toHarts_payload_address = logic_command_access_args_regno[4:0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    logic_toHarts_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_DebugModule_l205) begin
      logic_toHarts_payload_data = io_ctrl_cmd_payload_data;
    end
    case(logic_command_stateReg)
      logic_command_enumDef_IDLE : begin
      end
      logic_command_enumDef_DECODE : begin
      end
      logic_command_enumDef_READ_INT_REG : begin
        logic_toHarts_payload_data = (32'h7b401073 | _zz_logic_toHarts_payload_data);
      end
      logic_command_enumDef_WRITE_INT_REG : begin
        logic_toHarts_payload_data = (32'h7b402073 | _zz_logic_toHarts_payload_data_2);
      end
      logic_command_enumDef_WAIT_DONE : begin
      end
      logic_command_enumDef_POST_EXEC : begin
        logic_toHarts_payload_data = logic_progbufX_mem_spinal_port1;
      end
      logic_command_enumDef_POST_EXEC_WAIT : begin
      end
      logic_command_enumDef_READ_FPU_REG : begin
      end
      logic_command_enumDef_WRITE_FPU_REG : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    logic_toHarts_payload_size = 3'bxxx;
    logic_toHarts_payload_size = logic_command_access_args_aarsize;
  end

  assign logic_fromHarts_valid = (|{io_harts_1_hartToDm_valid,io_harts_0_hartToDm_valid});
  assign _zz_logic_fromHarts_payload_address = ((io_harts_0_hartToDm_valid ? {io_harts_0_hartToDm_payload_data,io_harts_0_hartToDm_payload_address} : 36'h0) | (io_harts_1_hartToDm_valid ? {io_harts_1_hartToDm_payload_data,io_harts_1_hartToDm_payload_address} : 36'h0));
  assign logic_fromHarts_payload_address = _zz_logic_fromHarts_payload_address[3 : 0];
  assign logic_fromHarts_payload_data = _zz_logic_fromHarts_payload_address[35 : 4];
  assign logic_harts_0_sel = (logic_dmcontrol_hartSel == 20'h0);
  assign logic_harts_0_resumeReady = ((! _zz_logic_harts_0_resumeReady) && _zz_logic_harts_0_resumeReady_1);
  assign logic_toHarts_takeWhen_valid = (logic_toHarts_valid && (! ((logic_toHarts_payload_op != DebugDmToHartOp_DATA) && (! logic_harts_0_sel))));
  assign logic_toHarts_takeWhen_payload_op = logic_toHarts_payload_op;
  assign logic_toHarts_takeWhen_payload_address = logic_toHarts_payload_address;
  assign logic_toHarts_takeWhen_payload_data = logic_toHarts_payload_data;
  assign logic_toHarts_takeWhen_payload_size = logic_toHarts_payload_size;
  assign io_harts_0_dmToHart_valid = logic_toHarts_takeWhen_valid;
  assign io_harts_0_dmToHart_payload_op = logic_toHarts_takeWhen_payload_op;
  assign io_harts_0_dmToHart_payload_address = logic_toHarts_takeWhen_payload_address;
  assign io_harts_0_dmToHart_payload_data = logic_toHarts_takeWhen_payload_data;
  assign io_harts_0_dmToHart_payload_size = logic_toHarts_takeWhen_payload_size;
  assign io_harts_0_ackReset = _zz_io_harts_0_ackReset;
  assign logic_harts_1_sel = (logic_dmcontrol_hartSel == 20'h00001);
  assign logic_harts_1_resumeReady = ((! _zz_logic_harts_1_resumeReady) && _zz_logic_harts_1_resumeReady_1);
  assign logic_toHarts_takeWhen_valid_1 = (logic_toHarts_valid && (! ((logic_toHarts_payload_op != DebugDmToHartOp_DATA) && (! logic_harts_1_sel))));
  assign logic_toHarts_takeWhen_payload_op_1 = logic_toHarts_payload_op;
  assign logic_toHarts_takeWhen_payload_address_1 = logic_toHarts_payload_address;
  assign logic_toHarts_takeWhen_payload_data_1 = logic_toHarts_payload_data;
  assign logic_toHarts_takeWhen_payload_size_1 = logic_toHarts_payload_size;
  assign io_harts_1_dmToHart_valid = logic_toHarts_takeWhen_valid_1;
  assign io_harts_1_dmToHart_payload_op = logic_toHarts_takeWhen_payload_op_1;
  assign io_harts_1_dmToHart_payload_address = logic_toHarts_takeWhen_payload_address_1;
  assign io_harts_1_dmToHart_payload_data = logic_toHarts_takeWhen_payload_data_1;
  assign io_harts_1_dmToHart_payload_size = logic_toHarts_takeWhen_payload_size_1;
  assign io_harts_1_ackReset = _zz_io_harts_1_ackReset;
  assign logic_selected_running = _zz_logic_selected_running;
  assign logic_selected_halted = _zz_logic_selected_halted;
  assign logic_selected_commit = _zz_logic_selected_commit;
  assign logic_selected_regSuccess = _zz_logic_selected_regSuccess;
  assign logic_selected_exception = _zz_logic_selected_exception;
  assign logic_selected_ebreak = _zz_logic_selected_ebreak;
  assign logic_selected_redo = _zz_logic_selected_redo;
  always @(*) begin
    logic_haltsum_value = 32'h0;
    if(when_DebugModule_l143) begin
      logic_haltsum_value[0] = io_harts_0_halted;
      logic_haltsum_value[1] = io_harts_1_halted;
    end
  end

  assign when_DebugModule_l143 = (_zz_when_DebugModule_l143 == 15'h0);
  assign logic_dmstatus_version = 4'b0010;
  assign logic_dmstatus_authenticated = 1'b1;
  assign logic_dmstatus_anyHalted = (|{(logic_harts_1_sel && io_harts_1_halted),(logic_harts_0_sel && io_harts_0_halted)});
  assign logic_dmstatus_allHalted = (&{((! logic_harts_1_sel) || io_harts_1_halted),((! logic_harts_0_sel) || io_harts_0_halted)});
  assign logic_dmstatus_anyRunning = (|{(logic_harts_1_sel && io_harts_1_running),(logic_harts_0_sel && io_harts_0_running)});
  assign logic_dmstatus_allRunning = (&{((! logic_harts_1_sel) || io_harts_1_running),((! logic_harts_0_sel) || io_harts_0_running)});
  assign logic_dmstatus_anyUnavail = (|{(logic_harts_1_sel && io_harts_1_unavailable),(logic_harts_0_sel && io_harts_0_unavailable)});
  assign logic_dmstatus_allUnavail = (&{((! logic_harts_1_sel) || io_harts_1_unavailable),((! logic_harts_0_sel) || io_harts_0_unavailable)});
  assign logic_dmstatus_anyNonExistent = (20'h00002 <= logic_dmcontrol_hartSel);
  assign logic_dmstatus_anyResumeAck = (|{(logic_harts_1_sel && logic_harts_1_resumeReady),(logic_harts_0_sel && logic_harts_0_resumeReady)});
  assign logic_dmstatus_allResumeAck = (&{((! logic_harts_1_sel) || logic_harts_1_resumeReady),((! logic_harts_0_sel) || logic_harts_0_resumeReady)});
  assign logic_dmstatus_anyHaveReset = (|{(logic_harts_1_sel && io_harts_1_haveReset),(logic_harts_0_sel && io_harts_0_haveReset)});
  assign logic_dmstatus_allHaveReset = (&{((! logic_harts_1_sel) || io_harts_1_haveReset),((! logic_harts_0_sel) || io_harts_0_haveReset)});
  assign logic_dmstatus_impebreak = 1'b1;
  assign logic_hartInfo_dataaddr = 4'b0000;
  assign logic_hartInfo_datasize = 4'b0000;
  assign logic_hartInfo_dataaccess = 1'b0;
  assign logic_hartInfo_nscratch = 4'b0000;
  assign logic_sbcs_sbversion = 3'b001;
  assign logic_sbcs_sbaccess = 3'b010;
  assign logic_progbufX_trigged = ((io_ctrl_cmd_valid && io_ctrl_cmd_payload_write) && ((io_ctrl_cmd_payload_address & 7'h70) == 7'h20));
  always @(*) begin
    logic_dataX_trigged = 1'b0;
    if(when_DebugModule_l205) begin
      logic_dataX_trigged = 1'b1;
    end
  end

  assign logic_dataX_cmdAddress = _zz_logic_dataX_cmdAddress[0:0];
  assign when_DebugModule_l205 = ((io_ctrl_cmd_valid && (7'h04 <= io_ctrl_cmd_payload_address)) && (io_ctrl_cmd_payload_address < 7'h06));
  assign _zz_factory_cmdToRsp_payload_data = logic_dataX_cmdAddress;
  assign logic_abstractcs_dataCount = 4'b0010;
  always @(*) begin
    when_BusSlaveFactory_l341 = 1'b0;
    case(io_ctrl_cmd_payload_address)
      7'h16 : begin
        if(factory_doWrite) begin
          when_BusSlaveFactory_l341 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign _zz_logic_abstractcs_cmdErr = (logic_abstractcs_cmdErr & (~ io_ctrl_cmd_payload_data[10 : 8]));
  assign logic_abstractcs_progBufSize = 5'h02;
  assign logic_abstractcs_noError = (logic_abstractcs_cmdErr == DebugModuleCmdErr_NONE);
  assign logic_abstractAuto_trigger = ((logic_progbufX_trigged && logic_abstractAuto_autoexecProgbuf[_zz_logic_abstractAuto_trigger]) || (logic_dataX_trigged && logic_abstractAuto_autoexecdata[logic_dataX_cmdAddress]));
  assign logic_command_wantExit = 1'b0;
  always @(*) begin
    logic_command_wantStart = 1'b0;
    case(logic_command_stateReg)
      logic_command_enumDef_IDLE : begin
      end
      logic_command_enumDef_DECODE : begin
      end
      logic_command_enumDef_READ_INT_REG : begin
      end
      logic_command_enumDef_WRITE_INT_REG : begin
      end
      logic_command_enumDef_WAIT_DONE : begin
      end
      logic_command_enumDef_POST_EXEC : begin
      end
      logic_command_enumDef_POST_EXEC_WAIT : begin
      end
      logic_command_enumDef_READ_FPU_REG : begin
      end
      logic_command_enumDef_WRITE_FPU_REG : begin
      end
      default : begin
        logic_command_wantStart = 1'b1;
      end
    endcase
  end

  assign logic_command_wantKill = 1'b0;
  always @(*) begin
    logic_command_commandRequest = 1'b0;
    case(io_ctrl_cmd_payload_address)
      7'h17 : begin
        if(factory_doWrite) begin
          logic_command_commandRequest = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign _zz_logic_command_access_args_regno = logic_command_data;
  assign logic_command_access_args_regno = _zz_logic_command_access_args_regno[15 : 0];
  assign logic_command_access_args_write = _zz_logic_command_access_args_regno[16];
  assign logic_command_access_args_transfer = _zz_logic_command_access_args_regno[17];
  assign logic_command_access_args_postExec = _zz_logic_command_access_args_regno[18];
  assign logic_command_access_args_aarpostincrement = _zz_logic_command_access_args_regno[19];
  assign logic_command_access_args_aarsize = _zz_logic_command_access_args_regno[22 : 20];
  assign logic_command_access_transferFloat = logic_command_access_args_regno[5];
  assign logic_command_access_notSupported = (((_zz_logic_command_access_notSupported < logic_command_access_args_aarsize) || logic_command_access_args_aarpostincrement) || (logic_command_access_args_transfer && (logic_command_access_args_regno[15 : 6] != 10'h040)));
  assign logic_command_request = (logic_command_commandRequest || logic_abstractAuto_trigger);
  assign when_DebugModule_l260 = ((logic_command_request && logic_abstractcs_busy) && logic_abstractcs_noError);
  assign when_DebugModule_l263 = (|{io_harts_1_exception,io_harts_0_exception});
  assign when_DebugModule_l266 = ((logic_abstractcs_busy && (logic_progbufX_trigged || logic_dataX_trigged)) && logic_abstractcs_noError);
  assign logic_dmcontrol_hartSelLoNew = io_ctrl_cmd_payload_data[25 : 16];
  assign logic_dmcontrol_hartSelHiNew = io_ctrl_cmd_payload_data[15 : 6];
  always @(*) begin
    logic_command_stateNext = logic_command_stateReg;
    case(logic_command_stateReg)
      logic_command_enumDef_IDLE : begin
        if(when_DebugModule_l275) begin
          if(!when_DebugModule_l276) begin
            logic_command_stateNext = logic_command_enumDef_DECODE;
          end
        end
      end
      logic_command_enumDef_DECODE : begin
        logic_command_stateNext = logic_command_enumDef_IDLE;
        case(switch_DebugModule_l287)
          8'h0 : begin
            if(!logic_command_access_notSupported) begin
              if(logic_command_access_args_postExec) begin
                logic_command_stateNext = logic_command_enumDef_POST_EXEC;
              end
              if(logic_command_access_args_transfer) begin
                if(when_DebugModule_l296) begin
                  if(logic_command_access_args_write) begin
                    logic_command_stateNext = logic_command_enumDef_WRITE_INT_REG;
                  end else begin
                    logic_command_stateNext = logic_command_enumDef_READ_INT_REG;
                  end
                end else begin
                  if(logic_command_access_args_write) begin
                    logic_command_stateNext = logic_command_enumDef_WRITE_FPU_REG;
                  end else begin
                    logic_command_stateNext = logic_command_enumDef_READ_FPU_REG;
                  end
                end
              end
            end
          end
          default : begin
          end
        endcase
      end
      logic_command_enumDef_READ_INT_REG : begin
        logic_command_stateNext = logic_command_enumDef_WAIT_DONE;
      end
      logic_command_enumDef_WRITE_INT_REG : begin
        logic_command_stateNext = logic_command_enumDef_WAIT_DONE;
      end
      logic_command_enumDef_WAIT_DONE : begin
        if(when_DebugModule_l350) begin
          logic_command_stateNext = logic_command_enumDef_IDLE;
          if(logic_command_access_args_postExec) begin
            logic_command_stateNext = logic_command_enumDef_POST_EXEC;
          end
        end
      end
      logic_command_enumDef_POST_EXEC : begin
        logic_command_stateNext = logic_command_enumDef_POST_EXEC_WAIT;
      end
      logic_command_enumDef_POST_EXEC_WAIT : begin
        if(when_DebugModule_l366) begin
          logic_command_stateNext = logic_command_enumDef_IDLE;
        end
        if(when_DebugModule_l370) begin
          logic_command_stateNext = logic_command_enumDef_POST_EXEC;
        end
      end
      logic_command_enumDef_READ_FPU_REG : begin
        logic_command_stateNext = logic_command_enumDef_WAIT_DONE;
      end
      logic_command_enumDef_WRITE_FPU_REG : begin
        logic_command_stateNext = logic_command_enumDef_WAIT_DONE;
      end
      default : begin
      end
    endcase
    if(logic_command_wantStart) begin
      logic_command_stateNext = logic_command_enumDef_IDLE;
    end
    if(logic_command_wantKill) begin
      logic_command_stateNext = logic_command_enumDef_BOOT;
    end
  end

  assign when_DebugModule_l275 = (logic_command_request && logic_abstractcs_noError);
  assign when_DebugModule_l276 = (! _zz_when_DebugModule_l276);
  assign switch_DebugModule_l287 = logic_command_data[31 : 24];
  assign when_DebugModule_l296 = (! logic_command_access_args_regno[5]);
  assign when_DebugModule_l350 = (logic_selected_commit || logic_selected_regSuccess);
  assign when_DebugModule_l366 = ((logic_selected_ebreak || logic_selected_exception) || logic_selected_commit);
  assign when_DebugModule_l370 = (logic_selected_redo || (logic_selected_commit && (logic_command_executionCounter != 1'b1)));
  assign when_StateMachine_l253 = ((! (logic_command_stateReg == logic_command_enumDef_IDLE)) && (logic_command_stateNext == logic_command_enumDef_IDLE));
  always @(posedge io_systemClk) begin
    if(debugCd_logic_outputReset) begin
      factory_rspBuffer_valid <= 1'b0;
      dmactive <= 1'b0;
    end else begin
      factory_rspBuffer_valid <= factory_cmdToRsp_valid;
      case(io_ctrl_cmd_payload_address)
        7'h10 : begin
          if(factory_doWrite) begin
            dmactive <= io_ctrl_cmd_payload_data[0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge io_systemClk) begin
    factory_rspBuffer_payload_error <= factory_cmdToRsp_payload_error;
    factory_rspBuffer_payload_data <= factory_cmdToRsp_payload_data;
  end

  always @(posedge io_systemClk or negedge dmactive) begin
    if(!dmactive) begin
      logic_dmcontrol_ndmreset <= 1'b0;
      logic_dmcontrol_hartSelLo <= 10'h0;
      logic_dmcontrol_hartSelHi <= 10'h0;
      logic_dmcontrol_harts_0_haltReq <= 1'b0;
      logic_dmcontrol_harts_1_haltReq <= 1'b0;
      _zz_logic_harts_0_resumeReady <= 1'b0;
      _zz_logic_harts_0_resumeReady_1 <= 1'b0;
      _zz_logic_harts_1_resumeReady <= 1'b0;
      _zz_logic_harts_1_resumeReady_1 <= 1'b0;
      logic_abstractcs_cmdErr <= DebugModuleCmdErr_NONE;
      logic_abstractcs_busy <= 1'b0;
      logic_abstractAuto_autoexecdata <= 2'b00;
      logic_abstractAuto_autoexecProgbuf <= 2'b00;
      logic_command_stateReg <= logic_command_enumDef_BOOT;
    end else begin
      if(when_DebugModule_l102) begin
        logic_dmcontrol_harts_0_haltReq <= ((logic_dmcontrol_harts_0_haltReq || logic_dmcontrol_haltSet) && (! logic_dmcontrol_haltClear));
      end
      if(when_DebugModule_l102_1) begin
        logic_dmcontrol_harts_1_haltReq <= ((logic_dmcontrol_harts_1_haltReq || logic_dmcontrol_haltSet) && (! logic_dmcontrol_haltClear));
      end
      if(io_harts_0_resume_cmd_valid) begin
        _zz_logic_harts_0_resumeReady <= 1'b1;
      end
      if(io_harts_0_resume_rsp_valid) begin
        _zz_logic_harts_0_resumeReady <= 1'b0;
      end
      if(io_harts_0_resume_cmd_valid) begin
        _zz_logic_harts_0_resumeReady_1 <= 1'b1;
      end
      if(io_harts_1_resume_cmd_valid) begin
        _zz_logic_harts_1_resumeReady <= 1'b1;
      end
      if(io_harts_1_resume_rsp_valid) begin
        _zz_logic_harts_1_resumeReady <= 1'b0;
      end
      if(io_harts_1_resume_cmd_valid) begin
        _zz_logic_harts_1_resumeReady_1 <= 1'b1;
      end
      if(when_BusSlaveFactory_l341) begin
        logic_abstractcs_cmdErr <= _zz_logic_abstractcs_cmdErr;
      end
      if(when_DebugModule_l260) begin
        logic_abstractcs_cmdErr <= DebugModuleCmdErr_BUSY;
      end
      if(when_DebugModule_l263) begin
        logic_abstractcs_cmdErr <= DebugModuleCmdErr_EXCEPTION;
      end
      if(when_DebugModule_l266) begin
        logic_abstractcs_cmdErr <= DebugModuleCmdErr_BUSY;
      end
      case(io_ctrl_cmd_payload_address)
        7'h10 : begin
          if(factory_doWrite) begin
            logic_dmcontrol_ndmreset <= io_ctrl_cmd_payload_data[1];
            logic_dmcontrol_hartSelLo <= io_ctrl_cmd_payload_data[25 : 16];
            logic_dmcontrol_hartSelHi <= io_ctrl_cmd_payload_data[15 : 6];
          end
        end
        7'h18 : begin
          if(factory_doWrite) begin
            logic_abstractAuto_autoexecdata <= io_ctrl_cmd_payload_data[1 : 0];
            logic_abstractAuto_autoexecProgbuf <= io_ctrl_cmd_payload_data[17 : 16];
          end
        end
        default : begin
        end
      endcase
      logic_command_stateReg <= logic_command_stateNext;
      case(logic_command_stateReg)
        logic_command_enumDef_IDLE : begin
          if(when_DebugModule_l275) begin
            if(when_DebugModule_l276) begin
              logic_abstractcs_cmdErr <= DebugModuleCmdErr_HALT_RESUME;
            end else begin
              logic_abstractcs_busy <= 1'b1;
            end
          end
        end
        logic_command_enumDef_DECODE : begin
          case(switch_DebugModule_l287)
            8'h0 : begin
              if(logic_command_access_notSupported) begin
                logic_abstractcs_cmdErr <= DebugModuleCmdErr_NOT_SUPPORTED;
              end
            end
            default : begin
              logic_abstractcs_cmdErr <= DebugModuleCmdErr_NOT_SUPPORTED;
            end
          endcase
        end
        logic_command_enumDef_READ_INT_REG : begin
        end
        logic_command_enumDef_WRITE_INT_REG : begin
        end
        logic_command_enumDef_WAIT_DONE : begin
        end
        logic_command_enumDef_POST_EXEC : begin
        end
        logic_command_enumDef_POST_EXEC_WAIT : begin
        end
        logic_command_enumDef_READ_FPU_REG : begin
        end
        logic_command_enumDef_WRITE_FPU_REG : begin
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l253) begin
        logic_abstractcs_busy <= 1'b0;
      end
    end
  end

  always @(posedge io_systemClk) begin
    _zz_io_harts_0_ackReset <= (logic_harts_0_sel && logic_dmcontrol_ackhavereset);
    _zz_io_harts_1_ackReset <= (logic_harts_1_sel && logic_dmcontrol_ackhavereset);
    case(io_ctrl_cmd_payload_address)
      7'h17 : begin
        if(factory_doWrite) begin
          logic_command_data <= io_ctrl_cmd_payload_data[31 : 0];
        end
      end
      default : begin
      end
    endcase
    case(logic_command_stateReg)
      logic_command_enumDef_IDLE : begin
        logic_command_executionCounter <= 1'b0;
        if(when_DebugModule_l275) begin
          if(!when_DebugModule_l276) begin
            logic_selected_hart <= logic_dmcontrol_hartSel[0:0];
          end
        end
      end
      logic_command_enumDef_DECODE : begin
      end
      logic_command_enumDef_READ_INT_REG : begin
      end
      logic_command_enumDef_WRITE_INT_REG : begin
      end
      logic_command_enumDef_WAIT_DONE : begin
      end
      logic_command_enumDef_POST_EXEC : begin
      end
      logic_command_enumDef_POST_EXEC_WAIT : begin
        if(when_DebugModule_l366) begin
          logic_command_executionCounter <= (logic_command_executionCounter + 1'b1);
        end
      end
      logic_command_enumDef_READ_FPU_REG : begin
      end
      logic_command_enumDef_WRITE_FPU_REG : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module FpuCore (
  input  wire          io_port_0_cmd_valid,
  output wire          io_port_0_cmd_ready,
  input  wire [3:0]    io_port_0_cmd_payload_opcode,
  input  wire [1:0]    io_port_0_cmd_payload_arg,
  input  wire [4:0]    io_port_0_cmd_payload_rs1,
  input  wire [4:0]    io_port_0_cmd_payload_rs2,
  input  wire [4:0]    io_port_0_cmd_payload_rs3,
  input  wire [4:0]    io_port_0_cmd_payload_rd,
  input  wire [0:0]    io_port_0_cmd_payload_format,
  input  wire [2:0]    io_port_0_cmd_payload_roundMode,
  input  wire          io_port_0_commit_valid,
  output wire          io_port_0_commit_ready,
  input  wire [3:0]    io_port_0_commit_payload_opcode,
  input  wire [4:0]    io_port_0_commit_payload_rd,
  input  wire          io_port_0_commit_payload_write,
  input  wire [63:0]   io_port_0_commit_payload_value,
  output wire          io_port_0_rsp_valid,
  input  wire          io_port_0_rsp_ready,
  output wire [63:0]   io_port_0_rsp_payload_value,
  output wire          io_port_0_rsp_payload_NV,
  output wire          io_port_0_rsp_payload_NX,
  output wire          io_port_0_completion_valid,
  output wire          io_port_0_completion_payload_flags_NX,
  output wire          io_port_0_completion_payload_flags_UF,
  output wire          io_port_0_completion_payload_flags_OF,
  output wire          io_port_0_completion_payload_flags_DZ,
  output wire          io_port_0_completion_payload_flags_NV,
  output wire          io_port_0_completion_payload_written,
  input  wire          io_port_1_cmd_valid,
  output wire          io_port_1_cmd_ready,
  input  wire [3:0]    io_port_1_cmd_payload_opcode,
  input  wire [1:0]    io_port_1_cmd_payload_arg,
  input  wire [4:0]    io_port_1_cmd_payload_rs1,
  input  wire [4:0]    io_port_1_cmd_payload_rs2,
  input  wire [4:0]    io_port_1_cmd_payload_rs3,
  input  wire [4:0]    io_port_1_cmd_payload_rd,
  input  wire [0:0]    io_port_1_cmd_payload_format,
  input  wire [2:0]    io_port_1_cmd_payload_roundMode,
  input  wire          io_port_1_commit_valid,
  output wire          io_port_1_commit_ready,
  input  wire [3:0]    io_port_1_commit_payload_opcode,
  input  wire [4:0]    io_port_1_commit_payload_rd,
  input  wire          io_port_1_commit_payload_write,
  input  wire [63:0]   io_port_1_commit_payload_value,
  output wire          io_port_1_rsp_valid,
  input  wire          io_port_1_rsp_ready,
  output wire [63:0]   io_port_1_rsp_payload_value,
  output wire          io_port_1_rsp_payload_NV,
  output wire          io_port_1_rsp_payload_NX,
  output wire          io_port_1_completion_valid,
  output wire          io_port_1_completion_payload_flags_NX,
  output wire          io_port_1_completion_payload_flags_UF,
  output wire          io_port_1_completion_payload_flags_OF,
  output wire          io_port_1_completion_payload_flags_DZ,
  output wire          io_port_1_completion_payload_flags_NV,
  output wire          io_port_1_completion_payload_written,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);
  localparam FpuOpcode_LOAD = 4'd0;
  localparam FpuOpcode_STORE = 4'd1;
  localparam FpuOpcode_MUL = 4'd2;
  localparam FpuOpcode_ADD = 4'd3;
  localparam FpuOpcode_FMA = 4'd4;
  localparam FpuOpcode_I2F = 4'd5;
  localparam FpuOpcode_F2I = 4'd6;
  localparam FpuOpcode_CMP = 4'd7;
  localparam FpuOpcode_DIV = 4'd8;
  localparam FpuOpcode_SQRT = 4'd9;
  localparam FpuOpcode_MIN_MAX = 4'd10;
  localparam FpuOpcode_SGNJ = 4'd11;
  localparam FpuOpcode_FMV_X_W = 4'd12;
  localparam FpuOpcode_FMV_W_X = 4'd13;
  localparam FpuOpcode_FCLASS = 4'd14;
  localparam FpuOpcode_FCVT_X_X = 4'd15;
  localparam FpuFormat_FLOAT = 1'd0;
  localparam FpuFormat_DOUBLE = 1'd1;
  localparam FpuRoundMode_RNE = 3'd0;
  localparam FpuRoundMode_RTZ = 3'd1;
  localparam FpuRoundMode_RDN = 3'd2;
  localparam FpuRoundMode_RUP = 3'd3;
  localparam FpuRoundMode_RMM = 3'd4;

  wire                div_divider_io_input_valid;
  wire                sqrt_sqrt_io_input_valid;
  wire       [53:0]   sqrt_sqrt_io_input_payload_a;
  reg        [66:0]   rf_ram_spinal_port0;
  reg        [66:0]   rf_ram_spinal_port1;
  reg        [66:0]   rf_ram_spinal_port2;
  wire       [0:0]    rf_scoreboards_0_target_spinal_port1;
  wire       [0:0]    rf_scoreboards_0_target_spinal_port2;
  wire       [0:0]    rf_scoreboards_0_target_spinal_port3;
  wire       [0:0]    rf_scoreboards_0_target_spinal_port4;
  wire       [0:0]    rf_scoreboards_0_hit_spinal_port1;
  wire       [0:0]    rf_scoreboards_0_hit_spinal_port2;
  wire       [0:0]    rf_scoreboards_0_hit_spinal_port3;
  wire       [0:0]    rf_scoreboards_0_hit_spinal_port4;
  wire       [0:0]    rf_scoreboards_0_hit_spinal_port5;
  wire       [0:0]    rf_scoreboards_0_writes_spinal_port1;
  wire       [0:0]    rf_scoreboards_1_target_spinal_port1;
  wire       [0:0]    rf_scoreboards_1_target_spinal_port2;
  wire       [0:0]    rf_scoreboards_1_target_spinal_port3;
  wire       [0:0]    rf_scoreboards_1_target_spinal_port4;
  wire       [0:0]    rf_scoreboards_1_hit_spinal_port1;
  wire       [0:0]    rf_scoreboards_1_hit_spinal_port2;
  wire       [0:0]    rf_scoreboards_1_hit_spinal_port3;
  wire       [0:0]    rf_scoreboards_1_hit_spinal_port4;
  wire       [0:0]    rf_scoreboards_1_hit_spinal_port5;
  wire       [0:0]    rf_scoreboards_1_writes_spinal_port1;
  wire                streamFork_3_io_input_ready;
  wire                streamFork_3_io_outputs_0_valid;
  wire       [3:0]    streamFork_3_io_outputs_0_payload_opcode;
  wire       [4:0]    streamFork_3_io_outputs_0_payload_rd;
  wire                streamFork_3_io_outputs_0_payload_write;
  wire       [63:0]   streamFork_3_io_outputs_0_payload_value;
  wire                streamFork_3_io_outputs_1_valid;
  wire       [3:0]    streamFork_3_io_outputs_1_payload_opcode;
  wire       [4:0]    streamFork_3_io_outputs_1_payload_rd;
  wire                streamFork_3_io_outputs_1_payload_write;
  wire       [63:0]   streamFork_3_io_outputs_1_payload_value;
  wire                streamFork_4_io_input_ready;
  wire                streamFork_4_io_outputs_0_valid;
  wire       [3:0]    streamFork_4_io_outputs_0_payload_opcode;
  wire       [4:0]    streamFork_4_io_outputs_0_payload_rd;
  wire                streamFork_4_io_outputs_0_payload_write;
  wire       [63:0]   streamFork_4_io_outputs_0_payload_value;
  wire                streamFork_4_io_outputs_1_valid;
  wire       [3:0]    streamFork_4_io_outputs_1_payload_opcode;
  wire       [4:0]    streamFork_4_io_outputs_1_payload_rd;
  wire                streamFork_4_io_outputs_1_payload_write;
  wire       [63:0]   streamFork_4_io_outputs_1_payload_value;
  wire                cmdArbiter_arbiter_io_inputs_0_ready;
  wire                cmdArbiter_arbiter_io_inputs_1_ready;
  wire                cmdArbiter_arbiter_io_output_valid;
  wire       [3:0]    cmdArbiter_arbiter_io_output_payload_opcode;
  wire       [1:0]    cmdArbiter_arbiter_io_output_payload_arg;
  wire       [4:0]    cmdArbiter_arbiter_io_output_payload_rs1;
  wire       [4:0]    cmdArbiter_arbiter_io_output_payload_rs2;
  wire       [4:0]    cmdArbiter_arbiter_io_output_payload_rs3;
  wire       [4:0]    cmdArbiter_arbiter_io_output_payload_rd;
  wire       [0:0]    cmdArbiter_arbiter_io_output_payload_format;
  wire       [2:0]    cmdArbiter_arbiter_io_output_payload_roundMode;
  wire       [0:0]    cmdArbiter_arbiter_io_chosen;
  wire       [1:0]    cmdArbiter_arbiter_io_chosenOH;
  wire                div_divider_io_input_ready;
  wire                div_divider_io_output_valid;
  wire       [54:0]   div_divider_io_output_payload_result;
  wire       [52:0]   div_divider_io_output_payload_remain;
  wire                sqrt_sqrt_io_input_ready;
  wire                sqrt_sqrt_io_output_valid;
  wire       [52:0]   sqrt_sqrt_io_output_payload_result;
  wire       [56:0]   sqrt_sqrt_io_output_payload_remain;
  wire                streamArbiter_10_io_inputs_0_ready;
  wire                streamArbiter_10_io_inputs_1_ready;
  wire                streamArbiter_10_io_inputs_2_ready;
  wire                streamArbiter_10_io_inputs_3_ready;
  wire                streamArbiter_10_io_inputs_4_ready;
  wire                streamArbiter_10_io_inputs_5_ready;
  wire                streamArbiter_10_io_output_valid;
  wire       [0:0]    streamArbiter_10_io_output_payload_source;
  wire       [4:0]    streamArbiter_10_io_output_payload_rd;
  wire       [52:0]   streamArbiter_10_io_output_payload_value_mantissa;
  wire       [11:0]   streamArbiter_10_io_output_payload_value_exponent;
  wire                streamArbiter_10_io_output_payload_value_sign;
  wire                streamArbiter_10_io_output_payload_value_special;
  wire                streamArbiter_10_io_output_payload_scrap;
  wire       [2:0]    streamArbiter_10_io_output_payload_roundMode;
  wire       [0:0]    streamArbiter_10_io_output_payload_format;
  wire                streamArbiter_10_io_output_payload_NV;
  wire                streamArbiter_10_io_output_payload_DZ;
  wire       [2:0]    streamArbiter_10_io_chosen;
  wire       [5:0]    streamArbiter_10_io_chosenOH;
  wire       [0:0]    _zz_rf_scoreboards_0_target_port;
  wire       [0:0]    _zz_rf_scoreboards_0_hit_port;
  wire       [0:0]    _zz_rf_scoreboards_1_target_port;
  wire       [0:0]    _zz_rf_scoreboards_1_hit_port;
  wire       [3:0]    _zz_commitLogic_0_pending_counter;
  wire       [3:0]    _zz_commitLogic_0_pending_counter_1;
  wire       [0:0]    _zz_commitLogic_0_pending_counter_2;
  wire       [3:0]    _zz_commitLogic_0_pending_counter_3;
  wire       [0:0]    _zz_commitLogic_0_pending_counter_4;
  wire       [3:0]    _zz_commitLogic_0_add_counter;
  wire       [3:0]    _zz_commitLogic_0_add_counter_1;
  wire       [0:0]    _zz_commitLogic_0_add_counter_2;
  wire       [3:0]    _zz_commitLogic_0_add_counter_3;
  wire       [0:0]    _zz_commitLogic_0_add_counter_4;
  wire       [3:0]    _zz_commitLogic_0_mul_counter;
  wire       [3:0]    _zz_commitLogic_0_mul_counter_1;
  wire       [0:0]    _zz_commitLogic_0_mul_counter_2;
  wire       [3:0]    _zz_commitLogic_0_mul_counter_3;
  wire       [0:0]    _zz_commitLogic_0_mul_counter_4;
  wire       [3:0]    _zz_commitLogic_0_div_counter;
  wire       [3:0]    _zz_commitLogic_0_div_counter_1;
  wire       [0:0]    _zz_commitLogic_0_div_counter_2;
  wire       [3:0]    _zz_commitLogic_0_div_counter_3;
  wire       [0:0]    _zz_commitLogic_0_div_counter_4;
  wire       [3:0]    _zz_commitLogic_0_sqrt_counter;
  wire       [3:0]    _zz_commitLogic_0_sqrt_counter_1;
  wire       [0:0]    _zz_commitLogic_0_sqrt_counter_2;
  wire       [3:0]    _zz_commitLogic_0_sqrt_counter_3;
  wire       [0:0]    _zz_commitLogic_0_sqrt_counter_4;
  wire       [3:0]    _zz_commitLogic_0_short_counter;
  wire       [3:0]    _zz_commitLogic_0_short_counter_1;
  wire       [0:0]    _zz_commitLogic_0_short_counter_2;
  wire       [3:0]    _zz_commitLogic_0_short_counter_3;
  wire       [0:0]    _zz_commitLogic_0_short_counter_4;
  wire       [0:0]    _zz_rf_scoreboards_0_writes_port;
  wire       [3:0]    _zz_commitLogic_1_pending_counter;
  wire       [3:0]    _zz_commitLogic_1_pending_counter_1;
  wire       [0:0]    _zz_commitLogic_1_pending_counter_2;
  wire       [3:0]    _zz_commitLogic_1_pending_counter_3;
  wire       [0:0]    _zz_commitLogic_1_pending_counter_4;
  wire       [3:0]    _zz_commitLogic_1_add_counter;
  wire       [3:0]    _zz_commitLogic_1_add_counter_1;
  wire       [0:0]    _zz_commitLogic_1_add_counter_2;
  wire       [3:0]    _zz_commitLogic_1_add_counter_3;
  wire       [0:0]    _zz_commitLogic_1_add_counter_4;
  wire       [3:0]    _zz_commitLogic_1_mul_counter;
  wire       [3:0]    _zz_commitLogic_1_mul_counter_1;
  wire       [0:0]    _zz_commitLogic_1_mul_counter_2;
  wire       [3:0]    _zz_commitLogic_1_mul_counter_3;
  wire       [0:0]    _zz_commitLogic_1_mul_counter_4;
  wire       [3:0]    _zz_commitLogic_1_div_counter;
  wire       [3:0]    _zz_commitLogic_1_div_counter_1;
  wire       [0:0]    _zz_commitLogic_1_div_counter_2;
  wire       [3:0]    _zz_commitLogic_1_div_counter_3;
  wire       [0:0]    _zz_commitLogic_1_div_counter_4;
  wire       [3:0]    _zz_commitLogic_1_sqrt_counter;
  wire       [3:0]    _zz_commitLogic_1_sqrt_counter_1;
  wire       [0:0]    _zz_commitLogic_1_sqrt_counter_2;
  wire       [3:0]    _zz_commitLogic_1_sqrt_counter_3;
  wire       [0:0]    _zz_commitLogic_1_sqrt_counter_4;
  wire       [3:0]    _zz_commitLogic_1_short_counter;
  wire       [3:0]    _zz_commitLogic_1_short_counter_1;
  wire       [0:0]    _zz_commitLogic_1_short_counter_2;
  wire       [3:0]    _zz_commitLogic_1_short_counter_3;
  wire       [0:0]    _zz_commitLogic_1_short_counter_4;
  wire       [0:0]    _zz_rf_scoreboards_1_writes_port;
  wire       [3:0]    _zz_decode_shortPipHit;
  wire                _zz_decode_shortPipHit_1;
  wire       [0:0]    _zz_decode_shortPipHit_2;
  wire       [0:0]    _zz_decode_shortPipHit_3;
  reg                 _zz_load_s0_hazard;
  reg        [63:0]   _zz_load_s0_output_payload_value;
  wire       [51:0]   _zz_load_s1_fsm_shift_input_1;
  wire       [51:0]   _zz_load_s1_fsm_shift_input_2;
  wire       [51:0]   _zz_load_s1_fsm_shift_input_3;
  wire       [51:0]   _zz_load_s1_fsm_shift_input_4;
  wire       [51:0]   _zz_load_s1_fsm_shift_input_5;
  wire       [51:0]   _zz_load_s1_fsm_shift_input_6;
  wire       [31:0]   _zz_load_s0_output_rData_value_2;
  wire       [64:0]   _zz_load_s0_output_rData_value_3;
  wire       [64:0]   _zz_load_s0_output_rData_value_4;
  wire       [64:0]   _zz_load_s0_output_rData_value_5;
  wire       [0:0]    _zz_load_s0_output_rData_value_6;
  wire                _zz__zz_load_s1_fsm_shift_by;
  wire       [0:0]    _zz__zz_load_s1_fsm_shift_by_1;
  wire       [42:0]   _zz__zz_load_s1_fsm_shift_by_2;
  wire                _zz__zz_load_s1_fsm_shift_by_3;
  wire       [0:0]    _zz__zz_load_s1_fsm_shift_by_4;
  wire       [31:0]   _zz__zz_load_s1_fsm_shift_by_5;
  wire                _zz__zz_load_s1_fsm_shift_by_6;
  wire       [0:0]    _zz__zz_load_s1_fsm_shift_by_7;
  wire       [20:0]   _zz__zz_load_s1_fsm_shift_by_8;
  wire                _zz__zz_load_s1_fsm_shift_by_9;
  wire       [0:0]    _zz__zz_load_s1_fsm_shift_by_10;
  wire       [9:0]    _zz__zz_load_s1_fsm_shift_by_11;
  wire       [51:0]   _zz__zz_load_s1_fsm_shift_by_1_1;
  wire                _zz__zz_load_s1_fsm_shift_by_47;
  wire                _zz__zz_load_s1_fsm_shift_by_48;
  wire                _zz__zz_load_s1_fsm_shift_by_49;
  wire                _zz__zz_load_s1_fsm_shift_by_50;
  wire                _zz__zz_load_s1_fsm_shift_by_51;
  wire                _zz__zz_load_s1_fsm_shift_by_52;
  wire       [12:0]   _zz_load_s1_recoded_exponent;
  wire       [12:0]   _zz_load_s1_recoded_exponent_1;
  wire       [12:0]   _zz_load_s1_recoded_exponent_2;
  wire       [11:0]   _zz_load_s1_output_payload_value_exponent;
  reg                 _zz_shortPip_isCommited;
  wire       [11:0]   _zz_shortPip_f32_exp;
  wire       [11:0]   _zz_shortPip_f64_exp;
  wire       [11:0]   _zz_shortPip_expInSubnormalRange;
  wire       [52:0]   _zz_shortPip_fsm_shift_input_1;
  wire       [52:0]   _zz_shortPip_fsm_shift_input_2;
  wire       [52:0]   _zz_shortPip_fsm_shift_input_3;
  wire       [52:0]   _zz_shortPip_fsm_shift_input_4;
  wire       [52:0]   _zz_shortPip_fsm_shift_input_5;
  wire       [52:0]   _zz_shortPip_fsm_shift_input_6;
  wire       [11:0]   _zz_shortPip_fsm_shift_by_2;
  wire       [11:0]   _zz_shortPip_fsm_shift_by_3;
  wire       [11:0]   _zz_shortPip_fsm_shift_by_4;
  wire       [11:0]   _zz_shortPip_fsm_shift_by_5;
  wire       [11:0]   _zz_shortPip_fsm_shift_by_6;
  wire       [31:0]   _zz_shortPip_f2i_result;
  wire       [0:0]    _zz_shortPip_f2i_result_1;
  wire       [30:0]   _zz_shortPip_f2i_underflow;
  wire       [30:0]   _zz_shortPip_f2i_underflow_1;
  reg                 _zz_shortPip_input_ready;
  wire       [105:0]  _zz_mul_sum1_sum;
  wire       [105:0]  _zz_mul_sum1_sum_1;
  wire       [105:0]  _zz_mul_sum1_sum_2;
  wire       [53:0]   _zz_mul_sum1_sum_3;
  wire       [105:0]  _zz_mul_sum1_sum_4;
  wire       [105:0]  _zz_mul_sum1_sum_5;
  wire       [53:0]   _zz_mul_sum1_sum_6;
  wire       [105:0]  _zz_mul_sum1_sum_7;
  wire       [70:0]   _zz_mul_sum1_sum_8;
  wire       [105:0]  _zz_mul_sum2_sum;
  wire       [105:0]  _zz_mul_sum2_sum_1;
  wire       [105:0]  _zz_mul_sum2_sum_2;
  wire       [105:0]  _zz_mul_sum2_sum_3;
  wire       [70:0]   _zz_mul_sum2_sum_4;
  wire       [105:0]  _zz_mul_sum2_sum_5;
  wire       [71:0]   _zz_mul_sum2_sum_6;
  wire       [105:0]  _zz_mul_sum2_sum_7;
  wire       [105:0]  _zz_mul_sum2_sum_8;
  wire       [88:0]   _zz_mul_sum2_sum_9;
  wire       [105:0]  _zz_mul_sum2_sum_10;
  wire       [88:0]   _zz_mul_sum2_sum_11;
  wire       [105:0]  _zz_mul_sum2_sum_12;
  reg                 _zz_mul_sum2_isCommited;
  wire       [12:0]   _zz_mul_norm_exp;
  wire       [0:0]    _zz_mul_norm_exp_1;
  wire       [12:0]   _zz_mul_norm_forceUnderflow;
  wire       [12:0]   _zz_mul_norm_output_exponent;
  reg                 _zz_div_isCommited;
  wire       [13:0]   _zz_div_exponent;
  wire       [13:0]   _zz_div_exponent_1;
  wire       [13:0]   _zz_div_exponent_2;
  wire       [13:0]   _zz_div_exponent_3;
  wire       [13:0]   _zz_div_exponent_4;
  wire       [0:0]    _zz_div_exponent_5;
  reg                 _zz_sqrt_isCommited;
  wire       [11:0]   _zz_sqrt_exponent;
  wire       [11:0]   _zz_sqrt_exponent_1;
  wire       [10:0]   _zz_sqrt_exponent_2;
  wire       [10:0]   _zz_sqrt_exponent_3;
  wire       [11:0]   _zz_sqrt_exponent_4;
  wire       [0:0]    _zz_sqrt_exponent_5;
  wire       [12:0]   _zz_add_shifter_shiftBy_1;
  wire       [12:0]   _zz_add_shifter_shiftBy_2;
  wire       [12:0]   _zz_add_shifter_shiftBy_3;
  wire       [0:0]    _zz_add_shifter_shiftBy_4;
  wire       [54:0]   _zz_add_shifter_yMantissa_1;
  wire       [54:0]   _zz_add_shifter_yMantissa_2;
  wire       [54:0]   _zz_add_shifter_yMantissa_3;
  wire       [54:0]   _zz_add_shifter_yMantissa_4;
  wire       [54:0]   _zz_add_shifter_yMantissa_5;
  wire       [54:0]   _zz_add_shifter_yMantissa_6;
  wire       [55:0]   _zz_add_math_xSigned;
  wire       [55:0]   _zz_add_math_xSigned_1;
  wire       [0:0]    _zz_add_math_xSigned_2;
  wire       [55:0]   _zz_add_math_ySigned;
  wire       [55:0]   _zz_add_math_ySigned_1;
  wire       [0:0]    _zz_add_math_ySigned_2;
  wire       [56:0]   _zz_add_math_output_payload_xyMantissa;
  wire       [56:0]   _zz_add_math_output_payload_xyMantissa_1;
  wire       [56:0]   _zz_add_math_output_payload_xyMantissa_2;
  wire       [56:0]   _zz_add_math_output_payload_xyMantissa_3;
  reg                 _zz_add_oh_isCommited;
  wire                _zz__zz_add_oh_shift;
  wire       [0:0]    _zz__zz_add_oh_shift_1;
  wire       [46:0]   _zz__zz_add_oh_shift_2;
  wire                _zz__zz_add_oh_shift_3;
  wire       [0:0]    _zz__zz_add_oh_shift_4;
  wire       [35:0]   _zz__zz_add_oh_shift_5;
  wire                _zz__zz_add_oh_shift_6;
  wire       [0:0]    _zz__zz_add_oh_shift_7;
  wire       [24:0]   _zz__zz_add_oh_shift_8;
  wire                _zz__zz_add_oh_shift_9;
  wire       [0:0]    _zz__zz_add_oh_shift_10;
  wire       [13:0]   _zz__zz_add_oh_shift_11;
  wire                _zz__zz_add_oh_shift_12;
  wire       [0:0]    _zz__zz_add_oh_shift_13;
  wire       [2:0]    _zz__zz_add_oh_shift_14;
  wire       [55:0]   _zz__zz_add_oh_shift_1_1;
  wire                _zz__zz_add_oh_shift_51;
  wire                _zz__zz_add_oh_shift_52;
  wire                _zz__zz_add_oh_shift_53;
  wire                _zz__zz_add_oh_shift_54;
  wire                _zz__zz_add_oh_shift_55;
  wire                _zz__zz_add_oh_shift_56;
  wire       [12:0]   _zz_add_norm_output_payload_exponent;
  wire       [12:0]   _zz_add_norm_output_payload_exponent_1;
  wire       [6:0]    _zz_add_norm_output_payload_exponent_2;
  wire       [53:0]   _zz_add_result_output_payload_value_mantissa;
  wire       [12:0]   _zz_roundFront_expDif;
  wire       [11:0]   _zz_roundFront_expDif_1;
  wire       [5:0]    _zz_roundFront_exactMask;
  wire                _zz_roundFront_exactMask_1;
  wire       [0:0]    _zz_roundFront_exactMask_2;
  wire       [46:0]   _zz_roundFront_exactMask_3;
  wire       [5:0]    _zz_roundFront_exactMask_4;
  wire                _zz_roundFront_exactMask_5;
  wire       [0:0]    _zz_roundFront_exactMask_6;
  wire       [38:0]   _zz_roundFront_exactMask_7;
  wire       [5:0]    _zz_roundFront_exactMask_8;
  wire                _zz_roundFront_exactMask_9;
  wire       [0:0]    _zz_roundFront_exactMask_10;
  wire       [30:0]   _zz_roundFront_exactMask_11;
  wire       [5:0]    _zz_roundFront_exactMask_12;
  wire                _zz_roundFront_exactMask_13;
  wire       [0:0]    _zz_roundFront_exactMask_14;
  wire       [22:0]   _zz_roundFront_exactMask_15;
  wire       [5:0]    _zz_roundFront_exactMask_16;
  wire                _zz_roundFront_exactMask_17;
  wire       [0:0]    _zz_roundFront_exactMask_18;
  wire       [14:0]   _zz_roundFront_exactMask_19;
  wire       [5:0]    _zz_roundFront_exactMask_20;
  wire                _zz_roundFront_exactMask_21;
  wire       [0:0]    _zz_roundFront_exactMask_22;
  wire       [6:0]    _zz_roundFront_exactMask_23;
  wire       [53:0]   _zz_roundFront_roundAdjusted;
  wire       [52:0]   _zz_roundFront_roundAdjusted_1;
  wire       [53:0]   _zz_roundFront_rneBit;
  wire       [51:0]   _zz_roundFront_rneBit_1;
  wire       [51:0]   _zz_roundBack_adderMantissa;
  wire       [52:0]   _zz_roundBack_adderRightOp;
  wire       [52:0]   _zz_roundBack_adderRightOp_1;
  wire       [63:0]   _zz_roundBack_adder_2;
  wire       [63:0]   _zz_roundBack_adder_3;
  wire       [63:0]   _zz_roundBack_adder_4;
  wire       [63:0]   _zz_roundBack_masked;
  wire       [51:0]   _zz_roundBack_masked_1;
  wire       [52:0]   _zz_roundBack_masked_2;
  wire       [11:0]   _zz_roundBack_borringCase;
  wire       [11:0]   _zz_when_FpuCore_l1616;
  wire       [11:0]   _zz_when_FpuCore_l1638;
  reg                 _zz_roundBack_write;
  wire       [66:0]   _zz_rf_ram_port;
  reg                 _zz_1;
  reg        [12:0]   roundFront_discardCount_1;
  reg        [54:0]   add_shifter_yMantissa_6;
  reg        [54:0]   add_shifter_yMantissa_5;
  reg        [54:0]   add_shifter_yMantissa_4;
  reg        [54:0]   add_shifter_yMantissa_3;
  reg        [54:0]   add_shifter_yMantissa_2;
  reg        [54:0]   add_shifter_yMantissa_1;
  reg        [52:0]   shortPip_fsm_shift_input_6;
  reg        [52:0]   shortPip_fsm_shift_input_5;
  reg        [52:0]   shortPip_fsm_shift_input_4;
  reg        [52:0]   shortPip_fsm_shift_input_3;
  reg        [52:0]   shortPip_fsm_shift_input_2;
  reg        [52:0]   shortPip_fsm_shift_input_1;
  reg        [51:0]   load_s1_fsm_shift_input_6;
  reg        [51:0]   load_s1_fsm_shift_input_5;
  reg        [51:0]   load_s1_fsm_shift_input_4;
  reg        [51:0]   load_s1_fsm_shift_input_3;
  reg        [51:0]   load_s1_fsm_shift_input_2;
  reg        [51:0]   load_s1_fsm_shift_input_1;
  reg                 _zz_2;
  reg                 _zz_3;
  reg                 _zz_4;
  reg                 _zz_5;
  reg                 _zz_6;
  reg                 _zz_7;
  reg        [5:0]    rf_init_counter;
  wire                rf_init_done;
  wire                when_FpuCore_l163;
  reg                 rf_scoreboards_0_targetWrite_valid;
  reg        [4:0]    rf_scoreboards_0_targetWrite_payload_address;
  reg                 rf_scoreboards_0_targetWrite_payload_data;
  reg                 rf_scoreboards_0_hitWrite_valid;
  reg        [4:0]    rf_scoreboards_0_hitWrite_payload_address;
  reg                 rf_scoreboards_0_hitWrite_payload_data;
  reg                 rf_scoreboards_1_targetWrite_valid;
  reg        [4:0]    rf_scoreboards_1_targetWrite_payload_address;
  reg                 rf_scoreboards_1_targetWrite_payload_data;
  reg                 rf_scoreboards_1_hitWrite_valid;
  reg        [4:0]    rf_scoreboards_1_hitWrite_payload_address;
  reg                 rf_scoreboards_1_hitWrite_payload_data;
  wire                commitFork_load_0_valid;
  reg                 commitFork_load_0_ready;
  wire       [3:0]    commitFork_load_0_payload_opcode;
  wire       [4:0]    commitFork_load_0_payload_rd;
  wire                commitFork_load_0_payload_write;
  wire       [63:0]   commitFork_load_0_payload_value;
  wire                commitFork_load_1_valid;
  reg                 commitFork_load_1_ready;
  wire       [3:0]    commitFork_load_1_payload_opcode;
  wire       [4:0]    commitFork_load_1_payload_rd;
  wire                commitFork_load_1_payload_write;
  wire       [63:0]   commitFork_load_1_payload_value;
  wire                commitFork_commit_0_valid;
  wire                commitFork_commit_0_ready;
  wire       [3:0]    commitFork_commit_0_payload_opcode;
  wire       [4:0]    commitFork_commit_0_payload_rd;
  wire                commitFork_commit_0_payload_write;
  wire       [63:0]   commitFork_commit_0_payload_value;
  wire                commitFork_commit_1_valid;
  wire                commitFork_commit_1_ready;
  wire       [3:0]    commitFork_commit_1_payload_opcode;
  wire       [4:0]    commitFork_commit_1_payload_rd;
  wire                commitFork_commit_1_payload_write;
  wire       [63:0]   commitFork_commit_1_payload_value;
  wire                streamFork_3_io_outputs_1_s2mPipe_valid;
  wire                streamFork_3_io_outputs_1_s2mPipe_ready;
  wire       [3:0]    streamFork_3_io_outputs_1_s2mPipe_payload_opcode;
  wire       [4:0]    streamFork_3_io_outputs_1_s2mPipe_payload_rd;
  wire                streamFork_3_io_outputs_1_s2mPipe_payload_write;
  wire       [63:0]   streamFork_3_io_outputs_1_s2mPipe_payload_value;
  reg                 streamFork_3_io_outputs_1_rValidN;
  reg        [3:0]    streamFork_3_io_outputs_1_rData_opcode;
  reg        [4:0]    streamFork_3_io_outputs_1_rData_rd;
  reg                 streamFork_3_io_outputs_1_rData_write;
  reg        [63:0]   streamFork_3_io_outputs_1_rData_value;
  wire       [3:0]    _zz_payload_opcode;
  wire                streamFork_4_io_outputs_1_s2mPipe_valid;
  wire                streamFork_4_io_outputs_1_s2mPipe_ready;
  wire       [3:0]    streamFork_4_io_outputs_1_s2mPipe_payload_opcode;
  wire       [4:0]    streamFork_4_io_outputs_1_s2mPipe_payload_rd;
  wire                streamFork_4_io_outputs_1_s2mPipe_payload_write;
  wire       [63:0]   streamFork_4_io_outputs_1_s2mPipe_payload_value;
  reg                 streamFork_4_io_outputs_1_rValidN;
  reg        [3:0]    streamFork_4_io_outputs_1_rData_opcode;
  reg        [4:0]    streamFork_4_io_outputs_1_rData_rd;
  reg                 streamFork_4_io_outputs_1_rData_write;
  reg        [63:0]   streamFork_4_io_outputs_1_rData_value;
  wire       [3:0]    _zz_payload_opcode_1;
  reg        [3:0]    commitLogic_0_pending_counter;
  wire                commitLogic_0_pending_full;
  wire                commitLogic_0_pending_notEmpty;
  reg                 commitLogic_0_pending_inc;
  reg                 commitLogic_0_pending_dec;
  reg        [3:0]    commitLogic_0_add_counter;
  wire                commitLogic_0_add_full;
  wire                commitLogic_0_add_notEmpty;
  reg                 commitLogic_0_add_inc;
  reg                 commitLogic_0_add_dec;
  reg        [3:0]    commitLogic_0_mul_counter;
  wire                commitLogic_0_mul_full;
  wire                commitLogic_0_mul_notEmpty;
  reg                 commitLogic_0_mul_inc;
  reg                 commitLogic_0_mul_dec;
  reg        [3:0]    commitLogic_0_div_counter;
  wire                commitLogic_0_div_full;
  wire                commitLogic_0_div_notEmpty;
  reg                 commitLogic_0_div_inc;
  reg                 commitLogic_0_div_dec;
  reg        [3:0]    commitLogic_0_sqrt_counter;
  wire                commitLogic_0_sqrt_full;
  wire                commitLogic_0_sqrt_notEmpty;
  reg                 commitLogic_0_sqrt_inc;
  reg                 commitLogic_0_sqrt_dec;
  reg        [3:0]    commitLogic_0_short_counter;
  wire                commitLogic_0_short_full;
  wire                commitLogic_0_short_notEmpty;
  reg                 commitLogic_0_short_inc;
  reg                 commitLogic_0_short_dec;
  wire                _zz_commitFork_commit_0_ready;
  wire       [3:0]    _zz_commitLogic_0_input_payload_opcode;
  wire                commitLogic_0_input_valid;
  wire       [3:0]    commitLogic_0_input_payload_opcode;
  wire       [4:0]    commitLogic_0_input_payload_rd;
  wire                commitLogic_0_input_payload_write;
  wire       [63:0]   commitLogic_0_input_payload_value;
  wire                when_FpuCore_l208;
  wire                when_FpuCore_l209;
  wire                when_FpuCore_l210;
  wire                when_FpuCore_l211;
  wire                when_FpuCore_l212;
  reg        [3:0]    commitLogic_1_pending_counter;
  wire                commitLogic_1_pending_full;
  wire                commitLogic_1_pending_notEmpty;
  reg                 commitLogic_1_pending_inc;
  reg                 commitLogic_1_pending_dec;
  reg        [3:0]    commitLogic_1_add_counter;
  wire                commitLogic_1_add_full;
  wire                commitLogic_1_add_notEmpty;
  reg                 commitLogic_1_add_inc;
  reg                 commitLogic_1_add_dec;
  reg        [3:0]    commitLogic_1_mul_counter;
  wire                commitLogic_1_mul_full;
  wire                commitLogic_1_mul_notEmpty;
  reg                 commitLogic_1_mul_inc;
  reg                 commitLogic_1_mul_dec;
  reg        [3:0]    commitLogic_1_div_counter;
  wire                commitLogic_1_div_full;
  wire                commitLogic_1_div_notEmpty;
  reg                 commitLogic_1_div_inc;
  reg                 commitLogic_1_div_dec;
  reg        [3:0]    commitLogic_1_sqrt_counter;
  wire                commitLogic_1_sqrt_full;
  wire                commitLogic_1_sqrt_notEmpty;
  reg                 commitLogic_1_sqrt_inc;
  reg                 commitLogic_1_sqrt_dec;
  reg        [3:0]    commitLogic_1_short_counter;
  wire                commitLogic_1_short_full;
  wire                commitLogic_1_short_notEmpty;
  reg                 commitLogic_1_short_inc;
  reg                 commitLogic_1_short_dec;
  wire                _zz_commitFork_commit_1_ready;
  wire       [3:0]    _zz_commitLogic_1_input_payload_opcode;
  wire                commitLogic_1_input_valid;
  wire       [3:0]    commitLogic_1_input_payload_opcode;
  wire       [4:0]    commitLogic_1_input_payload_rd;
  wire                commitLogic_1_input_payload_write;
  wire       [63:0]   commitLogic_1_input_payload_value;
  wire                when_FpuCore_l208_1;
  wire                when_FpuCore_l209_1;
  wire                when_FpuCore_l210_1;
  wire                when_FpuCore_l211_1;
  wire                when_FpuCore_l212_1;
  wire                scheduler_0_input_valid;
  wire                scheduler_0_input_ready;
  wire       [3:0]    scheduler_0_input_payload_opcode;
  wire       [1:0]    scheduler_0_input_payload_arg;
  wire       [4:0]    scheduler_0_input_payload_rs1;
  wire       [4:0]    scheduler_0_input_payload_rs2;
  wire       [4:0]    scheduler_0_input_payload_rs3;
  wire       [4:0]    scheduler_0_input_payload_rd;
  wire       [0:0]    scheduler_0_input_payload_format;
  wire       [2:0]    scheduler_0_input_payload_roundMode;
  reg                 io_port_0_cmd_rValidN;
  reg        [3:0]    io_port_0_cmd_rData_opcode;
  reg        [1:0]    io_port_0_cmd_rData_arg;
  reg        [4:0]    io_port_0_cmd_rData_rs1;
  reg        [4:0]    io_port_0_cmd_rData_rs2;
  reg        [4:0]    io_port_0_cmd_rData_rs3;
  reg        [4:0]    io_port_0_cmd_rData_rd;
  reg        [0:0]    io_port_0_cmd_rData_format;
  reg        [2:0]    io_port_0_cmd_rData_roundMode;
  wire       [3:0]    _zz_scheduler_0_input_payload_opcode;
  wire       [0:0]    _zz_scheduler_0_input_payload_format;
  wire       [2:0]    _zz_scheduler_0_input_payload_roundMode;
  reg                 scheduler_0_useRs1;
  reg                 scheduler_0_useRs2;
  reg                 scheduler_0_useRs3;
  reg                 scheduler_0_useRd;
  wire                scheduler_0_rfHits_0;
  wire                scheduler_0_rfHits_1;
  wire                scheduler_0_rfHits_2;
  wire                scheduler_0_rfHits_3;
  wire                scheduler_0_rfTargets_0;
  wire                scheduler_0_rfTargets_1;
  wire                scheduler_0_rfTargets_2;
  wire                scheduler_0_rfTargets_3;
  wire                scheduler_0_rfBusy_0;
  wire                scheduler_0_rfBusy_1;
  wire                scheduler_0_rfBusy_2;
  wire                scheduler_0_rfBusy_3;
  wire                scheduler_0_hits_0;
  wire                scheduler_0_hits_1;
  wire                scheduler_0_hits_2;
  wire                scheduler_0_hits_3;
  wire                scheduler_0_hazard;
  wire                _zz_scheduler_0_input_ready;
  wire                scheduler_0_output_valid;
  reg                 scheduler_0_output_ready;
  wire       [3:0]    scheduler_0_output_payload_opcode;
  wire       [1:0]    scheduler_0_output_payload_arg;
  reg        [4:0]    scheduler_0_output_payload_rs1;
  wire       [4:0]    scheduler_0_output_payload_rs2;
  wire       [4:0]    scheduler_0_output_payload_rs3;
  wire       [4:0]    scheduler_0_output_payload_rd;
  wire       [0:0]    scheduler_0_output_payload_format;
  wire       [2:0]    scheduler_0_output_payload_roundMode;
  wire                when_FpuCore_l258;
  wire                when_FpuCore_l261;
  wire                scheduler_0_output_fire;
  wire                when_FpuCore_l265;
  wire                scheduler_1_input_valid;
  wire                scheduler_1_input_ready;
  wire       [3:0]    scheduler_1_input_payload_opcode;
  wire       [1:0]    scheduler_1_input_payload_arg;
  wire       [4:0]    scheduler_1_input_payload_rs1;
  wire       [4:0]    scheduler_1_input_payload_rs2;
  wire       [4:0]    scheduler_1_input_payload_rs3;
  wire       [4:0]    scheduler_1_input_payload_rd;
  wire       [0:0]    scheduler_1_input_payload_format;
  wire       [2:0]    scheduler_1_input_payload_roundMode;
  reg                 io_port_1_cmd_rValidN;
  reg        [3:0]    io_port_1_cmd_rData_opcode;
  reg        [1:0]    io_port_1_cmd_rData_arg;
  reg        [4:0]    io_port_1_cmd_rData_rs1;
  reg        [4:0]    io_port_1_cmd_rData_rs2;
  reg        [4:0]    io_port_1_cmd_rData_rs3;
  reg        [4:0]    io_port_1_cmd_rData_rd;
  reg        [0:0]    io_port_1_cmd_rData_format;
  reg        [2:0]    io_port_1_cmd_rData_roundMode;
  wire       [3:0]    _zz_scheduler_1_input_payload_opcode;
  wire       [0:0]    _zz_scheduler_1_input_payload_format;
  wire       [2:0]    _zz_scheduler_1_input_payload_roundMode;
  reg                 scheduler_1_useRs1;
  reg                 scheduler_1_useRs2;
  reg                 scheduler_1_useRs3;
  reg                 scheduler_1_useRd;
  wire                scheduler_1_rfHits_0;
  wire                scheduler_1_rfHits_1;
  wire                scheduler_1_rfHits_2;
  wire                scheduler_1_rfHits_3;
  wire                scheduler_1_rfTargets_0;
  wire                scheduler_1_rfTargets_1;
  wire                scheduler_1_rfTargets_2;
  wire                scheduler_1_rfTargets_3;
  wire                scheduler_1_rfBusy_0;
  wire                scheduler_1_rfBusy_1;
  wire                scheduler_1_rfBusy_2;
  wire                scheduler_1_rfBusy_3;
  wire                scheduler_1_hits_0;
  wire                scheduler_1_hits_1;
  wire                scheduler_1_hits_2;
  wire                scheduler_1_hits_3;
  wire                scheduler_1_hazard;
  wire                _zz_scheduler_1_input_ready;
  wire                scheduler_1_output_valid;
  reg                 scheduler_1_output_ready;
  wire       [3:0]    scheduler_1_output_payload_opcode;
  wire       [1:0]    scheduler_1_output_payload_arg;
  reg        [4:0]    scheduler_1_output_payload_rs1;
  wire       [4:0]    scheduler_1_output_payload_rs2;
  wire       [4:0]    scheduler_1_output_payload_rs3;
  wire       [4:0]    scheduler_1_output_payload_rd;
  wire       [0:0]    scheduler_1_output_payload_format;
  wire       [2:0]    scheduler_1_output_payload_roundMode;
  wire                when_FpuCore_l258_1;
  wire                when_FpuCore_l261_1;
  wire                scheduler_1_output_fire;
  wire                when_FpuCore_l265_1;
  wire                scheduler_0_output_m2sPipe_valid;
  wire                scheduler_0_output_m2sPipe_ready;
  wire       [3:0]    scheduler_0_output_m2sPipe_payload_opcode;
  wire       [1:0]    scheduler_0_output_m2sPipe_payload_arg;
  wire       [4:0]    scheduler_0_output_m2sPipe_payload_rs1;
  wire       [4:0]    scheduler_0_output_m2sPipe_payload_rs2;
  wire       [4:0]    scheduler_0_output_m2sPipe_payload_rs3;
  wire       [4:0]    scheduler_0_output_m2sPipe_payload_rd;
  wire       [0:0]    scheduler_0_output_m2sPipe_payload_format;
  wire       [2:0]    scheduler_0_output_m2sPipe_payload_roundMode;
  reg                 scheduler_0_output_rValid;
  reg        [3:0]    scheduler_0_output_rData_opcode;
  reg        [1:0]    scheduler_0_output_rData_arg;
  reg        [4:0]    scheduler_0_output_rData_rs1;
  reg        [4:0]    scheduler_0_output_rData_rs2;
  reg        [4:0]    scheduler_0_output_rData_rs3;
  reg        [4:0]    scheduler_0_output_rData_rd;
  reg        [0:0]    scheduler_0_output_rData_format;
  reg        [2:0]    scheduler_0_output_rData_roundMode;
  wire                when_Stream_l375;
  wire                scheduler_1_output_m2sPipe_valid;
  wire                scheduler_1_output_m2sPipe_ready;
  wire       [3:0]    scheduler_1_output_m2sPipe_payload_opcode;
  wire       [1:0]    scheduler_1_output_m2sPipe_payload_arg;
  wire       [4:0]    scheduler_1_output_m2sPipe_payload_rs1;
  wire       [4:0]    scheduler_1_output_m2sPipe_payload_rs2;
  wire       [4:0]    scheduler_1_output_m2sPipe_payload_rs3;
  wire       [4:0]    scheduler_1_output_m2sPipe_payload_rd;
  wire       [0:0]    scheduler_1_output_m2sPipe_payload_format;
  wire       [2:0]    scheduler_1_output_m2sPipe_payload_roundMode;
  reg                 scheduler_1_output_rValid;
  reg        [3:0]    scheduler_1_output_rData_opcode;
  reg        [1:0]    scheduler_1_output_rData_arg;
  reg        [4:0]    scheduler_1_output_rData_rs1;
  reg        [4:0]    scheduler_1_output_rData_rs2;
  reg        [4:0]    scheduler_1_output_rData_rs3;
  reg        [4:0]    scheduler_1_output_rData_rd;
  reg        [0:0]    scheduler_1_output_rData_format;
  reg        [2:0]    scheduler_1_output_rData_roundMode;
  wire                when_Stream_l375_1;
  wire                cmdArbiter_output_valid;
  wire                cmdArbiter_output_ready;
  wire       [0:0]    cmdArbiter_output_payload_source;
  wire       [3:0]    cmdArbiter_output_payload_opcode;
  wire       [4:0]    cmdArbiter_output_payload_rs1;
  wire       [4:0]    cmdArbiter_output_payload_rs2;
  wire       [4:0]    cmdArbiter_output_payload_rs3;
  wire       [4:0]    cmdArbiter_output_payload_rd;
  wire       [1:0]    cmdArbiter_output_payload_arg;
  wire       [2:0]    cmdArbiter_output_payload_roundMode;
  wire       [0:0]    cmdArbiter_output_payload_format;
  wire                read_s0_valid;
  reg                 read_s0_ready;
  wire       [0:0]    read_s0_payload_source;
  wire       [3:0]    read_s0_payload_opcode;
  wire       [4:0]    read_s0_payload_rs1;
  wire       [4:0]    read_s0_payload_rs2;
  wire       [4:0]    read_s0_payload_rs3;
  wire       [4:0]    read_s0_payload_rd;
  wire       [1:0]    read_s0_payload_arg;
  wire       [2:0]    read_s0_payload_roundMode;
  wire       [0:0]    read_s0_payload_format;
  wire                read_s1_valid;
  wire                read_s1_ready;
  wire       [0:0]    read_s1_payload_source;
  wire       [3:0]    read_s1_payload_opcode;
  wire       [4:0]    read_s1_payload_rs1;
  wire       [4:0]    read_s1_payload_rs2;
  wire       [4:0]    read_s1_payload_rs3;
  wire       [4:0]    read_s1_payload_rd;
  wire       [1:0]    read_s1_payload_arg;
  wire       [2:0]    read_s1_payload_roundMode;
  wire       [0:0]    read_s1_payload_format;
  reg                 read_s0_rValid;
  reg        [0:0]    read_s0_rData_source;
  reg        [3:0]    read_s0_rData_opcode;
  reg        [4:0]    read_s0_rData_rs1;
  reg        [4:0]    read_s0_rData_rs2;
  reg        [4:0]    read_s0_rData_rs3;
  reg        [4:0]    read_s0_rData_rd;
  reg        [1:0]    read_s0_rData_arg;
  reg        [2:0]    read_s0_rData_roundMode;
  reg        [0:0]    read_s0_rData_format;
  wire                when_Stream_l375_2;
  wire                read_output_valid;
  wire                read_output_ready;
  wire       [0:0]    read_output_payload_source;
  wire       [3:0]    read_output_payload_opcode;
  reg        [51:0]   read_output_payload_rs1_mantissa;
  reg        [11:0]   read_output_payload_rs1_exponent;
  reg                 read_output_payload_rs1_sign;
  reg                 read_output_payload_rs1_special;
  reg        [51:0]   read_output_payload_rs2_mantissa;
  reg        [11:0]   read_output_payload_rs2_exponent;
  reg                 read_output_payload_rs2_sign;
  reg                 read_output_payload_rs2_special;
  reg        [51:0]   read_output_payload_rs3_mantissa;
  reg        [11:0]   read_output_payload_rs3_exponent;
  wire                read_output_payload_rs3_sign;
  reg                 read_output_payload_rs3_special;
  wire       [4:0]    read_output_payload_rd;
  wire       [1:0]    read_output_payload_arg;
  wire       [2:0]    read_output_payload_roundMode;
  reg        [0:0]    read_output_payload_format;
  wire                read_output_payload_rs1Boxed;
  wire                read_output_payload_rs2Boxed;
  wire       [5:0]    _zz_read_rs_0_boxed;
  wire                read_output_isStall;
  wire                _zz_read_rs_0_boxed_1;
  wire       [51:0]   read_rs_0_value_mantissa;
  wire       [11:0]   read_rs_0_value_exponent;
  wire                read_rs_0_value_sign;
  wire                read_rs_0_value_special;
  wire                read_rs_0_boxed;
  wire       [66:0]   _zz_read_rs_0_boxed_2;
  wire       [65:0]   _zz_read_rs_0_value_mantissa;
  wire       [5:0]    _zz_read_rs_1_boxed;
  wire                _zz_read_rs_1_boxed_1;
  wire       [51:0]   read_rs_1_value_mantissa;
  wire       [11:0]   read_rs_1_value_exponent;
  wire                read_rs_1_value_sign;
  wire                read_rs_1_value_special;
  wire                read_rs_1_boxed;
  wire       [66:0]   _zz_read_rs_1_boxed_2;
  wire       [65:0]   _zz_read_rs_1_value_mantissa;
  wire       [5:0]    _zz_read_rs_2_boxed;
  wire                _zz_read_rs_2_boxed_1;
  wire       [51:0]   read_rs_2_value_mantissa;
  wire       [11:0]   read_rs_2_value_exponent;
  wire                read_rs_2_value_sign;
  wire                read_rs_2_value_special;
  wire                read_rs_2_boxed;
  wire       [66:0]   _zz_read_rs_2_boxed_2;
  wire       [65:0]   _zz_read_rs_2_value_mantissa;
  wire                when_FpuCore_l305;
  wire                when_FpuCore_l304;
  wire       [0:0]    _zz_read_output_payload_format;
  wire                when_FpuCore_l307;
  wire                when_FpuCore_l312;
  wire                when_FpuCore_l316;
  wire                decode_input_valid;
  reg                 decode_input_ready;
  wire       [0:0]    decode_input_payload_source;
  wire       [3:0]    decode_input_payload_opcode;
  wire       [51:0]   decode_input_payload_rs1_mantissa;
  wire       [11:0]   decode_input_payload_rs1_exponent;
  wire                decode_input_payload_rs1_sign;
  wire                decode_input_payload_rs1_special;
  wire       [51:0]   decode_input_payload_rs2_mantissa;
  wire       [11:0]   decode_input_payload_rs2_exponent;
  wire                decode_input_payload_rs2_sign;
  wire                decode_input_payload_rs2_special;
  wire       [51:0]   decode_input_payload_rs3_mantissa;
  wire       [11:0]   decode_input_payload_rs3_exponent;
  wire                decode_input_payload_rs3_sign;
  wire                decode_input_payload_rs3_special;
  wire       [4:0]    decode_input_payload_rd;
  wire       [1:0]    decode_input_payload_arg;
  wire       [2:0]    decode_input_payload_roundMode;
  wire       [0:0]    decode_input_payload_format;
  wire                decode_input_payload_rs1Boxed;
  wire                decode_input_payload_rs2Boxed;
  wire                decode_loadHit;
  wire                decode_load_valid;
  wire                decode_load_ready;
  wire       [0:0]    decode_load_payload_source;
  wire       [4:0]    decode_load_payload_rd;
  wire                decode_load_payload_i2f;
  wire       [1:0]    decode_load_payload_arg;
  wire       [2:0]    decode_load_payload_roundMode;
  wire       [0:0]    decode_load_payload_format;
  wire                when_FpuCore_l329;
  wire                decode_shortPipHit;
  wire                decode_shortPip_valid;
  reg                 decode_shortPip_ready;
  wire       [0:0]    decode_shortPip_payload_source;
  wire       [3:0]    decode_shortPip_payload_opcode;
  wire       [51:0]   decode_shortPip_payload_rs1_mantissa;
  wire       [11:0]   decode_shortPip_payload_rs1_exponent;
  wire                decode_shortPip_payload_rs1_sign;
  wire                decode_shortPip_payload_rs1_special;
  wire       [51:0]   decode_shortPip_payload_rs2_mantissa;
  wire       [11:0]   decode_shortPip_payload_rs2_exponent;
  wire                decode_shortPip_payload_rs2_sign;
  wire                decode_shortPip_payload_rs2_special;
  wire       [4:0]    decode_shortPip_payload_rd;
  wire       [31:0]   decode_shortPip_payload_value;
  wire       [1:0]    decode_shortPip_payload_arg;
  wire       [2:0]    decode_shortPip_payload_roundMode;
  wire       [0:0]    decode_shortPip_payload_format;
  wire                decode_shortPip_payload_rs1Boxed;
  wire                decode_shortPip_payload_rs2Boxed;
  wire                when_FpuCore_l335;
  wire                decode_divSqrtHit;
  wire                decode_divSqrt_valid;
  wire                decode_divSqrt_ready;
  wire       [0:0]    decode_divSqrt_payload_source;
  wire       [51:0]   decode_divSqrt_payload_rs1_mantissa;
  wire       [11:0]   decode_divSqrt_payload_rs1_exponent;
  wire                decode_divSqrt_payload_rs1_sign;
  wire                decode_divSqrt_payload_rs1_special;
  wire       [51:0]   decode_divSqrt_payload_rs2_mantissa;
  wire       [11:0]   decode_divSqrt_payload_rs2_exponent;
  wire                decode_divSqrt_payload_rs2_sign;
  wire                decode_divSqrt_payload_rs2_special;
  wire       [4:0]    decode_divSqrt_payload_rd;
  wire                decode_divSqrt_payload_div;
  wire       [2:0]    decode_divSqrt_payload_roundMode;
  wire       [0:0]    decode_divSqrt_payload_format;
  wire                decode_divHit;
  wire                decode_div_valid;
  wire                decode_div_ready;
  wire       [0:0]    decode_div_payload_source;
  wire       [51:0]   decode_div_payload_rs1_mantissa;
  wire       [11:0]   decode_div_payload_rs1_exponent;
  wire                decode_div_payload_rs1_sign;
  wire                decode_div_payload_rs1_special;
  wire       [51:0]   decode_div_payload_rs2_mantissa;
  wire       [11:0]   decode_div_payload_rs2_exponent;
  wire                decode_div_payload_rs2_sign;
  wire                decode_div_payload_rs2_special;
  wire       [4:0]    decode_div_payload_rd;
  wire       [2:0]    decode_div_payload_roundMode;
  wire       [0:0]    decode_div_payload_format;
  wire                when_FpuCore_l351;
  wire                decode_sqrtHit;
  wire                decode_sqrt_valid;
  wire                decode_sqrt_ready;
  wire       [0:0]    decode_sqrt_payload_source;
  wire       [51:0]   decode_sqrt_payload_rs1_mantissa;
  wire       [11:0]   decode_sqrt_payload_rs1_exponent;
  wire                decode_sqrt_payload_rs1_sign;
  wire                decode_sqrt_payload_rs1_special;
  wire       [4:0]    decode_sqrt_payload_rd;
  wire       [2:0]    decode_sqrt_payload_roundMode;
  wire       [0:0]    decode_sqrt_payload_format;
  wire                when_FpuCore_l359;
  wire                decode_fmaHit;
  wire                decode_mulHit;
  wire                decode_mul_valid;
  reg                 decode_mul_ready;
  reg        [0:0]    decode_mul_payload_source;
  reg        [51:0]   decode_mul_payload_rs1_mantissa;
  reg        [11:0]   decode_mul_payload_rs1_exponent;
  reg                 decode_mul_payload_rs1_sign;
  reg                 decode_mul_payload_rs1_special;
  reg        [51:0]   decode_mul_payload_rs2_mantissa;
  reg        [11:0]   decode_mul_payload_rs2_exponent;
  reg                 decode_mul_payload_rs2_sign;
  reg                 decode_mul_payload_rs2_special;
  reg        [51:0]   decode_mul_payload_rs3_mantissa;
  reg        [11:0]   decode_mul_payload_rs3_exponent;
  reg                 decode_mul_payload_rs3_sign;
  reg                 decode_mul_payload_rs3_special;
  reg        [4:0]    decode_mul_payload_rd;
  reg                 decode_mul_payload_add;
  reg                 decode_mul_payload_divSqrt;
  reg                 decode_mul_payload_msb1;
  reg                 decode_mul_payload_msb2;
  reg        [2:0]    decode_mul_payload_roundMode;
  reg        [0:0]    decode_mul_payload_format;
  wire                decode_divSqrtToMul_valid;
  wire                decode_divSqrtToMul_ready;
  wire       [0:0]    decode_divSqrtToMul_payload_source;
  wire       [51:0]   decode_divSqrtToMul_payload_rs1_mantissa;
  wire       [11:0]   decode_divSqrtToMul_payload_rs1_exponent;
  wire                decode_divSqrtToMul_payload_rs1_sign;
  wire                decode_divSqrtToMul_payload_rs1_special;
  wire       [51:0]   decode_divSqrtToMul_payload_rs2_mantissa;
  wire       [11:0]   decode_divSqrtToMul_payload_rs2_exponent;
  wire                decode_divSqrtToMul_payload_rs2_sign;
  wire                decode_divSqrtToMul_payload_rs2_special;
  wire       [51:0]   decode_divSqrtToMul_payload_rs3_mantissa;
  wire       [11:0]   decode_divSqrtToMul_payload_rs3_exponent;
  wire                decode_divSqrtToMul_payload_rs3_sign;
  wire                decode_divSqrtToMul_payload_rs3_special;
  wire       [4:0]    decode_divSqrtToMul_payload_rd;
  wire                decode_divSqrtToMul_payload_add;
  wire                decode_divSqrtToMul_payload_divSqrt;
  wire                decode_divSqrtToMul_payload_msb1;
  wire                decode_divSqrtToMul_payload_msb2;
  wire       [2:0]    decode_divSqrtToMul_payload_roundMode;
  wire       [0:0]    decode_divSqrtToMul_payload_format;
  wire                when_FpuCore_l375;
  wire                when_FpuCore_l380;
  wire                decode_addHit;
  wire                decode_add_valid;
  wire                decode_add_ready;
  reg        [0:0]    decode_add_payload_source;
  reg        [53:0]   decode_add_payload_rs1_mantissa;
  reg        [11:0]   decode_add_payload_rs1_exponent;
  reg                 decode_add_payload_rs1_sign;
  reg                 decode_add_payload_rs1_special;
  reg        [53:0]   decode_add_payload_rs2_mantissa;
  reg        [11:0]   decode_add_payload_rs2_exponent;
  reg                 decode_add_payload_rs2_sign;
  reg                 decode_add_payload_rs2_special;
  reg        [4:0]    decode_add_payload_rd;
  reg        [2:0]    decode_add_payload_roundMode;
  reg        [0:0]    decode_add_payload_format;
  reg                 decode_add_payload_needCommit;
  wire                decode_mulToAdd_valid;
  wire                decode_mulToAdd_ready;
  wire       [0:0]    decode_mulToAdd_payload_source;
  wire       [53:0]   decode_mulToAdd_payload_rs1_mantissa;
  wire       [11:0]   decode_mulToAdd_payload_rs1_exponent;
  wire                decode_mulToAdd_payload_rs1_sign;
  wire                decode_mulToAdd_payload_rs1_special;
  wire       [53:0]   decode_mulToAdd_payload_rs2_mantissa;
  wire       [11:0]   decode_mulToAdd_payload_rs2_exponent;
  wire                decode_mulToAdd_payload_rs2_sign;
  wire                decode_mulToAdd_payload_rs2_special;
  wire       [4:0]    decode_mulToAdd_payload_rd;
  wire       [2:0]    decode_mulToAdd_payload_roundMode;
  wire       [0:0]    decode_mulToAdd_payload_format;
  wire                decode_mulToAdd_payload_needCommit;
  wire                when_FpuCore_l399;
  wire                when_FpuCore_l404;
  wire                decode_load_s2mPipe_valid;
  reg                 decode_load_s2mPipe_ready;
  wire       [0:0]    decode_load_s2mPipe_payload_source;
  wire       [4:0]    decode_load_s2mPipe_payload_rd;
  wire                decode_load_s2mPipe_payload_i2f;
  wire       [1:0]    decode_load_s2mPipe_payload_arg;
  wire       [2:0]    decode_load_s2mPipe_payload_roundMode;
  wire       [0:0]    decode_load_s2mPipe_payload_format;
  reg                 decode_load_rValidN;
  reg        [0:0]    decode_load_rData_source;
  reg        [4:0]    decode_load_rData_rd;
  reg                 decode_load_rData_i2f;
  reg        [1:0]    decode_load_rData_arg;
  reg        [2:0]    decode_load_rData_roundMode;
  reg        [0:0]    decode_load_rData_format;
  wire       [2:0]    _zz_decode_load_s2mPipe_payload_roundMode;
  wire       [0:0]    _zz_decode_load_s2mPipe_payload_format;
  wire                decode_load_s2mPipe_m2sPipe_valid;
  reg                 decode_load_s2mPipe_m2sPipe_ready;
  wire       [0:0]    decode_load_s2mPipe_m2sPipe_payload_source;
  wire       [4:0]    decode_load_s2mPipe_m2sPipe_payload_rd;
  wire                decode_load_s2mPipe_m2sPipe_payload_i2f;
  wire       [1:0]    decode_load_s2mPipe_m2sPipe_payload_arg;
  wire       [2:0]    decode_load_s2mPipe_m2sPipe_payload_roundMode;
  wire       [0:0]    decode_load_s2mPipe_m2sPipe_payload_format;
  reg                 decode_load_s2mPipe_rValid;
  reg        [0:0]    decode_load_s2mPipe_rData_source;
  reg        [4:0]    decode_load_s2mPipe_rData_rd;
  reg                 decode_load_s2mPipe_rData_i2f;
  reg        [1:0]    decode_load_s2mPipe_rData_arg;
  reg        [2:0]    decode_load_s2mPipe_rData_roundMode;
  reg        [0:0]    decode_load_s2mPipe_rData_format;
  wire                when_Stream_l375_3;
  wire                load_s0_input_valid;
  wire                load_s0_input_ready;
  wire       [0:0]    load_s0_input_payload_source;
  wire       [4:0]    load_s0_input_payload_rd;
  wire                load_s0_input_payload_i2f;
  wire       [1:0]    load_s0_input_payload_arg;
  wire       [2:0]    load_s0_input_payload_roundMode;
  wire       [0:0]    load_s0_input_payload_format;
  reg                 decode_load_s2mPipe_m2sPipe_rValid;
  reg        [0:0]    decode_load_s2mPipe_m2sPipe_rData_source;
  reg        [4:0]    decode_load_s2mPipe_m2sPipe_rData_rd;
  reg                 decode_load_s2mPipe_m2sPipe_rData_i2f;
  reg        [1:0]    decode_load_s2mPipe_m2sPipe_rData_arg;
  reg        [2:0]    decode_load_s2mPipe_m2sPipe_rData_roundMode;
  reg        [0:0]    decode_load_s2mPipe_m2sPipe_rData_format;
  wire                when_Stream_l375_4;
  wire                when_Stream_l445;
  reg                 load_s0_filtred_0_valid;
  reg                 load_s0_filtred_0_ready;
  wire       [3:0]    load_s0_filtred_0_payload_opcode;
  wire       [4:0]    load_s0_filtred_0_payload_rd;
  wire                load_s0_filtred_0_payload_write;
  wire       [63:0]   load_s0_filtred_0_payload_value;
  wire                when_Stream_l445_1;
  reg                 load_s0_filtred_1_valid;
  reg                 load_s0_filtred_1_ready;
  wire       [3:0]    load_s0_filtred_1_payload_opcode;
  wire       [4:0]    load_s0_filtred_1_payload_rd;
  wire                load_s0_filtred_1_payload_write;
  wire       [63:0]   load_s0_filtred_1_payload_value;
  wire                load_s0_hazard;
  wire                _zz_load_s0_input_ready;
  wire                load_s0_output_valid;
  reg                 load_s0_output_ready;
  wire       [0:0]    load_s0_output_payload_source;
  wire       [4:0]    load_s0_output_payload_rd;
  wire       [63:0]   load_s0_output_payload_value;
  wire                load_s0_output_payload_i2f;
  wire       [1:0]    load_s0_output_payload_arg;
  wire       [2:0]    load_s0_output_payload_roundMode;
  reg        [0:0]    load_s0_output_payload_format;
  wire       [1:0]    _zz_33;
  wire                _zz_load_s0_filtred_0_ready;
  wire                when_FpuCore_l452;
  wire                load_s1_input_valid;
  wire                load_s1_input_ready;
  wire       [0:0]    load_s1_input_payload_source;
  wire       [4:0]    load_s1_input_payload_rd;
  wire       [63:0]   load_s1_input_payload_value;
  wire                load_s1_input_payload_i2f;
  wire       [1:0]    load_s1_input_payload_arg;
  wire       [2:0]    load_s1_input_payload_roundMode;
  wire       [0:0]    load_s1_input_payload_format;
  reg                 load_s0_output_rValid;
  reg        [0:0]    load_s0_output_rData_source;
  reg        [4:0]    load_s0_output_rData_rd;
  reg        [63:0]   load_s0_output_rData_value;
  reg                 load_s0_output_rData_i2f;
  reg        [1:0]    load_s0_output_rData_arg;
  reg        [2:0]    load_s0_output_rData_roundMode;
  reg        [0:0]    load_s0_output_rData_format;
  wire                when_Stream_l375_5;
  reg                 load_s1_busy;
  wire       [22:0]   load_s1_f32_mantissa;
  wire       [7:0]    load_s1_f32_exponent;
  wire                load_s1_f32_sign;
  wire       [51:0]   load_s1_f64_mantissa;
  wire       [10:0]   load_s1_f64_exponent;
  wire                load_s1_f64_sign;
  reg        [11:0]   load_s1_recodedExpOffset;
  reg        [51:0]   load_s1_passThroughFloat_mantissa;
  reg        [11:0]   load_s1_passThroughFloat_exponent;
  reg                 load_s1_passThroughFloat_sign;
  wire                load_s1_passThroughFloat_special;
  wire                when_FpuCore_l31;
  wire                load_s1_manZero;
  reg                 load_s1_expZero;
  reg                 load_s1_expOne;
  wire                when_FpuCore_l494;
  wire                when_FpuCore_l495;
  wire                load_s1_isZero;
  wire                load_s1_isSubnormal;
  wire                load_s1_isInfinity;
  wire                load_s1_isNan;
  reg                 load_s1_fsm_done;
  reg                 load_s1_fsm_boot;
  reg                 load_s1_fsm_patched;
  reg        [51:0]   load_s1_fsm_ohInput;
  wire                when_FpuCore_l508;
  reg                 load_s1_fsm_i2fZero;
  reg        [5:0]    load_s1_fsm_shift_by;
  reg        [51:0]   load_s1_fsm_shift_input;
  wire                when_FpuCore_l525;
  reg        [51:0]   load_s1_fsm_shift_output;
  wire                when_FpuCore_l529;
  wire                when_FpuCore_l532;
  wire       [63:0]   _zz_load_s0_output_rData_value;
  wire                _zz_load_s0_output_rData_value_1;
  wire       [51:0]   _zz_load_s1_fsm_shift_by;
  wire       [51:0]   _zz_load_s1_fsm_shift_by_1;
  wire                _zz_load_s1_fsm_shift_by_2;
  wire                _zz_load_s1_fsm_shift_by_3;
  wire                _zz_load_s1_fsm_shift_by_4;
  wire                _zz_load_s1_fsm_shift_by_5;
  wire                _zz_load_s1_fsm_shift_by_6;
  wire                _zz_load_s1_fsm_shift_by_7;
  wire                _zz_load_s1_fsm_shift_by_8;
  wire                _zz_load_s1_fsm_shift_by_9;
  wire                _zz_load_s1_fsm_shift_by_10;
  wire                _zz_load_s1_fsm_shift_by_11;
  wire                _zz_load_s1_fsm_shift_by_12;
  wire                _zz_load_s1_fsm_shift_by_13;
  wire                _zz_load_s1_fsm_shift_by_14;
  wire                _zz_load_s1_fsm_shift_by_15;
  wire                _zz_load_s1_fsm_shift_by_16;
  wire                _zz_load_s1_fsm_shift_by_17;
  wire                _zz_load_s1_fsm_shift_by_18;
  wire                _zz_load_s1_fsm_shift_by_19;
  wire                _zz_load_s1_fsm_shift_by_20;
  wire                _zz_load_s1_fsm_shift_by_21;
  wire                _zz_load_s1_fsm_shift_by_22;
  wire                _zz_load_s1_fsm_shift_by_23;
  wire                _zz_load_s1_fsm_shift_by_24;
  wire                _zz_load_s1_fsm_shift_by_25;
  wire                _zz_load_s1_fsm_shift_by_26;
  wire                _zz_load_s1_fsm_shift_by_27;
  wire                _zz_load_s1_fsm_shift_by_28;
  wire                _zz_load_s1_fsm_shift_by_29;
  wire                _zz_load_s1_fsm_shift_by_30;
  wire                _zz_load_s1_fsm_shift_by_31;
  wire                _zz_load_s1_fsm_shift_by_32;
  wire                _zz_load_s1_fsm_shift_by_33;
  wire                _zz_load_s1_fsm_shift_by_34;
  wire                _zz_load_s1_fsm_shift_by_35;
  wire                _zz_load_s1_fsm_shift_by_36;
  wire                _zz_load_s1_fsm_shift_by_37;
  wire                _zz_load_s1_fsm_shift_by_38;
  wire                _zz_load_s1_fsm_shift_by_39;
  wire                _zz_load_s1_fsm_shift_by_40;
  wire                _zz_load_s1_fsm_shift_by_41;
  wire                _zz_load_s1_fsm_shift_by_42;
  wire                _zz_load_s1_fsm_shift_by_43;
  wire                _zz_load_s1_fsm_shift_by_44;
  wire                _zz_load_s1_fsm_shift_by_45;
  wire                _zz_load_s1_fsm_shift_by_46;
  wire                _zz_load_s1_fsm_shift_by_47;
  wire                _zz_load_s1_fsm_shift_by_48;
  wire                _zz_load_s1_fsm_shift_by_49;
  wire                _zz_load_s1_fsm_shift_by_50;
  wire                _zz_load_s1_fsm_shift_by_51;
  wire                _zz_load_s1_fsm_shift_by_52;
  reg        [11:0]   load_s1_fsm_expOffset;
  wire                load_s1_input_isStall;
  wire                when_FpuCore_l551;
  wire       [51:0]   load_s1_i2fHigh;
  wire                load_s1_scrap;
  wire       [51:0]   load_s1_recoded_mantissa;
  reg        [11:0]   load_s1_recoded_exponent;
  wire                load_s1_recoded_sign;
  reg                 load_s1_recoded_special;
  wire                _zz_load_s1_input_ready;
  wire                load_s1_output_valid;
  reg                 load_s1_output_ready;
  wire       [0:0]    load_s1_output_payload_source;
  wire       [4:0]    load_s1_output_payload_rd;
  reg        [52:0]   load_s1_output_payload_value_mantissa;
  reg        [11:0]   load_s1_output_payload_value_exponent;
  reg                 load_s1_output_payload_value_sign;
  reg                 load_s1_output_payload_value_special;
  reg                 load_s1_output_payload_scrap;
  wire       [2:0]    load_s1_output_payload_roundMode;
  wire       [0:0]    load_s1_output_payload_format;
  wire                load_s1_output_payload_NV;
  wire                load_s1_output_payload_DZ;
  wire                when_FpuCore_l594;
  wire                shortPip_input_valid;
  wire                shortPip_input_ready;
  wire       [0:0]    shortPip_input_payload_source;
  wire       [3:0]    shortPip_input_payload_opcode;
  wire       [51:0]   shortPip_input_payload_rs1_mantissa;
  wire       [11:0]   shortPip_input_payload_rs1_exponent;
  wire                shortPip_input_payload_rs1_sign;
  wire                shortPip_input_payload_rs1_special;
  wire       [51:0]   shortPip_input_payload_rs2_mantissa;
  wire       [11:0]   shortPip_input_payload_rs2_exponent;
  wire                shortPip_input_payload_rs2_sign;
  wire                shortPip_input_payload_rs2_special;
  wire       [4:0]    shortPip_input_payload_rd;
  wire       [31:0]   shortPip_input_payload_value;
  wire       [1:0]    shortPip_input_payload_arg;
  wire       [2:0]    shortPip_input_payload_roundMode;
  wire       [0:0]    shortPip_input_payload_format;
  wire                shortPip_input_payload_rs1Boxed;
  wire                shortPip_input_payload_rs2Boxed;
  reg                 decode_shortPip_rValid;
  reg        [0:0]    decode_shortPip_rData_source;
  reg        [3:0]    decode_shortPip_rData_opcode;
  reg        [51:0]   decode_shortPip_rData_rs1_mantissa;
  reg        [11:0]   decode_shortPip_rData_rs1_exponent;
  reg                 decode_shortPip_rData_rs1_sign;
  reg                 decode_shortPip_rData_rs1_special;
  reg        [51:0]   decode_shortPip_rData_rs2_mantissa;
  reg        [11:0]   decode_shortPip_rData_rs2_exponent;
  reg                 decode_shortPip_rData_rs2_sign;
  reg                 decode_shortPip_rData_rs2_special;
  reg        [4:0]    decode_shortPip_rData_rd;
  reg        [31:0]   decode_shortPip_rData_value;
  reg        [1:0]    decode_shortPip_rData_arg;
  reg        [2:0]    decode_shortPip_rData_roundMode;
  reg        [0:0]    decode_shortPip_rData_format;
  reg                 decode_shortPip_rData_rs1Boxed;
  reg                 decode_shortPip_rData_rs2Boxed;
  wire                when_Stream_l375_6;
  wire                shortPip_toFpuRf;
  wire                shortPip_rfOutput_valid;
  wire                shortPip_rfOutput_ready;
  wire       [0:0]    shortPip_rfOutput_payload_source;
  wire       [4:0]    shortPip_rfOutput_payload_rd;
  reg        [52:0]   shortPip_rfOutput_payload_value_mantissa;
  reg        [11:0]   shortPip_rfOutput_payload_value_exponent;
  reg                 shortPip_rfOutput_payload_value_sign;
  reg                 shortPip_rfOutput_payload_value_special;
  wire                shortPip_rfOutput_payload_scrap;
  wire       [2:0]    shortPip_rfOutput_payload_roundMode;
  reg        [0:0]    shortPip_rfOutput_payload_format;
  wire                shortPip_rfOutput_payload_NV;
  wire                shortPip_rfOutput_payload_DZ;
  wire                shortPip_input_fire;
  wire                _zz_when_FpuCore_l221;
  wire                when_FpuCore_l221;
  wire                when_FpuCore_l221_1;
  wire                shortPip_isCommited;
  wire                _zz_shortPip_rfOutput_ready;
  wire                shortPip_output_valid;
  reg                 shortPip_output_ready;
  wire       [0:0]    shortPip_output_payload_source;
  wire       [4:0]    shortPip_output_payload_rd;
  wire       [52:0]   shortPip_output_payload_value_mantissa;
  wire       [11:0]   shortPip_output_payload_value_exponent;
  wire                shortPip_output_payload_value_sign;
  wire                shortPip_output_payload_value_special;
  wire                shortPip_output_payload_scrap;
  wire       [2:0]    shortPip_output_payload_roundMode;
  wire       [0:0]    shortPip_output_payload_format;
  wire                shortPip_output_payload_NV;
  wire                shortPip_output_payload_DZ;
  reg        [63:0]   shortPip_result;
  reg                 shortPip_halt;
  reg        [63:0]   shortPip_recodedResult;
  wire       [7:0]    shortPip_f32_exp;
  wire       [22:0]   shortPip_f32_man;
  wire       [10:0]   shortPip_f64_exp;
  wire       [51:0]   shortPip_f64_man;
  wire                when_FpuCore_l31_1;
  wire       [10:0]   shortPip_expSubnormalThreshold;
  wire                shortPip_expInSubnormalRange;
  wire                shortPip_isSubnormal;
  wire                shortPip_isNormal;
  wire       [11:0]   shortPip_fsm_f2iShift;
  wire                shortPip_fsm_isF2i;
  wire                shortPip_fsm_needRecoding;
  reg                 shortPip_fsm_done;
  reg                 shortPip_fsm_boot;
  wire                shortPip_fsm_isZero;
  reg        [5:0]    shortPip_fsm_shift_by;
  reg        [52:0]   shortPip_fsm_shift_input;
  reg                 shortPip_fsm_shift_scrap;
  wire                when_FpuCore_l646;
  wire                when_FpuCore_l646_1;
  wire                when_FpuCore_l646_2;
  wire                when_FpuCore_l646_3;
  wire                when_FpuCore_l646_4;
  wire                when_FpuCore_l646_5;
  wire                when_FpuCore_l652;
  reg        [52:0]   shortPip_fsm_shift_output;
  wire       [10:0]   shortPip_fsm_formatShiftOffset;
  wire                when_FpuCore_l658;
  wire       [11:0]   _zz_shortPip_fsm_shift_by;
  wire       [5:0]    _zz_shortPip_fsm_shift_by_1;
  wire                shortPip_input_isStall;
  wire                when_FpuCore_l672;
  reg                 shortPip_mantissaForced;
  reg                 shortPip_exponentForced;
  reg                 shortPip_mantissaForcedValue;
  reg                 shortPip_exponentForcedValue;
  reg                 shortPip_cononicalForced;
  wire       [1:0]    switch_FpuCore_l686;
  wire                when_FpuCore_l702;
  wire                when_FpuCore_l31_2;
  wire                when_FpuCore_l31_3;
  wire                when_FpuCore_l31_4;
  wire                when_FpuCore_l31_5;
  reg                 shortPip_rspNv;
  reg                 shortPip_rspNx;
  wire       [31:0]   shortPip_f2i_unsigned;
  wire                shortPip_f2i_resign;
  wire       [1:0]    shortPip_f2i_round;
  reg                 shortPip_f2i_increment;
  reg        [31:0]   shortPip_f2i_result;
  reg                 shortPip_f2i_overflow;
  wire                shortPip_f2i_underflow;
  wire                shortPip_f2i_isZero;
  wire                when_FpuCore_l763;
  wire                when_FpuCore_l767;
  wire                shortPip_bothZero;
  reg                 shortPip_rs1Equal;
  reg                 shortPip_rs1AbsSmaller;
  wire                when_FpuCore_l780;
  wire                when_FpuCore_l781;
  wire                when_FpuCore_l782;
  wire                when_FpuCore_l783;
  wire                when_FpuCore_l784;
  wire       [1:0]    switch_Misc_l241;
  reg                 shortPip_rs1Smaller;
  wire                shortPip_minMaxSelectRs2;
  wire                shortPip_minMaxSelectNanQuiet;
  reg        [0:0]    shortPip_cmpResult;
  wire                when_FpuCore_l796;
  wire                shortPip_sgnjRs1Sign;
  reg                 shortPip_sgnjRs2Sign;
  wire                when_FpuCore_l800;
  wire                shortPip_sgnjResult;
  reg        [31:0]   shortPip_fclassResult;
  wire                shortPip_decoded_isNan;
  wire                shortPip_decoded_isNormal;
  wire                shortPip_decoded_isSubnormal;
  wire                shortPip_decoded_isZero;
  wire                shortPip_decoded_isInfinity;
  wire                shortPip_decoded_isQuiet;
  wire                when_FpuCore_l850;
  wire                when_FpuCore_l853;
  wire       [0:0]    _zz_shortPip_rfOutput_payload_format;
  wire                when_FpuCore_l860;
  wire                shortPip_signalQuiet;
  wire                shortPip_rs1Nan;
  wire                shortPip_rs2Nan;
  wire                shortPip_rs1NanNv;
  wire                shortPip_rs2NanNv;
  wire                shortPip_NV;
  wire                shortPip_rspStreams_0_valid;
  reg                 shortPip_rspStreams_0_ready;
  wire       [63:0]   shortPip_rspStreams_0_payload_value;
  wire                shortPip_rspStreams_0_payload_NV;
  wire                shortPip_rspStreams_0_payload_NX;
  wire                shortPip_rspStreams_1_valid;
  reg                 shortPip_rspStreams_1_ready;
  wire       [63:0]   shortPip_rspStreams_1_payload_value;
  wire                shortPip_rspStreams_1_payload_NV;
  wire                shortPip_rspStreams_1_payload_NX;
  wire                shortPip_rspStreams_0_m2sPipe_valid;
  wire                shortPip_rspStreams_0_m2sPipe_ready;
  wire       [63:0]   shortPip_rspStreams_0_m2sPipe_payload_value;
  wire                shortPip_rspStreams_0_m2sPipe_payload_NV;
  wire                shortPip_rspStreams_0_m2sPipe_payload_NX;
  reg                 shortPip_rspStreams_0_rValid;
  reg        [63:0]   shortPip_rspStreams_0_rData_value;
  reg                 shortPip_rspStreams_0_rData_NV;
  reg                 shortPip_rspStreams_0_rData_NX;
  wire                when_Stream_l375_7;
  wire                shortPip_rspStreams_1_m2sPipe_valid;
  wire                shortPip_rspStreams_1_m2sPipe_ready;
  wire       [63:0]   shortPip_rspStreams_1_m2sPipe_payload_value;
  wire                shortPip_rspStreams_1_m2sPipe_payload_NV;
  wire                shortPip_rspStreams_1_m2sPipe_payload_NX;
  reg                 shortPip_rspStreams_1_rValid;
  reg        [63:0]   shortPip_rspStreams_1_rData_value;
  reg                 shortPip_rspStreams_1_rData_NV;
  reg                 shortPip_rspStreams_1_rData_NX;
  wire                when_Stream_l375_8;
  wire                mul_preMul_input_valid;
  wire                mul_preMul_input_ready;
  wire       [0:0]    mul_preMul_input_payload_source;
  wire       [51:0]   mul_preMul_input_payload_rs1_mantissa;
  wire       [11:0]   mul_preMul_input_payload_rs1_exponent;
  wire                mul_preMul_input_payload_rs1_sign;
  wire                mul_preMul_input_payload_rs1_special;
  wire       [51:0]   mul_preMul_input_payload_rs2_mantissa;
  wire       [11:0]   mul_preMul_input_payload_rs2_exponent;
  wire                mul_preMul_input_payload_rs2_sign;
  wire                mul_preMul_input_payload_rs2_special;
  wire       [51:0]   mul_preMul_input_payload_rs3_mantissa;
  wire       [11:0]   mul_preMul_input_payload_rs3_exponent;
  wire                mul_preMul_input_payload_rs3_sign;
  wire                mul_preMul_input_payload_rs3_special;
  wire       [4:0]    mul_preMul_input_payload_rd;
  wire                mul_preMul_input_payload_add;
  wire                mul_preMul_input_payload_divSqrt;
  wire                mul_preMul_input_payload_msb1;
  wire                mul_preMul_input_payload_msb2;
  wire       [2:0]    mul_preMul_input_payload_roundMode;
  wire       [0:0]    mul_preMul_input_payload_format;
  reg                 decode_mul_rValid;
  reg        [0:0]    decode_mul_rData_source;
  reg        [51:0]   decode_mul_rData_rs1_mantissa;
  reg        [11:0]   decode_mul_rData_rs1_exponent;
  reg                 decode_mul_rData_rs1_sign;
  reg                 decode_mul_rData_rs1_special;
  reg        [51:0]   decode_mul_rData_rs2_mantissa;
  reg        [11:0]   decode_mul_rData_rs2_exponent;
  reg                 decode_mul_rData_rs2_sign;
  reg                 decode_mul_rData_rs2_special;
  reg        [51:0]   decode_mul_rData_rs3_mantissa;
  reg        [11:0]   decode_mul_rData_rs3_exponent;
  reg                 decode_mul_rData_rs3_sign;
  reg                 decode_mul_rData_rs3_special;
  reg        [4:0]    decode_mul_rData_rd;
  reg                 decode_mul_rData_add;
  reg                 decode_mul_rData_divSqrt;
  reg                 decode_mul_rData_msb1;
  reg                 decode_mul_rData_msb2;
  reg        [2:0]    decode_mul_rData_roundMode;
  reg        [0:0]    decode_mul_rData_format;
  wire                when_Stream_l375_9;
  wire                mul_preMul_output_valid;
  reg                 mul_preMul_output_ready;
  wire       [0:0]    mul_preMul_output_payload_source;
  wire       [51:0]   mul_preMul_output_payload_rs1_mantissa;
  wire       [11:0]   mul_preMul_output_payload_rs1_exponent;
  wire                mul_preMul_output_payload_rs1_sign;
  wire                mul_preMul_output_payload_rs1_special;
  wire       [51:0]   mul_preMul_output_payload_rs2_mantissa;
  wire       [11:0]   mul_preMul_output_payload_rs2_exponent;
  wire                mul_preMul_output_payload_rs2_sign;
  wire                mul_preMul_output_payload_rs2_special;
  wire       [51:0]   mul_preMul_output_payload_rs3_mantissa;
  wire       [11:0]   mul_preMul_output_payload_rs3_exponent;
  wire                mul_preMul_output_payload_rs3_sign;
  wire                mul_preMul_output_payload_rs3_special;
  wire       [4:0]    mul_preMul_output_payload_rd;
  wire                mul_preMul_output_payload_add;
  wire                mul_preMul_output_payload_divSqrt;
  wire                mul_preMul_output_payload_msb1;
  wire                mul_preMul_output_payload_msb2;
  wire       [2:0]    mul_preMul_output_payload_roundMode;
  wire       [0:0]    mul_preMul_output_payload_format;
  wire       [12:0]   mul_preMul_output_payload_exp;
  wire                mul_mul_input_valid;
  wire                mul_mul_input_ready;
  wire       [0:0]    mul_mul_input_payload_source;
  wire       [51:0]   mul_mul_input_payload_rs1_mantissa;
  wire       [11:0]   mul_mul_input_payload_rs1_exponent;
  wire                mul_mul_input_payload_rs1_sign;
  wire                mul_mul_input_payload_rs1_special;
  wire       [51:0]   mul_mul_input_payload_rs2_mantissa;
  wire       [11:0]   mul_mul_input_payload_rs2_exponent;
  wire                mul_mul_input_payload_rs2_sign;
  wire                mul_mul_input_payload_rs2_special;
  wire       [51:0]   mul_mul_input_payload_rs3_mantissa;
  wire       [11:0]   mul_mul_input_payload_rs3_exponent;
  wire                mul_mul_input_payload_rs3_sign;
  wire                mul_mul_input_payload_rs3_special;
  wire       [4:0]    mul_mul_input_payload_rd;
  wire                mul_mul_input_payload_add;
  wire                mul_mul_input_payload_divSqrt;
  wire                mul_mul_input_payload_msb1;
  wire                mul_mul_input_payload_msb2;
  wire       [2:0]    mul_mul_input_payload_roundMode;
  wire       [0:0]    mul_mul_input_payload_format;
  wire       [12:0]   mul_mul_input_payload_exp;
  reg                 mul_preMul_output_rValid;
  reg        [0:0]    mul_preMul_output_rData_source;
  reg        [51:0]   mul_preMul_output_rData_rs1_mantissa;
  reg        [11:0]   mul_preMul_output_rData_rs1_exponent;
  reg                 mul_preMul_output_rData_rs1_sign;
  reg                 mul_preMul_output_rData_rs1_special;
  reg        [51:0]   mul_preMul_output_rData_rs2_mantissa;
  reg        [11:0]   mul_preMul_output_rData_rs2_exponent;
  reg                 mul_preMul_output_rData_rs2_sign;
  reg                 mul_preMul_output_rData_rs2_special;
  reg        [51:0]   mul_preMul_output_rData_rs3_mantissa;
  reg        [11:0]   mul_preMul_output_rData_rs3_exponent;
  reg                 mul_preMul_output_rData_rs3_sign;
  reg                 mul_preMul_output_rData_rs3_special;
  reg        [4:0]    mul_preMul_output_rData_rd;
  reg                 mul_preMul_output_rData_add;
  reg                 mul_preMul_output_rData_divSqrt;
  reg                 mul_preMul_output_rData_msb1;
  reg                 mul_preMul_output_rData_msb2;
  reg        [2:0]    mul_preMul_output_rData_roundMode;
  reg        [0:0]    mul_preMul_output_rData_format;
  reg        [12:0]   mul_preMul_output_rData_exp;
  wire                when_Stream_l375_10;
  wire                mul_mul_output_valid;
  reg                 mul_mul_output_ready;
  wire       [0:0]    mul_mul_output_payload_source;
  wire       [51:0]   mul_mul_output_payload_rs1_mantissa;
  wire       [11:0]   mul_mul_output_payload_rs1_exponent;
  wire                mul_mul_output_payload_rs1_sign;
  wire                mul_mul_output_payload_rs1_special;
  wire       [51:0]   mul_mul_output_payload_rs2_mantissa;
  wire       [11:0]   mul_mul_output_payload_rs2_exponent;
  wire                mul_mul_output_payload_rs2_sign;
  wire                mul_mul_output_payload_rs2_special;
  wire       [51:0]   mul_mul_output_payload_rs3_mantissa;
  wire       [11:0]   mul_mul_output_payload_rs3_exponent;
  wire                mul_mul_output_payload_rs3_sign;
  wire                mul_mul_output_payload_rs3_special;
  wire       [4:0]    mul_mul_output_payload_rd;
  wire                mul_mul_output_payload_add;
  wire                mul_mul_output_payload_divSqrt;
  wire                mul_mul_output_payload_msb1;
  wire                mul_mul_output_payload_msb2;
  wire       [2:0]    mul_mul_output_payload_roundMode;
  wire       [0:0]    mul_mul_output_payload_format;
  wire       [12:0]   mul_mul_output_payload_exp;
  wire       [35:0]   mul_mul_output_payload_muls_0;
  wire       [35:0]   mul_mul_output_payload_muls_1;
  wire       [35:0]   mul_mul_output_payload_muls_2;
  wire       [34:0]   mul_mul_output_payload_muls_3;
  wire       [34:0]   mul_mul_output_payload_muls_4;
  wire       [35:0]   mul_mul_output_payload_muls_5;
  wire       [34:0]   mul_mul_output_payload_muls_6;
  wire       [34:0]   mul_mul_output_payload_muls_7;
  wire       [33:0]   mul_mul_output_payload_muls_8;
  wire       [52:0]   mul_mul_mulA;
  wire       [52:0]   mul_mul_mulB;
  wire                mul_sum1_input_valid;
  wire                mul_sum1_input_ready;
  wire       [0:0]    mul_sum1_input_payload_source;
  wire       [51:0]   mul_sum1_input_payload_rs1_mantissa;
  wire       [11:0]   mul_sum1_input_payload_rs1_exponent;
  wire                mul_sum1_input_payload_rs1_sign;
  wire                mul_sum1_input_payload_rs1_special;
  wire       [51:0]   mul_sum1_input_payload_rs2_mantissa;
  wire       [11:0]   mul_sum1_input_payload_rs2_exponent;
  wire                mul_sum1_input_payload_rs2_sign;
  wire                mul_sum1_input_payload_rs2_special;
  wire       [51:0]   mul_sum1_input_payload_rs3_mantissa;
  wire       [11:0]   mul_sum1_input_payload_rs3_exponent;
  wire                mul_sum1_input_payload_rs3_sign;
  wire                mul_sum1_input_payload_rs3_special;
  wire       [4:0]    mul_sum1_input_payload_rd;
  wire                mul_sum1_input_payload_add;
  wire                mul_sum1_input_payload_divSqrt;
  wire                mul_sum1_input_payload_msb1;
  wire                mul_sum1_input_payload_msb2;
  wire       [2:0]    mul_sum1_input_payload_roundMode;
  wire       [0:0]    mul_sum1_input_payload_format;
  wire       [12:0]   mul_sum1_input_payload_exp;
  wire       [35:0]   mul_sum1_input_payload_muls_0;
  wire       [35:0]   mul_sum1_input_payload_muls_1;
  wire       [35:0]   mul_sum1_input_payload_muls_2;
  wire       [34:0]   mul_sum1_input_payload_muls_3;
  wire       [34:0]   mul_sum1_input_payload_muls_4;
  wire       [35:0]   mul_sum1_input_payload_muls_5;
  wire       [34:0]   mul_sum1_input_payload_muls_6;
  wire       [34:0]   mul_sum1_input_payload_muls_7;
  wire       [33:0]   mul_sum1_input_payload_muls_8;
  reg                 mul_mul_output_rValid;
  reg        [0:0]    mul_mul_output_rData_source;
  reg        [51:0]   mul_mul_output_rData_rs1_mantissa;
  reg        [11:0]   mul_mul_output_rData_rs1_exponent;
  reg                 mul_mul_output_rData_rs1_sign;
  reg                 mul_mul_output_rData_rs1_special;
  reg        [51:0]   mul_mul_output_rData_rs2_mantissa;
  reg        [11:0]   mul_mul_output_rData_rs2_exponent;
  reg                 mul_mul_output_rData_rs2_sign;
  reg                 mul_mul_output_rData_rs2_special;
  reg        [51:0]   mul_mul_output_rData_rs3_mantissa;
  reg        [11:0]   mul_mul_output_rData_rs3_exponent;
  reg                 mul_mul_output_rData_rs3_sign;
  reg                 mul_mul_output_rData_rs3_special;
  reg        [4:0]    mul_mul_output_rData_rd;
  reg                 mul_mul_output_rData_add;
  reg                 mul_mul_output_rData_divSqrt;
  reg                 mul_mul_output_rData_msb1;
  reg                 mul_mul_output_rData_msb2;
  reg        [2:0]    mul_mul_output_rData_roundMode;
  reg        [0:0]    mul_mul_output_rData_format;
  reg        [12:0]   mul_mul_output_rData_exp;
  reg        [35:0]   mul_mul_output_rData_muls_0;
  reg        [35:0]   mul_mul_output_rData_muls_1;
  reg        [35:0]   mul_mul_output_rData_muls_2;
  reg        [34:0]   mul_mul_output_rData_muls_3;
  reg        [34:0]   mul_mul_output_rData_muls_4;
  reg        [35:0]   mul_mul_output_rData_muls_5;
  reg        [34:0]   mul_mul_output_rData_muls_6;
  reg        [34:0]   mul_mul_output_rData_muls_7;
  reg        [33:0]   mul_mul_output_rData_muls_8;
  wire                when_Stream_l375_11;
  wire       [105:0]  mul_sum1_sum;
  wire                mul_sum1_output_valid;
  reg                 mul_sum1_output_ready;
  wire       [0:0]    mul_sum1_output_payload_source;
  wire       [51:0]   mul_sum1_output_payload_rs1_mantissa;
  wire       [11:0]   mul_sum1_output_payload_rs1_exponent;
  wire                mul_sum1_output_payload_rs1_sign;
  wire                mul_sum1_output_payload_rs1_special;
  wire       [51:0]   mul_sum1_output_payload_rs2_mantissa;
  wire       [11:0]   mul_sum1_output_payload_rs2_exponent;
  wire                mul_sum1_output_payload_rs2_sign;
  wire                mul_sum1_output_payload_rs2_special;
  wire       [51:0]   mul_sum1_output_payload_rs3_mantissa;
  wire       [11:0]   mul_sum1_output_payload_rs3_exponent;
  wire                mul_sum1_output_payload_rs3_sign;
  wire                mul_sum1_output_payload_rs3_special;
  wire       [4:0]    mul_sum1_output_payload_rd;
  wire                mul_sum1_output_payload_add;
  wire                mul_sum1_output_payload_divSqrt;
  wire                mul_sum1_output_payload_msb1;
  wire                mul_sum1_output_payload_msb2;
  wire       [2:0]    mul_sum1_output_payload_roundMode;
  wire       [0:0]    mul_sum1_output_payload_format;
  wire       [12:0]   mul_sum1_output_payload_exp;
  wire       [34:0]   mul_sum1_output_payload_muls2_0;
  wire       [35:0]   mul_sum1_output_payload_muls2_1;
  wire       [34:0]   mul_sum1_output_payload_muls2_2;
  wire       [34:0]   mul_sum1_output_payload_muls2_3;
  wire       [33:0]   mul_sum1_output_payload_muls2_4;
  wire       [105:0]  mul_sum1_output_payload_mulC2;
  wire                mul_sum2_input_valid;
  wire                mul_sum2_input_ready;
  wire       [0:0]    mul_sum2_input_payload_source;
  wire       [51:0]   mul_sum2_input_payload_rs1_mantissa;
  wire       [11:0]   mul_sum2_input_payload_rs1_exponent;
  wire                mul_sum2_input_payload_rs1_sign;
  wire                mul_sum2_input_payload_rs1_special;
  wire       [51:0]   mul_sum2_input_payload_rs2_mantissa;
  wire       [11:0]   mul_sum2_input_payload_rs2_exponent;
  wire                mul_sum2_input_payload_rs2_sign;
  wire                mul_sum2_input_payload_rs2_special;
  wire       [51:0]   mul_sum2_input_payload_rs3_mantissa;
  wire       [11:0]   mul_sum2_input_payload_rs3_exponent;
  wire                mul_sum2_input_payload_rs3_sign;
  wire                mul_sum2_input_payload_rs3_special;
  wire       [4:0]    mul_sum2_input_payload_rd;
  wire                mul_sum2_input_payload_add;
  wire                mul_sum2_input_payload_divSqrt;
  wire                mul_sum2_input_payload_msb1;
  wire                mul_sum2_input_payload_msb2;
  wire       [2:0]    mul_sum2_input_payload_roundMode;
  wire       [0:0]    mul_sum2_input_payload_format;
  wire       [12:0]   mul_sum2_input_payload_exp;
  wire       [34:0]   mul_sum2_input_payload_muls2_0;
  wire       [35:0]   mul_sum2_input_payload_muls2_1;
  wire       [34:0]   mul_sum2_input_payload_muls2_2;
  wire       [34:0]   mul_sum2_input_payload_muls2_3;
  wire       [33:0]   mul_sum2_input_payload_muls2_4;
  wire       [105:0]  mul_sum2_input_payload_mulC2;
  reg                 mul_sum1_output_rValid;
  reg        [0:0]    mul_sum1_output_rData_source;
  reg        [51:0]   mul_sum1_output_rData_rs1_mantissa;
  reg        [11:0]   mul_sum1_output_rData_rs1_exponent;
  reg                 mul_sum1_output_rData_rs1_sign;
  reg                 mul_sum1_output_rData_rs1_special;
  reg        [51:0]   mul_sum1_output_rData_rs2_mantissa;
  reg        [11:0]   mul_sum1_output_rData_rs2_exponent;
  reg                 mul_sum1_output_rData_rs2_sign;
  reg                 mul_sum1_output_rData_rs2_special;
  reg        [51:0]   mul_sum1_output_rData_rs3_mantissa;
  reg        [11:0]   mul_sum1_output_rData_rs3_exponent;
  reg                 mul_sum1_output_rData_rs3_sign;
  reg                 mul_sum1_output_rData_rs3_special;
  reg        [4:0]    mul_sum1_output_rData_rd;
  reg                 mul_sum1_output_rData_add;
  reg                 mul_sum1_output_rData_divSqrt;
  reg                 mul_sum1_output_rData_msb1;
  reg                 mul_sum1_output_rData_msb2;
  reg        [2:0]    mul_sum1_output_rData_roundMode;
  reg        [0:0]    mul_sum1_output_rData_format;
  reg        [12:0]   mul_sum1_output_rData_exp;
  reg        [34:0]   mul_sum1_output_rData_muls2_0;
  reg        [35:0]   mul_sum1_output_rData_muls2_1;
  reg        [34:0]   mul_sum1_output_rData_muls2_2;
  reg        [34:0]   mul_sum1_output_rData_muls2_3;
  reg        [33:0]   mul_sum1_output_rData_muls2_4;
  reg        [105:0]  mul_sum1_output_rData_mulC2;
  wire                when_Stream_l375_12;
  wire       [105:0]  mul_sum2_sum;
  wire                mul_sum2_input_fire;
  wire                when_FpuCore_l221_2;
  wire                when_FpuCore_l221_3;
  wire                mul_sum2_isCommited;
  wire                _zz_mul_sum2_input_ready;
  wire                mul_sum2_output_valid;
  reg                 mul_sum2_output_ready;
  wire       [0:0]    mul_sum2_output_payload_source;
  wire       [51:0]   mul_sum2_output_payload_rs1_mantissa;
  wire       [11:0]   mul_sum2_output_payload_rs1_exponent;
  wire                mul_sum2_output_payload_rs1_sign;
  wire                mul_sum2_output_payload_rs1_special;
  wire       [51:0]   mul_sum2_output_payload_rs2_mantissa;
  wire       [11:0]   mul_sum2_output_payload_rs2_exponent;
  wire                mul_sum2_output_payload_rs2_sign;
  wire                mul_sum2_output_payload_rs2_special;
  wire       [51:0]   mul_sum2_output_payload_rs3_mantissa;
  wire       [11:0]   mul_sum2_output_payload_rs3_exponent;
  wire                mul_sum2_output_payload_rs3_sign;
  wire                mul_sum2_output_payload_rs3_special;
  wire       [4:0]    mul_sum2_output_payload_rd;
  wire                mul_sum2_output_payload_add;
  wire                mul_sum2_output_payload_divSqrt;
  wire                mul_sum2_output_payload_msb1;
  wire                mul_sum2_output_payload_msb2;
  wire       [2:0]    mul_sum2_output_payload_roundMode;
  wire       [0:0]    mul_sum2_output_payload_format;
  wire       [12:0]   mul_sum2_output_payload_exp;
  wire       [105:0]  mul_sum2_output_payload_mulC;
  wire                mul_norm_input_valid;
  wire                mul_norm_input_ready;
  wire       [0:0]    mul_norm_input_payload_source;
  wire       [51:0]   mul_norm_input_payload_rs1_mantissa;
  wire       [11:0]   mul_norm_input_payload_rs1_exponent;
  wire                mul_norm_input_payload_rs1_sign;
  wire                mul_norm_input_payload_rs1_special;
  wire       [51:0]   mul_norm_input_payload_rs2_mantissa;
  wire       [11:0]   mul_norm_input_payload_rs2_exponent;
  wire                mul_norm_input_payload_rs2_sign;
  wire                mul_norm_input_payload_rs2_special;
  wire       [51:0]   mul_norm_input_payload_rs3_mantissa;
  wire       [11:0]   mul_norm_input_payload_rs3_exponent;
  wire                mul_norm_input_payload_rs3_sign;
  wire                mul_norm_input_payload_rs3_special;
  wire       [4:0]    mul_norm_input_payload_rd;
  wire                mul_norm_input_payload_add;
  wire                mul_norm_input_payload_divSqrt;
  wire                mul_norm_input_payload_msb1;
  wire                mul_norm_input_payload_msb2;
  wire       [2:0]    mul_norm_input_payload_roundMode;
  wire       [0:0]    mul_norm_input_payload_format;
  wire       [12:0]   mul_norm_input_payload_exp;
  wire       [105:0]  mul_norm_input_payload_mulC;
  reg                 mul_sum2_output_rValid;
  reg        [0:0]    mul_sum2_output_rData_source;
  reg        [51:0]   mul_sum2_output_rData_rs1_mantissa;
  reg        [11:0]   mul_sum2_output_rData_rs1_exponent;
  reg                 mul_sum2_output_rData_rs1_sign;
  reg                 mul_sum2_output_rData_rs1_special;
  reg        [51:0]   mul_sum2_output_rData_rs2_mantissa;
  reg        [11:0]   mul_sum2_output_rData_rs2_exponent;
  reg                 mul_sum2_output_rData_rs2_sign;
  reg                 mul_sum2_output_rData_rs2_special;
  reg        [51:0]   mul_sum2_output_rData_rs3_mantissa;
  reg        [11:0]   mul_sum2_output_rData_rs3_exponent;
  reg                 mul_sum2_output_rData_rs3_sign;
  reg                 mul_sum2_output_rData_rs3_special;
  reg        [4:0]    mul_sum2_output_rData_rd;
  reg                 mul_sum2_output_rData_add;
  reg                 mul_sum2_output_rData_divSqrt;
  reg                 mul_sum2_output_rData_msb1;
  reg                 mul_sum2_output_rData_msb2;
  reg        [2:0]    mul_sum2_output_rData_roundMode;
  reg        [0:0]    mul_sum2_output_rData_format;
  reg        [12:0]   mul_sum2_output_rData_exp;
  reg        [105:0]  mul_sum2_output_rData_mulC;
  wire                when_Stream_l375_13;
  wire       [54:0]   mul_norm_mulHigh;
  wire       [50:0]   mul_norm_mulLow;
  reg                 mul_norm_scrap;
  wire                mul_norm_needShift;
  wire       [12:0]   mul_norm_exp;
  wire       [52:0]   mul_norm_man;
  wire                when_FpuCore_l967;
  wire                mul_norm_forceZero;
  wire       [11:0]   mul_norm_underflowThreshold;
  wire       [10:0]   mul_norm_underflowExp;
  wire                mul_norm_forceUnderflow;
  wire                mul_norm_forceOverflow;
  wire                mul_norm_infinitynan;
  wire                mul_norm_forceNan;
  reg        [52:0]   mul_norm_output_mantissa;
  reg        [11:0]   mul_norm_output_exponent;
  wire                mul_norm_output_sign;
  reg                 mul_norm_output_special;
  reg                 mul_norm_NV;
  wire                when_FpuCore_l983;
  wire                when_FpuCore_l987;
  wire                mul_result_notMul_output_valid;
  wire       [52:0]   mul_result_notMul_output_payload;
  wire                mul_result_output_valid;
  wire                mul_result_output_ready;
  wire       [0:0]    mul_result_output_payload_source;
  wire       [4:0]    mul_result_output_payload_rd;
  wire       [52:0]   mul_result_output_payload_value_mantissa;
  wire       [11:0]   mul_result_output_payload_value_exponent;
  wire                mul_result_output_payload_value_sign;
  wire                mul_result_output_payload_value_special;
  wire                mul_result_output_payload_scrap;
  wire       [2:0]    mul_result_output_payload_roundMode;
  wire       [0:0]    mul_result_output_payload_format;
  wire                mul_result_output_payload_NV;
  wire                mul_result_output_payload_DZ;
  wire                mul_result_mulToAdd_valid;
  reg                 mul_result_mulToAdd_ready;
  wire       [0:0]    mul_result_mulToAdd_payload_source;
  reg        [53:0]   mul_result_mulToAdd_payload_rs1_mantissa;
  wire       [11:0]   mul_result_mulToAdd_payload_rs1_exponent;
  wire                mul_result_mulToAdd_payload_rs1_sign;
  wire                mul_result_mulToAdd_payload_rs1_special;
  wire       [53:0]   mul_result_mulToAdd_payload_rs2_mantissa;
  wire       [11:0]   mul_result_mulToAdd_payload_rs2_exponent;
  wire                mul_result_mulToAdd_payload_rs2_sign;
  wire                mul_result_mulToAdd_payload_rs2_special;
  wire       [4:0]    mul_result_mulToAdd_payload_rd;
  wire       [2:0]    mul_result_mulToAdd_payload_roundMode;
  wire       [0:0]    mul_result_mulToAdd_payload_format;
  wire                mul_result_mulToAdd_payload_needCommit;
  wire                mul_result_mulToAdd_m2sPipe_valid;
  wire                mul_result_mulToAdd_m2sPipe_ready;
  wire       [0:0]    mul_result_mulToAdd_m2sPipe_payload_source;
  wire       [53:0]   mul_result_mulToAdd_m2sPipe_payload_rs1_mantissa;
  wire       [11:0]   mul_result_mulToAdd_m2sPipe_payload_rs1_exponent;
  wire                mul_result_mulToAdd_m2sPipe_payload_rs1_sign;
  wire                mul_result_mulToAdd_m2sPipe_payload_rs1_special;
  wire       [53:0]   mul_result_mulToAdd_m2sPipe_payload_rs2_mantissa;
  wire       [11:0]   mul_result_mulToAdd_m2sPipe_payload_rs2_exponent;
  wire                mul_result_mulToAdd_m2sPipe_payload_rs2_sign;
  wire                mul_result_mulToAdd_m2sPipe_payload_rs2_special;
  wire       [4:0]    mul_result_mulToAdd_m2sPipe_payload_rd;
  wire       [2:0]    mul_result_mulToAdd_m2sPipe_payload_roundMode;
  wire       [0:0]    mul_result_mulToAdd_m2sPipe_payload_format;
  wire                mul_result_mulToAdd_m2sPipe_payload_needCommit;
  reg                 mul_result_mulToAdd_rValid;
  reg        [0:0]    mul_result_mulToAdd_rData_source;
  reg        [53:0]   mul_result_mulToAdd_rData_rs1_mantissa;
  reg        [11:0]   mul_result_mulToAdd_rData_rs1_exponent;
  reg                 mul_result_mulToAdd_rData_rs1_sign;
  reg                 mul_result_mulToAdd_rData_rs1_special;
  reg        [53:0]   mul_result_mulToAdd_rData_rs2_mantissa;
  reg        [11:0]   mul_result_mulToAdd_rData_rs2_exponent;
  reg                 mul_result_mulToAdd_rData_rs2_sign;
  reg                 mul_result_mulToAdd_rData_rs2_special;
  reg        [4:0]    mul_result_mulToAdd_rData_rd;
  reg        [2:0]    mul_result_mulToAdd_rData_roundMode;
  reg        [0:0]    mul_result_mulToAdd_rData_format;
  reg                 mul_result_mulToAdd_rData_needCommit;
  wire                when_Stream_l375_14;
  wire                div_input_valid;
  wire                div_input_ready;
  wire       [0:0]    div_input_payload_source;
  wire       [51:0]   div_input_payload_rs1_mantissa;
  wire       [11:0]   div_input_payload_rs1_exponent;
  wire                div_input_payload_rs1_sign;
  wire                div_input_payload_rs1_special;
  wire       [51:0]   div_input_payload_rs2_mantissa;
  wire       [11:0]   div_input_payload_rs2_exponent;
  wire                div_input_payload_rs2_sign;
  wire                div_input_payload_rs2_special;
  wire       [4:0]    div_input_payload_rd;
  wire       [2:0]    div_input_payload_roundMode;
  wire       [0:0]    div_input_payload_format;
  reg                 decode_div_rValid;
  wire                div_input_fire;
  reg        [0:0]    decode_div_rData_source;
  reg        [51:0]   decode_div_rData_rs1_mantissa;
  reg        [11:0]   decode_div_rData_rs1_exponent;
  reg                 decode_div_rData_rs1_sign;
  reg                 decode_div_rData_rs1_special;
  reg        [51:0]   decode_div_rData_rs2_mantissa;
  reg        [11:0]   decode_div_rData_rs2_exponent;
  reg                 decode_div_rData_rs2_sign;
  reg                 decode_div_rData_rs2_special;
  reg        [4:0]    decode_div_rData_rd;
  reg        [2:0]    decode_div_rData_roundMode;
  reg        [0:0]    decode_div_rData_format;
  reg                 div_haltIt;
  wire                when_FpuCore_l221_4;
  wire                when_FpuCore_l221_5;
  reg                 div_isCommited;
  wire                _zz_div_input_ready;
  wire                div_output_valid;
  wire                div_output_ready;
  wire       [0:0]    div_output_payload_source;
  wire       [4:0]    div_output_payload_rd;
  reg        [52:0]   div_output_payload_value_mantissa;
  reg        [11:0]   div_output_payload_value_exponent;
  wire                div_output_payload_value_sign;
  reg                 div_output_payload_value_special;
  wire                div_output_payload_scrap;
  wire       [2:0]    div_output_payload_roundMode;
  wire       [0:0]    div_output_payload_format;
  reg                 div_output_payload_NV;
  wire                div_output_payload_DZ;
  wire       [54:0]   div_dividerResult;
  wire                div_dividerScrap;
  reg                 div_cmdSent;
  wire                div_divider_io_input_fire;
  wire                when_FpuCore_l1056;
  wire                div_needShift;
  wire       [52:0]   div_mantissa;
  wire                div_scrap;
  wire       [13:0]   div_exponent;
  wire                when_FpuCore_l1072;
  wire       [13:0]   div_underflowThreshold;
  wire       [13:0]   div_underflowExp;
  wire                div_forceUnderflow;
  wire                div_forceOverflow;
  wire                div_infinitynan;
  wire                div_forceNan;
  wire                div_forceZero;
  wire                when_FpuCore_l1089;
  wire                when_FpuCore_l1093;
  wire                sqrt_input_valid;
  wire                sqrt_input_ready;
  wire       [0:0]    sqrt_input_payload_source;
  wire       [51:0]   sqrt_input_payload_rs1_mantissa;
  wire       [11:0]   sqrt_input_payload_rs1_exponent;
  wire                sqrt_input_payload_rs1_sign;
  wire                sqrt_input_payload_rs1_special;
  wire       [4:0]    sqrt_input_payload_rd;
  wire       [2:0]    sqrt_input_payload_roundMode;
  wire       [0:0]    sqrt_input_payload_format;
  reg                 decode_sqrt_rValid;
  wire                sqrt_input_fire;
  reg        [0:0]    decode_sqrt_rData_source;
  reg        [51:0]   decode_sqrt_rData_rs1_mantissa;
  reg        [11:0]   decode_sqrt_rData_rs1_exponent;
  reg                 decode_sqrt_rData_rs1_sign;
  reg                 decode_sqrt_rData_rs1_special;
  reg        [4:0]    decode_sqrt_rData_rd;
  reg        [2:0]    decode_sqrt_rData_roundMode;
  reg        [0:0]    decode_sqrt_rData_format;
  reg                 sqrt_haltIt;
  wire                when_FpuCore_l221_6;
  wire                when_FpuCore_l221_7;
  reg                 sqrt_isCommited;
  wire                _zz_sqrt_input_ready;
  wire                sqrt_output_valid;
  wire                sqrt_output_ready;
  wire       [0:0]    sqrt_output_payload_source;
  wire       [4:0]    sqrt_output_payload_rd;
  reg        [52:0]   sqrt_output_payload_value_mantissa;
  reg        [11:0]   sqrt_output_payload_value_exponent;
  wire                sqrt_output_payload_value_sign;
  reg                 sqrt_output_payload_value_special;
  wire                sqrt_output_payload_scrap;
  wire       [2:0]    sqrt_output_payload_roundMode;
  wire       [0:0]    sqrt_output_payload_format;
  reg                 sqrt_output_payload_NV;
  wire                sqrt_output_payload_DZ;
  wire                sqrt_needShift;
  reg                 sqrt_cmdSent;
  wire                sqrt_sqrt_io_input_fire;
  wire                when_FpuCore_l1118;
  wire                sqrt_scrap;
  reg        [11:0]   sqrt_exponent;
  wire                sqrt_negative;
  wire                when_FpuCore_l1137;
  wire                when_FpuCore_l1144;
  wire                when_FpuCore_l1148;
  wire                add_preShifter_input_valid;
  wire                add_preShifter_input_ready;
  wire       [0:0]    add_preShifter_input_payload_source;
  wire       [53:0]   add_preShifter_input_payload_rs1_mantissa;
  wire       [11:0]   add_preShifter_input_payload_rs1_exponent;
  wire                add_preShifter_input_payload_rs1_sign;
  wire                add_preShifter_input_payload_rs1_special;
  wire       [53:0]   add_preShifter_input_payload_rs2_mantissa;
  wire       [11:0]   add_preShifter_input_payload_rs2_exponent;
  wire                add_preShifter_input_payload_rs2_sign;
  wire                add_preShifter_input_payload_rs2_special;
  wire       [4:0]    add_preShifter_input_payload_rd;
  wire       [2:0]    add_preShifter_input_payload_roundMode;
  wire       [0:0]    add_preShifter_input_payload_format;
  wire                add_preShifter_input_payload_needCommit;
  wire                add_preShifter_output_valid;
  reg                 add_preShifter_output_ready;
  wire       [0:0]    add_preShifter_output_payload_source;
  wire       [53:0]   add_preShifter_output_payload_rs1_mantissa;
  wire       [11:0]   add_preShifter_output_payload_rs1_exponent;
  wire                add_preShifter_output_payload_rs1_sign;
  wire                add_preShifter_output_payload_rs1_special;
  wire       [53:0]   add_preShifter_output_payload_rs2_mantissa;
  wire       [11:0]   add_preShifter_output_payload_rs2_exponent;
  wire                add_preShifter_output_payload_rs2_sign;
  wire                add_preShifter_output_payload_rs2_special;
  wire       [4:0]    add_preShifter_output_payload_rd;
  wire       [2:0]    add_preShifter_output_payload_roundMode;
  wire       [0:0]    add_preShifter_output_payload_format;
  wire                add_preShifter_output_payload_needCommit;
  wire                add_preShifter_output_payload_absRs1Bigger;
  wire                add_preShifter_output_payload_rs1ExponentBigger;
  wire       [12:0]   add_preShifter_exp21;
  wire                add_preShifter_rs1ExponentBigger;
  wire                add_preShifter_rs1ExponentEqual;
  wire                add_preShifter_rs1MantissaBigger;
  wire                add_preShifter_absRs1Bigger;
  wire                add_shifter_input_valid;
  wire                add_shifter_input_ready;
  wire       [0:0]    add_shifter_input_payload_source;
  wire       [53:0]   add_shifter_input_payload_rs1_mantissa;
  wire       [11:0]   add_shifter_input_payload_rs1_exponent;
  wire                add_shifter_input_payload_rs1_sign;
  wire                add_shifter_input_payload_rs1_special;
  wire       [53:0]   add_shifter_input_payload_rs2_mantissa;
  wire       [11:0]   add_shifter_input_payload_rs2_exponent;
  wire                add_shifter_input_payload_rs2_sign;
  wire                add_shifter_input_payload_rs2_special;
  wire       [4:0]    add_shifter_input_payload_rd;
  wire       [2:0]    add_shifter_input_payload_roundMode;
  wire       [0:0]    add_shifter_input_payload_format;
  wire                add_shifter_input_payload_needCommit;
  wire                add_shifter_input_payload_absRs1Bigger;
  wire                add_shifter_input_payload_rs1ExponentBigger;
  reg                 add_preShifter_output_rValid;
  reg        [0:0]    add_preShifter_output_rData_source;
  reg        [53:0]   add_preShifter_output_rData_rs1_mantissa;
  reg        [11:0]   add_preShifter_output_rData_rs1_exponent;
  reg                 add_preShifter_output_rData_rs1_sign;
  reg                 add_preShifter_output_rData_rs1_special;
  reg        [53:0]   add_preShifter_output_rData_rs2_mantissa;
  reg        [11:0]   add_preShifter_output_rData_rs2_exponent;
  reg                 add_preShifter_output_rData_rs2_sign;
  reg                 add_preShifter_output_rData_rs2_special;
  reg        [4:0]    add_preShifter_output_rData_rd;
  reg        [2:0]    add_preShifter_output_rData_roundMode;
  reg        [0:0]    add_preShifter_output_rData_format;
  reg                 add_preShifter_output_rData_needCommit;
  reg                 add_preShifter_output_rData_absRs1Bigger;
  reg                 add_preShifter_output_rData_rs1ExponentBigger;
  wire                when_Stream_l375_15;
  wire                add_shifter_output_valid;
  reg                 add_shifter_output_ready;
  wire       [0:0]    add_shifter_output_payload_source;
  wire       [53:0]   add_shifter_output_payload_rs1_mantissa;
  wire       [11:0]   add_shifter_output_payload_rs1_exponent;
  wire                add_shifter_output_payload_rs1_sign;
  wire                add_shifter_output_payload_rs1_special;
  wire       [53:0]   add_shifter_output_payload_rs2_mantissa;
  wire       [11:0]   add_shifter_output_payload_rs2_exponent;
  wire                add_shifter_output_payload_rs2_sign;
  wire                add_shifter_output_payload_rs2_special;
  wire       [4:0]    add_shifter_output_payload_rd;
  wire       [2:0]    add_shifter_output_payload_roundMode;
  wire       [0:0]    add_shifter_output_payload_format;
  wire                add_shifter_output_payload_needCommit;
  wire                add_shifter_output_payload_xSign;
  wire                add_shifter_output_payload_ySign;
  wire       [54:0]   add_shifter_output_payload_xMantissa;
  wire       [54:0]   add_shifter_output_payload_yMantissa;
  wire       [11:0]   add_shifter_output_payload_xyExponent;
  wire                add_shifter_output_payload_xySign;
  wire                add_shifter_output_payload_roundingScrap;
  wire       [12:0]   add_shifter_exp21;
  wire       [12:0]   _zz_add_shifter_shiftBy;
  wire       [12:0]   add_shifter_shiftBy;
  wire                add_shifter_shiftOverflow;
  wire                add_shifter_passThrough;
  wire                add_shifter_xySign;
  wire       [54:0]   add_shifter_xMantissa;
  wire       [54:0]   add_shifter_yMantissaUnshifted;
  wire       [54:0]   add_shifter_yMantissa;
  reg                 add_shifter_roundingScrap;
  wire                when_FpuCore_l1419;
  wire                when_FpuCore_l1419_1;
  wire                when_FpuCore_l1419_2;
  wire                when_FpuCore_l1419_3;
  wire                when_FpuCore_l1419_4;
  wire                when_FpuCore_l1419_5;
  wire                when_FpuCore_l1424;
  wire                add_math_input_valid;
  wire                add_math_input_ready;
  wire       [0:0]    add_math_input_payload_source;
  wire       [53:0]   add_math_input_payload_rs1_mantissa;
  wire       [11:0]   add_math_input_payload_rs1_exponent;
  wire                add_math_input_payload_rs1_sign;
  wire                add_math_input_payload_rs1_special;
  wire       [53:0]   add_math_input_payload_rs2_mantissa;
  wire       [11:0]   add_math_input_payload_rs2_exponent;
  wire                add_math_input_payload_rs2_sign;
  wire                add_math_input_payload_rs2_special;
  wire       [4:0]    add_math_input_payload_rd;
  wire       [2:0]    add_math_input_payload_roundMode;
  wire       [0:0]    add_math_input_payload_format;
  wire                add_math_input_payload_needCommit;
  wire                add_math_input_payload_xSign;
  wire                add_math_input_payload_ySign;
  wire       [54:0]   add_math_input_payload_xMantissa;
  wire       [54:0]   add_math_input_payload_yMantissa;
  wire       [11:0]   add_math_input_payload_xyExponent;
  wire                add_math_input_payload_xySign;
  wire                add_math_input_payload_roundingScrap;
  reg                 add_shifter_output_rValid;
  reg        [0:0]    add_shifter_output_rData_source;
  reg        [53:0]   add_shifter_output_rData_rs1_mantissa;
  reg        [11:0]   add_shifter_output_rData_rs1_exponent;
  reg                 add_shifter_output_rData_rs1_sign;
  reg                 add_shifter_output_rData_rs1_special;
  reg        [53:0]   add_shifter_output_rData_rs2_mantissa;
  reg        [11:0]   add_shifter_output_rData_rs2_exponent;
  reg                 add_shifter_output_rData_rs2_sign;
  reg                 add_shifter_output_rData_rs2_special;
  reg        [4:0]    add_shifter_output_rData_rd;
  reg        [2:0]    add_shifter_output_rData_roundMode;
  reg        [0:0]    add_shifter_output_rData_format;
  reg                 add_shifter_output_rData_needCommit;
  reg                 add_shifter_output_rData_xSign;
  reg                 add_shifter_output_rData_ySign;
  reg        [54:0]   add_shifter_output_rData_xMantissa;
  reg        [54:0]   add_shifter_output_rData_yMantissa;
  reg        [11:0]   add_shifter_output_rData_xyExponent;
  reg                 add_shifter_output_rData_xySign;
  reg                 add_shifter_output_rData_roundingScrap;
  wire                when_Stream_l375_16;
  wire                add_math_output_valid;
  reg                 add_math_output_ready;
  wire       [0:0]    add_math_output_payload_source;
  wire       [53:0]   add_math_output_payload_rs1_mantissa;
  wire       [11:0]   add_math_output_payload_rs1_exponent;
  wire                add_math_output_payload_rs1_sign;
  wire                add_math_output_payload_rs1_special;
  wire       [53:0]   add_math_output_payload_rs2_mantissa;
  wire       [11:0]   add_math_output_payload_rs2_exponent;
  wire                add_math_output_payload_rs2_sign;
  wire                add_math_output_payload_rs2_special;
  wire       [4:0]    add_math_output_payload_rd;
  wire       [2:0]    add_math_output_payload_roundMode;
  wire       [0:0]    add_math_output_payload_format;
  wire                add_math_output_payload_needCommit;
  wire                add_math_output_payload_xSign;
  wire                add_math_output_payload_ySign;
  wire       [54:0]   add_math_output_payload_xMantissa;
  wire       [54:0]   add_math_output_payload_yMantissa;
  wire       [11:0]   add_math_output_payload_xyExponent;
  wire                add_math_output_payload_xySign;
  wire                add_math_output_payload_roundingScrap;
  wire       [55:0]   add_math_output_payload_xyMantissa;
  wire       [55:0]   add_math_xSigned;
  wire       [55:0]   add_math_ySigned;
  wire                add_oh_input_valid;
  wire                add_oh_input_ready;
  wire       [0:0]    add_oh_input_payload_source;
  wire       [53:0]   add_oh_input_payload_rs1_mantissa;
  wire       [11:0]   add_oh_input_payload_rs1_exponent;
  wire                add_oh_input_payload_rs1_sign;
  wire                add_oh_input_payload_rs1_special;
  wire       [53:0]   add_oh_input_payload_rs2_mantissa;
  wire       [11:0]   add_oh_input_payload_rs2_exponent;
  wire                add_oh_input_payload_rs2_sign;
  wire                add_oh_input_payload_rs2_special;
  wire       [4:0]    add_oh_input_payload_rd;
  wire       [2:0]    add_oh_input_payload_roundMode;
  wire       [0:0]    add_oh_input_payload_format;
  wire                add_oh_input_payload_needCommit;
  wire                add_oh_input_payload_xSign;
  wire                add_oh_input_payload_ySign;
  wire       [54:0]   add_oh_input_payload_xMantissa;
  wire       [54:0]   add_oh_input_payload_yMantissa;
  wire       [11:0]   add_oh_input_payload_xyExponent;
  wire                add_oh_input_payload_xySign;
  wire                add_oh_input_payload_roundingScrap;
  wire       [55:0]   add_oh_input_payload_xyMantissa;
  reg                 add_math_output_rValid;
  reg        [0:0]    add_math_output_rData_source;
  reg        [53:0]   add_math_output_rData_rs1_mantissa;
  reg        [11:0]   add_math_output_rData_rs1_exponent;
  reg                 add_math_output_rData_rs1_sign;
  reg                 add_math_output_rData_rs1_special;
  reg        [53:0]   add_math_output_rData_rs2_mantissa;
  reg        [11:0]   add_math_output_rData_rs2_exponent;
  reg                 add_math_output_rData_rs2_sign;
  reg                 add_math_output_rData_rs2_special;
  reg        [4:0]    add_math_output_rData_rd;
  reg        [2:0]    add_math_output_rData_roundMode;
  reg        [0:0]    add_math_output_rData_format;
  reg                 add_math_output_rData_needCommit;
  reg                 add_math_output_rData_xSign;
  reg                 add_math_output_rData_ySign;
  reg        [54:0]   add_math_output_rData_xMantissa;
  reg        [54:0]   add_math_output_rData_yMantissa;
  reg        [11:0]   add_math_output_rData_xyExponent;
  reg                 add_math_output_rData_xySign;
  reg                 add_math_output_rData_roundingScrap;
  reg        [55:0]   add_math_output_rData_xyMantissa;
  wire                when_Stream_l375_17;
  wire                add_oh_input_fire;
  wire                _zz_when_FpuCore_l221_1;
  wire                when_FpuCore_l221_8;
  wire                when_FpuCore_l221_9;
  wire                add_oh_isCommited;
  wire                _zz_add_oh_input_ready;
  wire                add_oh_output_valid;
  reg                 add_oh_output_ready;
  wire       [0:0]    add_oh_output_payload_source;
  wire       [53:0]   add_oh_output_payload_rs1_mantissa;
  wire       [11:0]   add_oh_output_payload_rs1_exponent;
  wire                add_oh_output_payload_rs1_sign;
  wire                add_oh_output_payload_rs1_special;
  wire       [53:0]   add_oh_output_payload_rs2_mantissa;
  wire       [11:0]   add_oh_output_payload_rs2_exponent;
  wire                add_oh_output_payload_rs2_sign;
  wire                add_oh_output_payload_rs2_special;
  wire       [4:0]    add_oh_output_payload_rd;
  wire       [2:0]    add_oh_output_payload_roundMode;
  wire       [0:0]    add_oh_output_payload_format;
  wire                add_oh_output_payload_needCommit;
  wire                add_oh_output_payload_xSign;
  wire                add_oh_output_payload_ySign;
  wire       [54:0]   add_oh_output_payload_xMantissa;
  wire       [54:0]   add_oh_output_payload_yMantissa;
  wire       [11:0]   add_oh_output_payload_xyExponent;
  wire                add_oh_output_payload_xySign;
  wire                add_oh_output_payload_roundingScrap;
  wire       [55:0]   add_oh_output_payload_xyMantissa;
  wire       [5:0]    add_oh_output_payload_shift;
  wire       [55:0]   _zz_add_oh_shift;
  wire       [55:0]   _zz_add_oh_shift_1;
  wire                _zz_add_oh_shift_2;
  wire                _zz_add_oh_shift_3;
  wire                _zz_add_oh_shift_4;
  wire                _zz_add_oh_shift_5;
  wire                _zz_add_oh_shift_6;
  wire                _zz_add_oh_shift_7;
  wire                _zz_add_oh_shift_8;
  wire                _zz_add_oh_shift_9;
  wire                _zz_add_oh_shift_10;
  wire                _zz_add_oh_shift_11;
  wire                _zz_add_oh_shift_12;
  wire                _zz_add_oh_shift_13;
  wire                _zz_add_oh_shift_14;
  wire                _zz_add_oh_shift_15;
  wire                _zz_add_oh_shift_16;
  wire                _zz_add_oh_shift_17;
  wire                _zz_add_oh_shift_18;
  wire                _zz_add_oh_shift_19;
  wire                _zz_add_oh_shift_20;
  wire                _zz_add_oh_shift_21;
  wire                _zz_add_oh_shift_22;
  wire                _zz_add_oh_shift_23;
  wire                _zz_add_oh_shift_24;
  wire                _zz_add_oh_shift_25;
  wire                _zz_add_oh_shift_26;
  wire                _zz_add_oh_shift_27;
  wire                _zz_add_oh_shift_28;
  wire                _zz_add_oh_shift_29;
  wire                _zz_add_oh_shift_30;
  wire                _zz_add_oh_shift_31;
  wire                _zz_add_oh_shift_32;
  wire                _zz_add_oh_shift_33;
  wire                _zz_add_oh_shift_34;
  wire                _zz_add_oh_shift_35;
  wire                _zz_add_oh_shift_36;
  wire                _zz_add_oh_shift_37;
  wire                _zz_add_oh_shift_38;
  wire                _zz_add_oh_shift_39;
  wire                _zz_add_oh_shift_40;
  wire                _zz_add_oh_shift_41;
  wire                _zz_add_oh_shift_42;
  wire                _zz_add_oh_shift_43;
  wire                _zz_add_oh_shift_44;
  wire                _zz_add_oh_shift_45;
  wire                _zz_add_oh_shift_46;
  wire                _zz_add_oh_shift_47;
  wire                _zz_add_oh_shift_48;
  wire                _zz_add_oh_shift_49;
  wire                _zz_add_oh_shift_50;
  wire                _zz_add_oh_shift_51;
  wire                _zz_add_oh_shift_52;
  wire                _zz_add_oh_shift_53;
  wire                _zz_add_oh_shift_54;
  wire                _zz_add_oh_shift_55;
  wire                _zz_add_oh_shift_56;
  wire       [5:0]    add_oh_shift;
  wire                add_norm_input_valid;
  wire                add_norm_input_ready;
  wire       [0:0]    add_norm_input_payload_source;
  wire       [53:0]   add_norm_input_payload_rs1_mantissa;
  wire       [11:0]   add_norm_input_payload_rs1_exponent;
  wire                add_norm_input_payload_rs1_sign;
  wire                add_norm_input_payload_rs1_special;
  wire       [53:0]   add_norm_input_payload_rs2_mantissa;
  wire       [11:0]   add_norm_input_payload_rs2_exponent;
  wire                add_norm_input_payload_rs2_sign;
  wire                add_norm_input_payload_rs2_special;
  wire       [4:0]    add_norm_input_payload_rd;
  wire       [2:0]    add_norm_input_payload_roundMode;
  wire       [0:0]    add_norm_input_payload_format;
  wire                add_norm_input_payload_needCommit;
  wire                add_norm_input_payload_xSign;
  wire                add_norm_input_payload_ySign;
  wire       [54:0]   add_norm_input_payload_xMantissa;
  wire       [54:0]   add_norm_input_payload_yMantissa;
  wire       [11:0]   add_norm_input_payload_xyExponent;
  wire                add_norm_input_payload_xySign;
  wire                add_norm_input_payload_roundingScrap;
  wire       [55:0]   add_norm_input_payload_xyMantissa;
  wire       [5:0]    add_norm_input_payload_shift;
  reg                 add_oh_output_rValid;
  reg        [0:0]    add_oh_output_rData_source;
  reg        [53:0]   add_oh_output_rData_rs1_mantissa;
  reg        [11:0]   add_oh_output_rData_rs1_exponent;
  reg                 add_oh_output_rData_rs1_sign;
  reg                 add_oh_output_rData_rs1_special;
  reg        [53:0]   add_oh_output_rData_rs2_mantissa;
  reg        [11:0]   add_oh_output_rData_rs2_exponent;
  reg                 add_oh_output_rData_rs2_sign;
  reg                 add_oh_output_rData_rs2_special;
  reg        [4:0]    add_oh_output_rData_rd;
  reg        [2:0]    add_oh_output_rData_roundMode;
  reg        [0:0]    add_oh_output_rData_format;
  reg                 add_oh_output_rData_needCommit;
  reg                 add_oh_output_rData_xSign;
  reg                 add_oh_output_rData_ySign;
  reg        [54:0]   add_oh_output_rData_xMantissa;
  reg        [54:0]   add_oh_output_rData_yMantissa;
  reg        [11:0]   add_oh_output_rData_xyExponent;
  reg                 add_oh_output_rData_xySign;
  reg                 add_oh_output_rData_roundingScrap;
  reg        [55:0]   add_oh_output_rData_xyMantissa;
  reg        [5:0]    add_oh_output_rData_shift;
  wire                when_Stream_l375_18;
  wire                add_norm_output_valid;
  wire                add_norm_output_ready;
  wire       [0:0]    add_norm_output_payload_source;
  wire       [53:0]   add_norm_output_payload_rs1_mantissa;
  wire       [11:0]   add_norm_output_payload_rs1_exponent;
  wire                add_norm_output_payload_rs1_sign;
  wire                add_norm_output_payload_rs1_special;
  wire       [53:0]   add_norm_output_payload_rs2_mantissa;
  wire       [11:0]   add_norm_output_payload_rs2_exponent;
  wire                add_norm_output_payload_rs2_sign;
  wire                add_norm_output_payload_rs2_special;
  wire       [4:0]    add_norm_output_payload_rd;
  wire       [2:0]    add_norm_output_payload_roundMode;
  wire       [0:0]    add_norm_output_payload_format;
  wire                add_norm_output_payload_needCommit;
  wire       [55:0]   add_norm_output_payload_mantissa;
  wire       [12:0]   add_norm_output_payload_exponent;
  wire                add_norm_output_payload_infinityNan;
  wire                add_norm_output_payload_forceNan;
  wire                add_norm_output_payload_forceZero;
  wire                add_norm_output_payload_forceInfinity;
  wire                add_norm_output_payload_xySign;
  wire                add_norm_output_payload_roundingScrap;
  wire                add_norm_output_payload_xyMantissaZero;
  wire                add_result_input_valid;
  wire                add_result_input_ready;
  wire       [0:0]    add_result_input_payload_source;
  wire       [53:0]   add_result_input_payload_rs1_mantissa;
  wire       [11:0]   add_result_input_payload_rs1_exponent;
  wire                add_result_input_payload_rs1_sign;
  wire                add_result_input_payload_rs1_special;
  wire       [53:0]   add_result_input_payload_rs2_mantissa;
  wire       [11:0]   add_result_input_payload_rs2_exponent;
  wire                add_result_input_payload_rs2_sign;
  wire                add_result_input_payload_rs2_special;
  wire       [4:0]    add_result_input_payload_rd;
  wire       [2:0]    add_result_input_payload_roundMode;
  wire       [0:0]    add_result_input_payload_format;
  wire                add_result_input_payload_needCommit;
  wire       [55:0]   add_result_input_payload_mantissa;
  wire       [12:0]   add_result_input_payload_exponent;
  wire                add_result_input_payload_infinityNan;
  wire                add_result_input_payload_forceNan;
  wire                add_result_input_payload_forceZero;
  wire                add_result_input_payload_forceInfinity;
  wire                add_result_input_payload_xySign;
  wire                add_result_input_payload_roundingScrap;
  wire                add_result_input_payload_xyMantissaZero;
  wire                add_result_output_valid;
  wire                add_result_output_ready;
  wire       [0:0]    add_result_output_payload_source;
  wire       [4:0]    add_result_output_payload_rd;
  reg        [52:0]   add_result_output_payload_value_mantissa;
  reg        [11:0]   add_result_output_payload_value_exponent;
  reg                 add_result_output_payload_value_sign;
  reg                 add_result_output_payload_value_special;
  wire                add_result_output_payload_scrap;
  wire       [2:0]    add_result_output_payload_roundMode;
  wire       [0:0]    add_result_output_payload_format;
  wire                add_result_output_payload_NV;
  wire                add_result_output_payload_DZ;
  wire                when_FpuCore_l1513;
  wire                when_FpuCore_l1516;
  wire                load_s1_output_m2sPipe_valid;
  wire                load_s1_output_m2sPipe_ready;
  wire       [0:0]    load_s1_output_m2sPipe_payload_source;
  wire       [4:0]    load_s1_output_m2sPipe_payload_rd;
  wire       [52:0]   load_s1_output_m2sPipe_payload_value_mantissa;
  wire       [11:0]   load_s1_output_m2sPipe_payload_value_exponent;
  wire                load_s1_output_m2sPipe_payload_value_sign;
  wire                load_s1_output_m2sPipe_payload_value_special;
  wire                load_s1_output_m2sPipe_payload_scrap;
  wire       [2:0]    load_s1_output_m2sPipe_payload_roundMode;
  wire       [0:0]    load_s1_output_m2sPipe_payload_format;
  wire                load_s1_output_m2sPipe_payload_NV;
  wire                load_s1_output_m2sPipe_payload_DZ;
  reg                 load_s1_output_rValid;
  reg        [0:0]    load_s1_output_rData_source;
  reg        [4:0]    load_s1_output_rData_rd;
  reg        [52:0]   load_s1_output_rData_value_mantissa;
  reg        [11:0]   load_s1_output_rData_value_exponent;
  reg                 load_s1_output_rData_value_sign;
  reg                 load_s1_output_rData_value_special;
  reg                 load_s1_output_rData_scrap;
  reg        [2:0]    load_s1_output_rData_roundMode;
  reg        [0:0]    load_s1_output_rData_format;
  reg                 load_s1_output_rData_NV;
  reg                 load_s1_output_rData_DZ;
  wire                when_Stream_l375_19;
  wire                shortPip_output_m2sPipe_valid;
  wire                shortPip_output_m2sPipe_ready;
  wire       [0:0]    shortPip_output_m2sPipe_payload_source;
  wire       [4:0]    shortPip_output_m2sPipe_payload_rd;
  wire       [52:0]   shortPip_output_m2sPipe_payload_value_mantissa;
  wire       [11:0]   shortPip_output_m2sPipe_payload_value_exponent;
  wire                shortPip_output_m2sPipe_payload_value_sign;
  wire                shortPip_output_m2sPipe_payload_value_special;
  wire                shortPip_output_m2sPipe_payload_scrap;
  wire       [2:0]    shortPip_output_m2sPipe_payload_roundMode;
  wire       [0:0]    shortPip_output_m2sPipe_payload_format;
  wire                shortPip_output_m2sPipe_payload_NV;
  wire                shortPip_output_m2sPipe_payload_DZ;
  reg                 shortPip_output_rValid;
  reg        [0:0]    shortPip_output_rData_source;
  reg        [4:0]    shortPip_output_rData_rd;
  reg        [52:0]   shortPip_output_rData_value_mantissa;
  reg        [11:0]   shortPip_output_rData_value_exponent;
  reg                 shortPip_output_rData_value_sign;
  reg                 shortPip_output_rData_value_special;
  reg                 shortPip_output_rData_scrap;
  reg        [2:0]    shortPip_output_rData_roundMode;
  reg        [0:0]    shortPip_output_rData_format;
  reg                 shortPip_output_rData_NV;
  reg                 shortPip_output_rData_DZ;
  wire                when_Stream_l375_20;
  wire                streamArbiter_10_io_output_combStage_valid;
  wire                streamArbiter_10_io_output_combStage_ready;
  wire       [0:0]    streamArbiter_10_io_output_combStage_payload_source;
  wire       [4:0]    streamArbiter_10_io_output_combStage_payload_rd;
  wire       [52:0]   streamArbiter_10_io_output_combStage_payload_value_mantissa;
  wire       [11:0]   streamArbiter_10_io_output_combStage_payload_value_exponent;
  wire                streamArbiter_10_io_output_combStage_payload_value_sign;
  wire                streamArbiter_10_io_output_combStage_payload_value_special;
  wire                streamArbiter_10_io_output_combStage_payload_scrap;
  wire       [2:0]    streamArbiter_10_io_output_combStage_payload_roundMode;
  wire       [0:0]    streamArbiter_10_io_output_combStage_payload_format;
  wire                streamArbiter_10_io_output_combStage_payload_NV;
  wire                streamArbiter_10_io_output_combStage_payload_DZ;
  wire                merge_arbitrated_valid;
  wire       [0:0]    merge_arbitrated_payload_source;
  wire       [4:0]    merge_arbitrated_payload_rd;
  wire       [52:0]   merge_arbitrated_payload_value_mantissa;
  wire       [11:0]   merge_arbitrated_payload_value_exponent;
  wire                merge_arbitrated_payload_value_sign;
  wire                merge_arbitrated_payload_value_special;
  wire                merge_arbitrated_payload_scrap;
  wire       [2:0]    merge_arbitrated_payload_roundMode;
  wire       [0:0]    merge_arbitrated_payload_format;
  wire                merge_arbitrated_payload_NV;
  wire                merge_arbitrated_payload_DZ;
  reg                 roundFront_input_valid;
  reg        [0:0]    roundFront_input_payload_source;
  reg        [4:0]    roundFront_input_payload_rd;
  reg        [52:0]   roundFront_input_payload_value_mantissa;
  reg        [11:0]   roundFront_input_payload_value_exponent;
  reg                 roundFront_input_payload_value_sign;
  reg                 roundFront_input_payload_value_special;
  reg                 roundFront_input_payload_scrap;
  reg        [2:0]    roundFront_input_payload_roundMode;
  reg        [0:0]    roundFront_input_payload_format;
  reg                 roundFront_input_payload_NV;
  reg                 roundFront_input_payload_DZ;
  wire                roundFront_output_valid;
  wire       [0:0]    roundFront_output_payload_source;
  wire       [4:0]    roundFront_output_payload_rd;
  wire       [52:0]   roundFront_output_payload_value_mantissa;
  wire       [11:0]   roundFront_output_payload_value_exponent;
  wire                roundFront_output_payload_value_sign;
  wire                roundFront_output_payload_value_special;
  wire                roundFront_output_payload_scrap;
  wire       [2:0]    roundFront_output_payload_roundMode;
  wire       [0:0]    roundFront_output_payload_format;
  wire                roundFront_output_payload_NV;
  wire                roundFront_output_payload_DZ;
  wire                roundFront_output_payload_mantissaIncrement;
  wire       [1:0]    roundFront_output_payload_roundAdjusted;
  wire       [53:0]   roundFront_output_payload_exactMask;
  wire       [53:0]   roundFront_manAggregate;
  wire       [10:0]   roundFront_expBase;
  wire       [12:0]   roundFront_expDif;
  wire                roundFront_expSubnormal;
  wire       [12:0]   roundFront_discardCount;
  wire                when_FpuCore_l1551;
  wire       [5:0]    roundFront_discardCountTrunk;
  reg        [53:0]   roundFront_exactMask;
  reg        [1:0]    roundFront_roundAdjusted;
  reg                 roundFront_rneBit;
  wire                when_FpuCore_l1559;
  reg                 _zz_roundFront_mantissaIncrement;
  wire                roundFront_mantissaIncrement;
  reg                 roundBack_input_valid;
  reg        [0:0]    roundBack_input_payload_source;
  reg        [4:0]    roundBack_input_payload_rd;
  reg        [52:0]   roundBack_input_payload_value_mantissa;
  reg        [11:0]   roundBack_input_payload_value_exponent;
  reg                 roundBack_input_payload_value_sign;
  reg                 roundBack_input_payload_value_special;
  reg                 roundBack_input_payload_scrap;
  reg        [2:0]    roundBack_input_payload_roundMode;
  reg        [0:0]    roundBack_input_payload_format;
  reg                 roundBack_input_payload_NV;
  reg                 roundBack_input_payload_DZ;
  reg                 roundBack_input_payload_mantissaIncrement;
  reg        [1:0]    roundBack_input_payload_roundAdjusted;
  reg        [53:0]   roundBack_input_payload_exactMask;
  wire                roundBack_output_valid;
  wire       [0:0]    roundBack_output_payload_source;
  wire       [4:0]    roundBack_output_payload_rd;
  wire       [51:0]   roundBack_output_payload_value_mantissa;
  wire       [11:0]   roundBack_output_payload_value_exponent;
  wire                roundBack_output_payload_value_sign;
  wire                roundBack_output_payload_value_special;
  wire       [0:0]    roundBack_output_payload_format;
  wire                roundBack_output_payload_NV;
  wire                roundBack_output_payload_NX;
  wire                roundBack_output_payload_OF;
  wire                roundBack_output_payload_UF;
  wire                roundBack_output_payload_DZ;
  wire                roundBack_output_payload_write;
  wire       [51:0]   roundBack_math_mantissa;
  wire       [11:0]   roundBack_math_exponent;
  wire                roundBack_math_sign;
  wire                roundBack_math_special;
  wire       [51:0]   roundBack_adderMantissa;
  (* keep , syn_keep *) wire       [51:0]   roundBack_adderRightOp /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [63:0]   _zz_roundBack_adder /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [0:0]    _zz_roundBack_adder_1 /* synthesis syn_keep = 1 */ ;
  (* keep , syn_keep *) wire       [63:0]   roundBack_adder /* synthesis syn_keep = 1 */ ;
  wire       [63:0]   roundBack_masked;
  reg        [51:0]   roundBack_patched_mantissa;
  reg        [11:0]   roundBack_patched_exponent;
  wire                roundBack_patched_sign;
  reg                 roundBack_patched_special;
  reg                 roundBack_nx;
  reg                 roundBack_of;
  reg                 roundBack_uf;
  wire       [10:0]   roundBack_ufSubnormalThreshold;
  wire       [10:0]   roundBack_ufThreshold;
  wire       [11:0]   roundBack_ofThreshold;
  reg        [2:0]    roundBack_threshold;
  reg        [2:0]    roundBack_borringRound;
  wire                when_FpuCore_l1613;
  wire                roundBack_borringCase;
  wire                when_FpuCore_l1616;
  wire                when_FpuCore_l1619;
  reg                 when_FpuCore_l1629;
  wire                when_FpuCore_l1638;
  reg                 when_FpuCore_l1648;
  wire                when_FpuCore_l1657;
  wire                roundBack_writes_0;
  wire                roundBack_writes_1;
  wire                roundBack_write;
  reg                 writeback_input_valid;
  reg        [0:0]    writeback_input_payload_source;
  reg        [4:0]    writeback_input_payload_rd;
  reg        [51:0]   writeback_input_payload_value_mantissa;
  reg        [11:0]   writeback_input_payload_value_exponent;
  reg                 writeback_input_payload_value_sign;
  reg                 writeback_input_payload_value_special;
  reg        [0:0]    writeback_input_payload_format;
  reg                 writeback_input_payload_NV;
  reg                 writeback_input_payload_NX;
  reg                 writeback_input_payload_OF;
  reg                 writeback_input_payload_UF;
  reg                 writeback_input_payload_DZ;
  reg                 writeback_input_payload_write;
  wire                when_FpuCore_l1689;
  wire                when_FpuCore_l1689_1;
  wire                writeback_port_valid;
  wire       [5:0]    writeback_port_payload_address;
  reg        [51:0]   writeback_port_payload_data_value_mantissa;
  wire       [11:0]   writeback_port_payload_data_value_exponent;
  wire                writeback_port_payload_data_value_sign;
  wire                writeback_port_payload_data_value_special;
  wire                writeback_port_payload_data_boxed;
  `ifndef SYNTHESIS
  reg [63:0] io_port_0_cmd_payload_opcode_string;
  reg [47:0] io_port_0_cmd_payload_format_string;
  reg [23:0] io_port_0_cmd_payload_roundMode_string;
  reg [63:0] io_port_0_commit_payload_opcode_string;
  reg [63:0] io_port_1_cmd_payload_opcode_string;
  reg [47:0] io_port_1_cmd_payload_format_string;
  reg [23:0] io_port_1_cmd_payload_roundMode_string;
  reg [63:0] io_port_1_commit_payload_opcode_string;
  reg [63:0] commitFork_load_0_payload_opcode_string;
  reg [63:0] commitFork_load_1_payload_opcode_string;
  reg [63:0] commitFork_commit_0_payload_opcode_string;
  reg [63:0] commitFork_commit_1_payload_opcode_string;
  reg [63:0] streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string;
  reg [63:0] streamFork_3_io_outputs_1_rData_opcode_string;
  reg [63:0] _zz_payload_opcode_string;
  reg [63:0] streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string;
  reg [63:0] streamFork_4_io_outputs_1_rData_opcode_string;
  reg [63:0] _zz_payload_opcode_1_string;
  reg [63:0] _zz_commitLogic_0_input_payload_opcode_string;
  reg [63:0] commitLogic_0_input_payload_opcode_string;
  reg [63:0] _zz_commitLogic_1_input_payload_opcode_string;
  reg [63:0] commitLogic_1_input_payload_opcode_string;
  reg [63:0] scheduler_0_input_payload_opcode_string;
  reg [47:0] scheduler_0_input_payload_format_string;
  reg [23:0] scheduler_0_input_payload_roundMode_string;
  reg [63:0] io_port_0_cmd_rData_opcode_string;
  reg [47:0] io_port_0_cmd_rData_format_string;
  reg [23:0] io_port_0_cmd_rData_roundMode_string;
  reg [63:0] _zz_scheduler_0_input_payload_opcode_string;
  reg [47:0] _zz_scheduler_0_input_payload_format_string;
  reg [23:0] _zz_scheduler_0_input_payload_roundMode_string;
  reg [63:0] scheduler_0_output_payload_opcode_string;
  reg [47:0] scheduler_0_output_payload_format_string;
  reg [23:0] scheduler_0_output_payload_roundMode_string;
  reg [63:0] scheduler_1_input_payload_opcode_string;
  reg [47:0] scheduler_1_input_payload_format_string;
  reg [23:0] scheduler_1_input_payload_roundMode_string;
  reg [63:0] io_port_1_cmd_rData_opcode_string;
  reg [47:0] io_port_1_cmd_rData_format_string;
  reg [23:0] io_port_1_cmd_rData_roundMode_string;
  reg [63:0] _zz_scheduler_1_input_payload_opcode_string;
  reg [47:0] _zz_scheduler_1_input_payload_format_string;
  reg [23:0] _zz_scheduler_1_input_payload_roundMode_string;
  reg [63:0] scheduler_1_output_payload_opcode_string;
  reg [47:0] scheduler_1_output_payload_format_string;
  reg [23:0] scheduler_1_output_payload_roundMode_string;
  reg [63:0] scheduler_0_output_m2sPipe_payload_opcode_string;
  reg [47:0] scheduler_0_output_m2sPipe_payload_format_string;
  reg [23:0] scheduler_0_output_m2sPipe_payload_roundMode_string;
  reg [63:0] scheduler_0_output_rData_opcode_string;
  reg [47:0] scheduler_0_output_rData_format_string;
  reg [23:0] scheduler_0_output_rData_roundMode_string;
  reg [63:0] scheduler_1_output_m2sPipe_payload_opcode_string;
  reg [47:0] scheduler_1_output_m2sPipe_payload_format_string;
  reg [23:0] scheduler_1_output_m2sPipe_payload_roundMode_string;
  reg [63:0] scheduler_1_output_rData_opcode_string;
  reg [47:0] scheduler_1_output_rData_format_string;
  reg [23:0] scheduler_1_output_rData_roundMode_string;
  reg [63:0] cmdArbiter_output_payload_opcode_string;
  reg [23:0] cmdArbiter_output_payload_roundMode_string;
  reg [47:0] cmdArbiter_output_payload_format_string;
  reg [63:0] read_s0_payload_opcode_string;
  reg [23:0] read_s0_payload_roundMode_string;
  reg [47:0] read_s0_payload_format_string;
  reg [63:0] read_s1_payload_opcode_string;
  reg [23:0] read_s1_payload_roundMode_string;
  reg [47:0] read_s1_payload_format_string;
  reg [63:0] read_s0_rData_opcode_string;
  reg [23:0] read_s0_rData_roundMode_string;
  reg [47:0] read_s0_rData_format_string;
  reg [63:0] read_output_payload_opcode_string;
  reg [23:0] read_output_payload_roundMode_string;
  reg [47:0] read_output_payload_format_string;
  reg [47:0] _zz_read_output_payload_format_string;
  reg [63:0] decode_input_payload_opcode_string;
  reg [23:0] decode_input_payload_roundMode_string;
  reg [47:0] decode_input_payload_format_string;
  reg [23:0] decode_load_payload_roundMode_string;
  reg [47:0] decode_load_payload_format_string;
  reg [63:0] decode_shortPip_payload_opcode_string;
  reg [23:0] decode_shortPip_payload_roundMode_string;
  reg [47:0] decode_shortPip_payload_format_string;
  reg [23:0] decode_divSqrt_payload_roundMode_string;
  reg [47:0] decode_divSqrt_payload_format_string;
  reg [23:0] decode_div_payload_roundMode_string;
  reg [47:0] decode_div_payload_format_string;
  reg [23:0] decode_sqrt_payload_roundMode_string;
  reg [47:0] decode_sqrt_payload_format_string;
  reg [23:0] decode_mul_payload_roundMode_string;
  reg [47:0] decode_mul_payload_format_string;
  reg [23:0] decode_divSqrtToMul_payload_roundMode_string;
  reg [47:0] decode_divSqrtToMul_payload_format_string;
  reg [23:0] decode_add_payload_roundMode_string;
  reg [47:0] decode_add_payload_format_string;
  reg [23:0] decode_mulToAdd_payload_roundMode_string;
  reg [47:0] decode_mulToAdd_payload_format_string;
  reg [23:0] decode_load_s2mPipe_payload_roundMode_string;
  reg [47:0] decode_load_s2mPipe_payload_format_string;
  reg [23:0] decode_load_rData_roundMode_string;
  reg [47:0] decode_load_rData_format_string;
  reg [23:0] _zz_decode_load_s2mPipe_payload_roundMode_string;
  reg [47:0] _zz_decode_load_s2mPipe_payload_format_string;
  reg [23:0] decode_load_s2mPipe_m2sPipe_payload_roundMode_string;
  reg [47:0] decode_load_s2mPipe_m2sPipe_payload_format_string;
  reg [23:0] decode_load_s2mPipe_rData_roundMode_string;
  reg [47:0] decode_load_s2mPipe_rData_format_string;
  reg [23:0] load_s0_input_payload_roundMode_string;
  reg [47:0] load_s0_input_payload_format_string;
  reg [23:0] decode_load_s2mPipe_m2sPipe_rData_roundMode_string;
  reg [47:0] decode_load_s2mPipe_m2sPipe_rData_format_string;
  reg [63:0] load_s0_filtred_0_payload_opcode_string;
  reg [63:0] load_s0_filtred_1_payload_opcode_string;
  reg [23:0] load_s0_output_payload_roundMode_string;
  reg [47:0] load_s0_output_payload_format_string;
  reg [23:0] load_s1_input_payload_roundMode_string;
  reg [47:0] load_s1_input_payload_format_string;
  reg [23:0] load_s0_output_rData_roundMode_string;
  reg [47:0] load_s0_output_rData_format_string;
  reg [23:0] load_s1_output_payload_roundMode_string;
  reg [47:0] load_s1_output_payload_format_string;
  reg [63:0] shortPip_input_payload_opcode_string;
  reg [23:0] shortPip_input_payload_roundMode_string;
  reg [47:0] shortPip_input_payload_format_string;
  reg [63:0] decode_shortPip_rData_opcode_string;
  reg [23:0] decode_shortPip_rData_roundMode_string;
  reg [47:0] decode_shortPip_rData_format_string;
  reg [23:0] shortPip_rfOutput_payload_roundMode_string;
  reg [47:0] shortPip_rfOutput_payload_format_string;
  reg [23:0] shortPip_output_payload_roundMode_string;
  reg [47:0] shortPip_output_payload_format_string;
  reg [47:0] _zz_shortPip_rfOutput_payload_format_string;
  reg [23:0] mul_preMul_input_payload_roundMode_string;
  reg [47:0] mul_preMul_input_payload_format_string;
  reg [23:0] decode_mul_rData_roundMode_string;
  reg [47:0] decode_mul_rData_format_string;
  reg [23:0] mul_preMul_output_payload_roundMode_string;
  reg [47:0] mul_preMul_output_payload_format_string;
  reg [23:0] mul_mul_input_payload_roundMode_string;
  reg [47:0] mul_mul_input_payload_format_string;
  reg [23:0] mul_preMul_output_rData_roundMode_string;
  reg [47:0] mul_preMul_output_rData_format_string;
  reg [23:0] mul_mul_output_payload_roundMode_string;
  reg [47:0] mul_mul_output_payload_format_string;
  reg [23:0] mul_sum1_input_payload_roundMode_string;
  reg [47:0] mul_sum1_input_payload_format_string;
  reg [23:0] mul_mul_output_rData_roundMode_string;
  reg [47:0] mul_mul_output_rData_format_string;
  reg [23:0] mul_sum1_output_payload_roundMode_string;
  reg [47:0] mul_sum1_output_payload_format_string;
  reg [23:0] mul_sum2_input_payload_roundMode_string;
  reg [47:0] mul_sum2_input_payload_format_string;
  reg [23:0] mul_sum1_output_rData_roundMode_string;
  reg [47:0] mul_sum1_output_rData_format_string;
  reg [23:0] mul_sum2_output_payload_roundMode_string;
  reg [47:0] mul_sum2_output_payload_format_string;
  reg [23:0] mul_norm_input_payload_roundMode_string;
  reg [47:0] mul_norm_input_payload_format_string;
  reg [23:0] mul_sum2_output_rData_roundMode_string;
  reg [47:0] mul_sum2_output_rData_format_string;
  reg [23:0] mul_result_output_payload_roundMode_string;
  reg [47:0] mul_result_output_payload_format_string;
  reg [23:0] mul_result_mulToAdd_payload_roundMode_string;
  reg [47:0] mul_result_mulToAdd_payload_format_string;
  reg [23:0] mul_result_mulToAdd_m2sPipe_payload_roundMode_string;
  reg [47:0] mul_result_mulToAdd_m2sPipe_payload_format_string;
  reg [23:0] mul_result_mulToAdd_rData_roundMode_string;
  reg [47:0] mul_result_mulToAdd_rData_format_string;
  reg [23:0] div_input_payload_roundMode_string;
  reg [47:0] div_input_payload_format_string;
  reg [23:0] decode_div_rData_roundMode_string;
  reg [47:0] decode_div_rData_format_string;
  reg [23:0] div_output_payload_roundMode_string;
  reg [47:0] div_output_payload_format_string;
  reg [23:0] sqrt_input_payload_roundMode_string;
  reg [47:0] sqrt_input_payload_format_string;
  reg [23:0] decode_sqrt_rData_roundMode_string;
  reg [47:0] decode_sqrt_rData_format_string;
  reg [23:0] sqrt_output_payload_roundMode_string;
  reg [47:0] sqrt_output_payload_format_string;
  reg [23:0] add_preShifter_input_payload_roundMode_string;
  reg [47:0] add_preShifter_input_payload_format_string;
  reg [23:0] add_preShifter_output_payload_roundMode_string;
  reg [47:0] add_preShifter_output_payload_format_string;
  reg [23:0] add_shifter_input_payload_roundMode_string;
  reg [47:0] add_shifter_input_payload_format_string;
  reg [23:0] add_preShifter_output_rData_roundMode_string;
  reg [47:0] add_preShifter_output_rData_format_string;
  reg [23:0] add_shifter_output_payload_roundMode_string;
  reg [47:0] add_shifter_output_payload_format_string;
  reg [23:0] add_math_input_payload_roundMode_string;
  reg [47:0] add_math_input_payload_format_string;
  reg [23:0] add_shifter_output_rData_roundMode_string;
  reg [47:0] add_shifter_output_rData_format_string;
  reg [23:0] add_math_output_payload_roundMode_string;
  reg [47:0] add_math_output_payload_format_string;
  reg [23:0] add_oh_input_payload_roundMode_string;
  reg [47:0] add_oh_input_payload_format_string;
  reg [23:0] add_math_output_rData_roundMode_string;
  reg [47:0] add_math_output_rData_format_string;
  reg [23:0] add_oh_output_payload_roundMode_string;
  reg [47:0] add_oh_output_payload_format_string;
  reg [23:0] add_norm_input_payload_roundMode_string;
  reg [47:0] add_norm_input_payload_format_string;
  reg [23:0] add_oh_output_rData_roundMode_string;
  reg [47:0] add_oh_output_rData_format_string;
  reg [23:0] add_norm_output_payload_roundMode_string;
  reg [47:0] add_norm_output_payload_format_string;
  reg [23:0] add_result_input_payload_roundMode_string;
  reg [47:0] add_result_input_payload_format_string;
  reg [23:0] add_result_output_payload_roundMode_string;
  reg [47:0] add_result_output_payload_format_string;
  reg [23:0] load_s1_output_m2sPipe_payload_roundMode_string;
  reg [47:0] load_s1_output_m2sPipe_payload_format_string;
  reg [23:0] load_s1_output_rData_roundMode_string;
  reg [47:0] load_s1_output_rData_format_string;
  reg [23:0] shortPip_output_m2sPipe_payload_roundMode_string;
  reg [47:0] shortPip_output_m2sPipe_payload_format_string;
  reg [23:0] shortPip_output_rData_roundMode_string;
  reg [47:0] shortPip_output_rData_format_string;
  reg [23:0] streamArbiter_10_io_output_combStage_payload_roundMode_string;
  reg [47:0] streamArbiter_10_io_output_combStage_payload_format_string;
  reg [23:0] merge_arbitrated_payload_roundMode_string;
  reg [47:0] merge_arbitrated_payload_format_string;
  reg [23:0] roundFront_input_payload_roundMode_string;
  reg [47:0] roundFront_input_payload_format_string;
  reg [23:0] roundFront_output_payload_roundMode_string;
  reg [47:0] roundFront_output_payload_format_string;
  reg [23:0] roundBack_input_payload_roundMode_string;
  reg [47:0] roundBack_input_payload_format_string;
  reg [47:0] roundBack_output_payload_format_string;
  reg [47:0] writeback_input_payload_format_string;
  `endif

  reg [66:0] rf_ram [0:63];
  (* ram_style = "distributed" *) reg [0:0] rf_scoreboards_0_target [0:31];
  (* ram_style = "distributed" *) reg [0:0] rf_scoreboards_0_hit [0:31];
  (* ram_style = "distributed" *) reg [0:0] rf_scoreboards_0_writes [0:31];
  (* ram_style = "distributed" *) reg [0:0] rf_scoreboards_1_target [0:31];
  (* ram_style = "distributed" *) reg [0:0] rf_scoreboards_1_hit [0:31];
  (* ram_style = "distributed" *) reg [0:0] rf_scoreboards_1_writes [0:31];

  assign _zz_commitLogic_0_pending_counter = (commitLogic_0_pending_counter + _zz_commitLogic_0_pending_counter_1);
  assign _zz_commitLogic_0_pending_counter_2 = commitLogic_0_pending_inc;
  assign _zz_commitLogic_0_pending_counter_1 = {3'd0, _zz_commitLogic_0_pending_counter_2};
  assign _zz_commitLogic_0_pending_counter_4 = commitLogic_0_pending_dec;
  assign _zz_commitLogic_0_pending_counter_3 = {3'd0, _zz_commitLogic_0_pending_counter_4};
  assign _zz_commitLogic_0_add_counter = (commitLogic_0_add_counter + _zz_commitLogic_0_add_counter_1);
  assign _zz_commitLogic_0_add_counter_2 = commitLogic_0_add_inc;
  assign _zz_commitLogic_0_add_counter_1 = {3'd0, _zz_commitLogic_0_add_counter_2};
  assign _zz_commitLogic_0_add_counter_4 = commitLogic_0_add_dec;
  assign _zz_commitLogic_0_add_counter_3 = {3'd0, _zz_commitLogic_0_add_counter_4};
  assign _zz_commitLogic_0_mul_counter = (commitLogic_0_mul_counter + _zz_commitLogic_0_mul_counter_1);
  assign _zz_commitLogic_0_mul_counter_2 = commitLogic_0_mul_inc;
  assign _zz_commitLogic_0_mul_counter_1 = {3'd0, _zz_commitLogic_0_mul_counter_2};
  assign _zz_commitLogic_0_mul_counter_4 = commitLogic_0_mul_dec;
  assign _zz_commitLogic_0_mul_counter_3 = {3'd0, _zz_commitLogic_0_mul_counter_4};
  assign _zz_commitLogic_0_div_counter = (commitLogic_0_div_counter + _zz_commitLogic_0_div_counter_1);
  assign _zz_commitLogic_0_div_counter_2 = commitLogic_0_div_inc;
  assign _zz_commitLogic_0_div_counter_1 = {3'd0, _zz_commitLogic_0_div_counter_2};
  assign _zz_commitLogic_0_div_counter_4 = commitLogic_0_div_dec;
  assign _zz_commitLogic_0_div_counter_3 = {3'd0, _zz_commitLogic_0_div_counter_4};
  assign _zz_commitLogic_0_sqrt_counter = (commitLogic_0_sqrt_counter + _zz_commitLogic_0_sqrt_counter_1);
  assign _zz_commitLogic_0_sqrt_counter_2 = commitLogic_0_sqrt_inc;
  assign _zz_commitLogic_0_sqrt_counter_1 = {3'd0, _zz_commitLogic_0_sqrt_counter_2};
  assign _zz_commitLogic_0_sqrt_counter_4 = commitLogic_0_sqrt_dec;
  assign _zz_commitLogic_0_sqrt_counter_3 = {3'd0, _zz_commitLogic_0_sqrt_counter_4};
  assign _zz_commitLogic_0_short_counter = (commitLogic_0_short_counter + _zz_commitLogic_0_short_counter_1);
  assign _zz_commitLogic_0_short_counter_2 = commitLogic_0_short_inc;
  assign _zz_commitLogic_0_short_counter_1 = {3'd0, _zz_commitLogic_0_short_counter_2};
  assign _zz_commitLogic_0_short_counter_4 = commitLogic_0_short_dec;
  assign _zz_commitLogic_0_short_counter_3 = {3'd0, _zz_commitLogic_0_short_counter_4};
  assign _zz_commitLogic_1_pending_counter = (commitLogic_1_pending_counter + _zz_commitLogic_1_pending_counter_1);
  assign _zz_commitLogic_1_pending_counter_2 = commitLogic_1_pending_inc;
  assign _zz_commitLogic_1_pending_counter_1 = {3'd0, _zz_commitLogic_1_pending_counter_2};
  assign _zz_commitLogic_1_pending_counter_4 = commitLogic_1_pending_dec;
  assign _zz_commitLogic_1_pending_counter_3 = {3'd0, _zz_commitLogic_1_pending_counter_4};
  assign _zz_commitLogic_1_add_counter = (commitLogic_1_add_counter + _zz_commitLogic_1_add_counter_1);
  assign _zz_commitLogic_1_add_counter_2 = commitLogic_1_add_inc;
  assign _zz_commitLogic_1_add_counter_1 = {3'd0, _zz_commitLogic_1_add_counter_2};
  assign _zz_commitLogic_1_add_counter_4 = commitLogic_1_add_dec;
  assign _zz_commitLogic_1_add_counter_3 = {3'd0, _zz_commitLogic_1_add_counter_4};
  assign _zz_commitLogic_1_mul_counter = (commitLogic_1_mul_counter + _zz_commitLogic_1_mul_counter_1);
  assign _zz_commitLogic_1_mul_counter_2 = commitLogic_1_mul_inc;
  assign _zz_commitLogic_1_mul_counter_1 = {3'd0, _zz_commitLogic_1_mul_counter_2};
  assign _zz_commitLogic_1_mul_counter_4 = commitLogic_1_mul_dec;
  assign _zz_commitLogic_1_mul_counter_3 = {3'd0, _zz_commitLogic_1_mul_counter_4};
  assign _zz_commitLogic_1_div_counter = (commitLogic_1_div_counter + _zz_commitLogic_1_div_counter_1);
  assign _zz_commitLogic_1_div_counter_2 = commitLogic_1_div_inc;
  assign _zz_commitLogic_1_div_counter_1 = {3'd0, _zz_commitLogic_1_div_counter_2};
  assign _zz_commitLogic_1_div_counter_4 = commitLogic_1_div_dec;
  assign _zz_commitLogic_1_div_counter_3 = {3'd0, _zz_commitLogic_1_div_counter_4};
  assign _zz_commitLogic_1_sqrt_counter = (commitLogic_1_sqrt_counter + _zz_commitLogic_1_sqrt_counter_1);
  assign _zz_commitLogic_1_sqrt_counter_2 = commitLogic_1_sqrt_inc;
  assign _zz_commitLogic_1_sqrt_counter_1 = {3'd0, _zz_commitLogic_1_sqrt_counter_2};
  assign _zz_commitLogic_1_sqrt_counter_4 = commitLogic_1_sqrt_dec;
  assign _zz_commitLogic_1_sqrt_counter_3 = {3'd0, _zz_commitLogic_1_sqrt_counter_4};
  assign _zz_commitLogic_1_short_counter = (commitLogic_1_short_counter + _zz_commitLogic_1_short_counter_1);
  assign _zz_commitLogic_1_short_counter_2 = commitLogic_1_short_inc;
  assign _zz_commitLogic_1_short_counter_1 = {3'd0, _zz_commitLogic_1_short_counter_2};
  assign _zz_commitLogic_1_short_counter_4 = commitLogic_1_short_dec;
  assign _zz_commitLogic_1_short_counter_3 = {3'd0, _zz_commitLogic_1_short_counter_4};
  assign _zz_load_s1_fsm_shift_input_1 = (load_s1_fsm_shift_input <<< 1'b1);
  assign _zz_load_s1_fsm_shift_input_2 = (load_s1_fsm_shift_input_1 <<< 2'b10);
  assign _zz_load_s1_fsm_shift_input_3 = (load_s1_fsm_shift_input_2 <<< 3'b100);
  assign _zz_load_s1_fsm_shift_input_4 = (load_s1_fsm_shift_input_3 <<< 4'b1000);
  assign _zz_load_s1_fsm_shift_input_5 = (load_s1_fsm_shift_input_4 <<< 5'h10);
  assign _zz_load_s1_fsm_shift_input_6 = (load_s1_fsm_shift_input_5 <<< 6'h20);
  assign _zz_load_s0_output_rData_value_3 = _zz_load_s0_output_rData_value_4;
  assign _zz_load_s0_output_rData_value_2 = _zz_load_s0_output_rData_value_3[31:0];
  assign _zz_load_s0_output_rData_value_4 = ({_zz_load_s0_output_rData_value_1,(_zz_load_s0_output_rData_value_1 ? (~ _zz_load_s0_output_rData_value) : _zz_load_s0_output_rData_value)} + _zz_load_s0_output_rData_value_5);
  assign _zz_load_s0_output_rData_value_6 = _zz_load_s0_output_rData_value_1;
  assign _zz_load_s0_output_rData_value_5 = {64'd0, _zz_load_s0_output_rData_value_6};
  assign _zz__zz_load_s1_fsm_shift_by_1_1 = (_zz_load_s1_fsm_shift_by - 52'h0000000000001);
  assign _zz_load_s1_recoded_exponent = (_zz_load_s1_recoded_exponent_1 + _zz_load_s1_recoded_exponent_2);
  assign _zz_load_s1_recoded_exponent_1 = ({1'b0,load_s1_passThroughFloat_exponent} - {1'b0,load_s1_fsm_expOffset});
  assign _zz_load_s1_recoded_exponent_2 = {1'd0, load_s1_recodedExpOffset};
  assign _zz_load_s1_output_payload_value_exponent = {6'd0, load_s1_fsm_shift_by};
  assign _zz_shortPip_f32_exp = (shortPip_input_payload_rs1_exponent - 12'h780);
  assign _zz_shortPip_f64_exp = (shortPip_input_payload_rs1_exponent - 12'h400);
  assign _zz_shortPip_expInSubnormalRange = {1'd0, shortPip_expSubnormalThreshold};
  assign _zz_shortPip_fsm_shift_input_1 = (shortPip_fsm_shift_input >>> 6'h20);
  assign _zz_shortPip_fsm_shift_input_2 = (shortPip_fsm_shift_input_1 >>> 5'h10);
  assign _zz_shortPip_fsm_shift_input_3 = (shortPip_fsm_shift_input_2 >>> 4'b1000);
  assign _zz_shortPip_fsm_shift_input_4 = (shortPip_fsm_shift_input_3 >>> 3'b100);
  assign _zz_shortPip_fsm_shift_input_5 = (shortPip_fsm_shift_input_4 >>> 2'b10);
  assign _zz_shortPip_fsm_shift_input_6 = (shortPip_fsm_shift_input_5 >>> 1'b1);
  assign _zz_shortPip_fsm_shift_by_2 = (((_zz_shortPip_fsm_shift_by < _zz_shortPip_fsm_shift_by_3) ? _zz_shortPip_fsm_shift_by : _zz_shortPip_fsm_shift_by_4) + 12'h014);
  assign _zz_shortPip_fsm_shift_by_3 = {6'd0, _zz_shortPip_fsm_shift_by_1};
  assign _zz_shortPip_fsm_shift_by_4 = {6'd0, _zz_shortPip_fsm_shift_by_1};
  assign _zz_shortPip_fsm_shift_by_5 = (_zz_shortPip_fsm_shift_by_6 - shortPip_input_payload_rs1_exponent);
  assign _zz_shortPip_fsm_shift_by_6 = {1'd0, shortPip_fsm_formatShiftOffset};
  assign _zz_shortPip_f2i_result_1 = (shortPip_f2i_resign ^ shortPip_f2i_increment);
  assign _zz_shortPip_f2i_result = {31'd0, _zz_shortPip_f2i_result_1};
  assign _zz_mul_sum1_sum = (_zz_mul_sum1_sum_1 + _zz_mul_sum1_sum_2);
  assign _zz_mul_sum1_sum_1 = {70'd0, mul_sum1_input_payload_muls_0};
  assign _zz_mul_sum1_sum_3 = ({18'd0,mul_sum1_input_payload_muls_1} <<< 5'd18);
  assign _zz_mul_sum1_sum_2 = {52'd0, _zz_mul_sum1_sum_3};
  assign _zz_mul_sum1_sum_4 = (_zz_mul_sum1_sum_5 + _zz_mul_sum1_sum_7);
  assign _zz_mul_sum1_sum_6 = ({18'd0,mul_sum1_input_payload_muls_2} <<< 5'd18);
  assign _zz_mul_sum1_sum_5 = {52'd0, _zz_mul_sum1_sum_6};
  assign _zz_mul_sum1_sum_8 = ({36'd0,mul_sum1_input_payload_muls_3} <<< 6'd36);
  assign _zz_mul_sum1_sum_7 = {35'd0, _zz_mul_sum1_sum_8};
  assign _zz_mul_sum2_sum = (_zz_mul_sum2_sum_1 + _zz_mul_sum2_sum_12);
  assign _zz_mul_sum2_sum_1 = (_zz_mul_sum2_sum_2 + _zz_mul_sum2_sum_7);
  assign _zz_mul_sum2_sum_2 = (_zz_mul_sum2_sum_3 + _zz_mul_sum2_sum_5);
  assign _zz_mul_sum2_sum_4 = ({36'd0,mul_sum2_input_payload_muls2_0} <<< 6'd36);
  assign _zz_mul_sum2_sum_3 = {35'd0, _zz_mul_sum2_sum_4};
  assign _zz_mul_sum2_sum_6 = ({36'd0,mul_sum2_input_payload_muls2_1} <<< 6'd36);
  assign _zz_mul_sum2_sum_5 = {34'd0, _zz_mul_sum2_sum_6};
  assign _zz_mul_sum2_sum_7 = (_zz_mul_sum2_sum_8 + _zz_mul_sum2_sum_10);
  assign _zz_mul_sum2_sum_9 = ({54'd0,mul_sum2_input_payload_muls2_2} <<< 6'd54);
  assign _zz_mul_sum2_sum_8 = {17'd0, _zz_mul_sum2_sum_9};
  assign _zz_mul_sum2_sum_11 = ({54'd0,mul_sum2_input_payload_muls2_3} <<< 6'd54);
  assign _zz_mul_sum2_sum_10 = {17'd0, _zz_mul_sum2_sum_11};
  assign _zz_mul_sum2_sum_12 = ({72'd0,mul_sum2_input_payload_muls2_4} <<< 7'd72);
  assign _zz_mul_norm_exp_1 = mul_norm_needShift;
  assign _zz_mul_norm_exp = {12'd0, _zz_mul_norm_exp_1};
  assign _zz_mul_norm_forceUnderflow = {1'd0, mul_norm_underflowThreshold};
  assign _zz_mul_norm_output_exponent = (mul_norm_exp - 13'h07ff);
  assign _zz_div_exponent = (_zz_div_exponent_1 - _zz_div_exponent_3);
  assign _zz_div_exponent_1 = (_zz_div_exponent_2 + 14'h27ff);
  assign _zz_div_exponent_2 = {2'd0, div_input_payload_rs1_exponent};
  assign _zz_div_exponent_3 = {2'd0, div_input_payload_rs2_exponent};
  assign _zz_div_exponent_5 = div_needShift;
  assign _zz_div_exponent_4 = {13'd0, _zz_div_exponent_5};
  assign _zz_sqrt_exponent = (_zz_sqrt_exponent_1 + {1'b0,_zz_sqrt_exponent_3});
  assign _zz_sqrt_exponent_2 = {1'b0,10'h3ff};
  assign _zz_sqrt_exponent_1 = {1'd0, _zz_sqrt_exponent_2};
  assign _zz_sqrt_exponent_3 = (sqrt_input_payload_rs1_exponent >>> 1'd1);
  assign _zz_sqrt_exponent_5 = sqrt_input_payload_rs1_exponent[0];
  assign _zz_sqrt_exponent_4 = {11'd0, _zz_sqrt_exponent_5};
  assign _zz_add_shifter_shiftBy_1 = (_zz_add_shifter_shiftBy[12] ? _zz_add_shifter_shiftBy_2 : _zz_add_shifter_shiftBy);
  assign _zz_add_shifter_shiftBy_2 = (~ _zz_add_shifter_shiftBy);
  assign _zz_add_shifter_shiftBy_4 = _zz_add_shifter_shiftBy[12];
  assign _zz_add_shifter_shiftBy_3 = {12'd0, _zz_add_shifter_shiftBy_4};
  assign _zz_add_shifter_yMantissa_1 = (add_shifter_yMantissa >>> 6'h20);
  assign _zz_add_shifter_yMantissa_2 = (add_shifter_yMantissa_1 >>> 5'h10);
  assign _zz_add_shifter_yMantissa_3 = (add_shifter_yMantissa_2 >>> 4'b1000);
  assign _zz_add_shifter_yMantissa_4 = (add_shifter_yMantissa_3 >>> 3'b100);
  assign _zz_add_shifter_yMantissa_5 = (add_shifter_yMantissa_4 >>> 2'b10);
  assign _zz_add_shifter_yMantissa_6 = (add_shifter_yMantissa_5 >>> 1'b1);
  assign _zz_add_math_xSigned = ({add_math_input_payload_xSign,(add_math_input_payload_xSign ? (~ add_math_input_payload_xMantissa) : add_math_input_payload_xMantissa)} + _zz_add_math_xSigned_1);
  assign _zz_add_math_xSigned_2 = add_math_input_payload_xSign;
  assign _zz_add_math_xSigned_1 = {55'd0, _zz_add_math_xSigned_2};
  assign _zz_add_math_ySigned = ({add_math_input_payload_ySign,(add_math_input_payload_ySign ? (~ add_math_input_payload_yMantissa) : add_math_input_payload_yMantissa)} + _zz_add_math_ySigned_1);
  assign _zz_add_math_ySigned_2 = (add_math_input_payload_ySign && (! add_math_input_payload_roundingScrap));
  assign _zz_add_math_ySigned_1 = {55'd0, _zz_add_math_ySigned_2};
  assign _zz_add_math_output_payload_xyMantissa = _zz_add_math_output_payload_xyMantissa_1;
  assign _zz_add_math_output_payload_xyMantissa_1 = ($signed(_zz_add_math_output_payload_xyMantissa_2) + $signed(_zz_add_math_output_payload_xyMantissa_3));
  assign _zz_add_math_output_payload_xyMantissa_2 = {add_math_xSigned[55],add_math_xSigned};
  assign _zz_add_math_output_payload_xyMantissa_3 = {add_math_ySigned[55],add_math_ySigned};
  assign _zz__zz_add_oh_shift_1_1 = (_zz_add_oh_shift - 56'h00000000000001);
  assign _zz_add_norm_output_payload_exponent = ({1'b0,add_norm_input_payload_xyExponent} - _zz_add_norm_output_payload_exponent_1);
  assign _zz_add_norm_output_payload_exponent_2 = {1'b0,add_norm_input_payload_shift};
  assign _zz_add_norm_output_payload_exponent_1 = {6'd0, _zz_add_norm_output_payload_exponent_2};
  assign _zz_add_result_output_payload_value_mantissa = (add_result_input_payload_mantissa >>> 2'd2);
  assign _zz_roundFront_expDif_1 = {1'b0,roundFront_expBase};
  assign _zz_roundFront_expDif = {1'd0, _zz_roundFront_expDif_1};
  assign _zz_roundFront_roundAdjusted = {1'b1,_zz_roundFront_roundAdjusted_1};
  assign _zz_roundFront_roundAdjusted_1 = (roundFront_manAggregate >>> 1'd1);
  assign _zz_roundFront_rneBit = {2'b01,_zz_roundFront_rneBit_1};
  assign _zz_roundFront_rneBit_1 = (roundFront_manAggregate >>> 2'd2);
  assign _zz_roundBack_adderMantissa = (roundBack_input_payload_exactMask[52 : 0] >>> 1'd1);
  assign _zz_roundBack_adderRightOp = (roundBack_input_payload_mantissaIncrement ? _zz_roundBack_adderRightOp_1 : 53'h0);
  assign _zz_roundBack_adderRightOp_1 = (roundBack_input_payload_exactMask >>> 1'd1);
  assign _zz_roundBack_adder_2 = (_zz_roundBack_adder + _zz_roundBack_adder_3);
  assign _zz_roundBack_adder_3 = {12'd0, roundBack_adderRightOp};
  assign _zz_roundBack_adder_4 = {63'd0, _zz_roundBack_adder_1};
  assign _zz_roundBack_masked_1 = _zz_roundBack_masked_2[51:0];
  assign _zz_roundBack_masked = {12'd0, _zz_roundBack_masked_1};
  assign _zz_roundBack_masked_2 = (roundBack_input_payload_exactMask >>> 1'd1);
  assign _zz_roundBack_borringCase = {1'd0, roundBack_ufSubnormalThreshold};
  assign _zz_when_FpuCore_l1616 = {1'd0, roundBack_ufSubnormalThreshold};
  assign _zz_when_FpuCore_l1638 = {1'd0, roundBack_ufThreshold};
  assign _zz_rf_ram_port = {writeback_port_payload_data_boxed,{writeback_port_payload_data_value_special,{writeback_port_payload_data_value_sign,{writeback_port_payload_data_value_exponent,writeback_port_payload_data_value_mantissa}}}};
  assign _zz_rf_scoreboards_0_target_port = rf_scoreboards_0_targetWrite_payload_data;
  assign _zz_rf_scoreboards_0_hit_port = rf_scoreboards_0_hitWrite_payload_data;
  assign _zz_rf_scoreboards_0_writes_port = commitLogic_0_input_payload_write;
  assign _zz_rf_scoreboards_1_target_port = rf_scoreboards_1_targetWrite_payload_data;
  assign _zz_rf_scoreboards_1_hit_port = rf_scoreboards_1_hitWrite_payload_data;
  assign _zz_rf_scoreboards_1_writes_port = commitLogic_1_input_payload_write;
  assign _zz_decode_shortPipHit = FpuOpcode_MIN_MAX;
  assign _zz_decode_shortPipHit_1 = (decode_input_payload_opcode == FpuOpcode_CMP);
  assign _zz_decode_shortPipHit_2 = (decode_input_payload_opcode == FpuOpcode_F2I);
  assign _zz_decode_shortPipHit_3 = (decode_input_payload_opcode == FpuOpcode_STORE);
  assign _zz__zz_load_s1_fsm_shift_by = load_s1_fsm_ohInput[7];
  assign _zz__zz_load_s1_fsm_shift_by_1 = load_s1_fsm_ohInput[8];
  assign _zz__zz_load_s1_fsm_shift_by_2 = {load_s1_fsm_ohInput[9],{load_s1_fsm_ohInput[10],{load_s1_fsm_ohInput[11],{load_s1_fsm_ohInput[12],{load_s1_fsm_ohInput[13],{load_s1_fsm_ohInput[14],{load_s1_fsm_ohInput[15],{load_s1_fsm_ohInput[16],{load_s1_fsm_ohInput[17],{_zz__zz_load_s1_fsm_shift_by_3,{_zz__zz_load_s1_fsm_shift_by_4,_zz__zz_load_s1_fsm_shift_by_5}}}}}}}}}}};
  assign _zz__zz_load_s1_fsm_shift_by_3 = load_s1_fsm_ohInput[18];
  assign _zz__zz_load_s1_fsm_shift_by_4 = load_s1_fsm_ohInput[19];
  assign _zz__zz_load_s1_fsm_shift_by_5 = {load_s1_fsm_ohInput[20],{load_s1_fsm_ohInput[21],{load_s1_fsm_ohInput[22],{load_s1_fsm_ohInput[23],{load_s1_fsm_ohInput[24],{load_s1_fsm_ohInput[25],{load_s1_fsm_ohInput[26],{load_s1_fsm_ohInput[27],{load_s1_fsm_ohInput[28],{_zz__zz_load_s1_fsm_shift_by_6,{_zz__zz_load_s1_fsm_shift_by_7,_zz__zz_load_s1_fsm_shift_by_8}}}}}}}}}}};
  assign _zz__zz_load_s1_fsm_shift_by_6 = load_s1_fsm_ohInput[29];
  assign _zz__zz_load_s1_fsm_shift_by_7 = load_s1_fsm_ohInput[30];
  assign _zz__zz_load_s1_fsm_shift_by_8 = {load_s1_fsm_ohInput[31],{load_s1_fsm_ohInput[32],{load_s1_fsm_ohInput[33],{load_s1_fsm_ohInput[34],{load_s1_fsm_ohInput[35],{load_s1_fsm_ohInput[36],{load_s1_fsm_ohInput[37],{load_s1_fsm_ohInput[38],{load_s1_fsm_ohInput[39],{_zz__zz_load_s1_fsm_shift_by_9,{_zz__zz_load_s1_fsm_shift_by_10,_zz__zz_load_s1_fsm_shift_by_11}}}}}}}}}}};
  assign _zz__zz_load_s1_fsm_shift_by_9 = load_s1_fsm_ohInput[40];
  assign _zz__zz_load_s1_fsm_shift_by_10 = load_s1_fsm_ohInput[41];
  assign _zz__zz_load_s1_fsm_shift_by_11 = {load_s1_fsm_ohInput[42],{load_s1_fsm_ohInput[43],{load_s1_fsm_ohInput[44],{load_s1_fsm_ohInput[45],{load_s1_fsm_ohInput[46],{load_s1_fsm_ohInput[47],{load_s1_fsm_ohInput[48],{load_s1_fsm_ohInput[49],{load_s1_fsm_ohInput[50],load_s1_fsm_ohInput[51]}}}}}}}}};
  assign _zz__zz_load_s1_fsm_shift_by_47 = (((((((((_zz_load_s1_fsm_shift_by_1[1] || _zz_load_s1_fsm_shift_by_2) || _zz_load_s1_fsm_shift_by_3) || _zz_load_s1_fsm_shift_by_5) || _zz_load_s1_fsm_shift_by_6) || _zz_load_s1_fsm_shift_by_8) || _zz_load_s1_fsm_shift_by_10) || _zz_load_s1_fsm_shift_by_12) || _zz_load_s1_fsm_shift_by_13) || _zz_load_s1_fsm_shift_by_15);
  assign _zz__zz_load_s1_fsm_shift_by_48 = (((((((((_zz_load_s1_fsm_shift_by_1[2] || _zz_load_s1_fsm_shift_by_2) || _zz_load_s1_fsm_shift_by_4) || _zz_load_s1_fsm_shift_by_5) || _zz_load_s1_fsm_shift_by_7) || _zz_load_s1_fsm_shift_by_8) || _zz_load_s1_fsm_shift_by_11) || _zz_load_s1_fsm_shift_by_12) || _zz_load_s1_fsm_shift_by_14) || _zz_load_s1_fsm_shift_by_15);
  assign _zz__zz_load_s1_fsm_shift_by_49 = ((((((_zz_load_s1_fsm_shift_by_1[4] || _zz_load_s1_fsm_shift_by_3) || _zz_load_s1_fsm_shift_by_4) || _zz_load_s1_fsm_shift_by_5) || _zz_load_s1_fsm_shift_by_9) || _zz_load_s1_fsm_shift_by_10) || _zz_load_s1_fsm_shift_by_11);
  assign _zz__zz_load_s1_fsm_shift_by_50 = (((((((_zz_load_s1_fsm_shift_by_1[8] || _zz_load_s1_fsm_shift_by_6) || _zz_load_s1_fsm_shift_by_7) || _zz_load_s1_fsm_shift_by_8) || _zz_load_s1_fsm_shift_by_9) || _zz_load_s1_fsm_shift_by_10) || _zz_load_s1_fsm_shift_by_11) || _zz_load_s1_fsm_shift_by_12);
  assign _zz__zz_load_s1_fsm_shift_by_51 = ((_zz_load_s1_fsm_shift_by_1[16] || _zz_load_s1_fsm_shift_by_13) || _zz_load_s1_fsm_shift_by_14);
  assign _zz__zz_load_s1_fsm_shift_by_52 = (((_zz_load_s1_fsm_shift_by_1[32] || _zz_load_s1_fsm_shift_by_28) || _zz_load_s1_fsm_shift_by_29) || _zz_load_s1_fsm_shift_by_30);
  assign _zz_shortPip_f2i_underflow = shortPip_f2i_unsigned[30 : 0];
  assign _zz_shortPip_f2i_underflow_1 = 31'h0;
  assign _zz__zz_add_oh_shift = add_oh_output_payload_xyMantissa[7];
  assign _zz__zz_add_oh_shift_1 = add_oh_output_payload_xyMantissa[8];
  assign _zz__zz_add_oh_shift_2 = {add_oh_output_payload_xyMantissa[9],{add_oh_output_payload_xyMantissa[10],{add_oh_output_payload_xyMantissa[11],{add_oh_output_payload_xyMantissa[12],{add_oh_output_payload_xyMantissa[13],{add_oh_output_payload_xyMantissa[14],{add_oh_output_payload_xyMantissa[15],{add_oh_output_payload_xyMantissa[16],{add_oh_output_payload_xyMantissa[17],{_zz__zz_add_oh_shift_3,{_zz__zz_add_oh_shift_4,_zz__zz_add_oh_shift_5}}}}}}}}}}};
  assign _zz__zz_add_oh_shift_3 = add_oh_output_payload_xyMantissa[18];
  assign _zz__zz_add_oh_shift_4 = add_oh_output_payload_xyMantissa[19];
  assign _zz__zz_add_oh_shift_5 = {add_oh_output_payload_xyMantissa[20],{add_oh_output_payload_xyMantissa[21],{add_oh_output_payload_xyMantissa[22],{add_oh_output_payload_xyMantissa[23],{add_oh_output_payload_xyMantissa[24],{add_oh_output_payload_xyMantissa[25],{add_oh_output_payload_xyMantissa[26],{add_oh_output_payload_xyMantissa[27],{add_oh_output_payload_xyMantissa[28],{_zz__zz_add_oh_shift_6,{_zz__zz_add_oh_shift_7,_zz__zz_add_oh_shift_8}}}}}}}}}}};
  assign _zz__zz_add_oh_shift_6 = add_oh_output_payload_xyMantissa[29];
  assign _zz__zz_add_oh_shift_7 = add_oh_output_payload_xyMantissa[30];
  assign _zz__zz_add_oh_shift_8 = {add_oh_output_payload_xyMantissa[31],{add_oh_output_payload_xyMantissa[32],{add_oh_output_payload_xyMantissa[33],{add_oh_output_payload_xyMantissa[34],{add_oh_output_payload_xyMantissa[35],{add_oh_output_payload_xyMantissa[36],{add_oh_output_payload_xyMantissa[37],{add_oh_output_payload_xyMantissa[38],{add_oh_output_payload_xyMantissa[39],{_zz__zz_add_oh_shift_9,{_zz__zz_add_oh_shift_10,_zz__zz_add_oh_shift_11}}}}}}}}}}};
  assign _zz__zz_add_oh_shift_9 = add_oh_output_payload_xyMantissa[40];
  assign _zz__zz_add_oh_shift_10 = add_oh_output_payload_xyMantissa[41];
  assign _zz__zz_add_oh_shift_11 = {add_oh_output_payload_xyMantissa[42],{add_oh_output_payload_xyMantissa[43],{add_oh_output_payload_xyMantissa[44],{add_oh_output_payload_xyMantissa[45],{add_oh_output_payload_xyMantissa[46],{add_oh_output_payload_xyMantissa[47],{add_oh_output_payload_xyMantissa[48],{add_oh_output_payload_xyMantissa[49],{add_oh_output_payload_xyMantissa[50],{_zz__zz_add_oh_shift_12,{_zz__zz_add_oh_shift_13,_zz__zz_add_oh_shift_14}}}}}}}}}}};
  assign _zz__zz_add_oh_shift_12 = add_oh_output_payload_xyMantissa[51];
  assign _zz__zz_add_oh_shift_13 = add_oh_output_payload_xyMantissa[52];
  assign _zz__zz_add_oh_shift_14 = {add_oh_output_payload_xyMantissa[53],{add_oh_output_payload_xyMantissa[54],add_oh_output_payload_xyMantissa[55]}};
  assign _zz__zz_add_oh_shift_51 = (((((((((((_zz_add_oh_shift_1[1] || _zz_add_oh_shift_2) || _zz_add_oh_shift_3) || _zz_add_oh_shift_5) || _zz_add_oh_shift_6) || _zz_add_oh_shift_8) || _zz_add_oh_shift_10) || _zz_add_oh_shift_12) || _zz_add_oh_shift_13) || _zz_add_oh_shift_15) || _zz_add_oh_shift_17) || _zz_add_oh_shift_19);
  assign _zz__zz_add_oh_shift_52 = (((((((((((_zz_add_oh_shift_1[2] || _zz_add_oh_shift_2) || _zz_add_oh_shift_4) || _zz_add_oh_shift_5) || _zz_add_oh_shift_7) || _zz_add_oh_shift_8) || _zz_add_oh_shift_11) || _zz_add_oh_shift_12) || _zz_add_oh_shift_14) || _zz_add_oh_shift_15) || _zz_add_oh_shift_18) || _zz_add_oh_shift_19);
  assign _zz__zz_add_oh_shift_53 = (((((((((((_zz_add_oh_shift_1[4] || _zz_add_oh_shift_3) || _zz_add_oh_shift_4) || _zz_add_oh_shift_5) || _zz_add_oh_shift_9) || _zz_add_oh_shift_10) || _zz_add_oh_shift_11) || _zz_add_oh_shift_12) || _zz_add_oh_shift_16) || _zz_add_oh_shift_17) || _zz_add_oh_shift_18) || _zz_add_oh_shift_19);
  assign _zz__zz_add_oh_shift_54 = ((((((_zz_add_oh_shift_1[8] || _zz_add_oh_shift_6) || _zz_add_oh_shift_7) || _zz_add_oh_shift_8) || _zz_add_oh_shift_9) || _zz_add_oh_shift_10) || _zz_add_oh_shift_11);
  assign _zz__zz_add_oh_shift_55 = ((((((_zz_add_oh_shift_1[16] || _zz_add_oh_shift_13) || _zz_add_oh_shift_14) || _zz_add_oh_shift_15) || _zz_add_oh_shift_16) || _zz_add_oh_shift_17) || _zz_add_oh_shift_18);
  assign _zz__zz_add_oh_shift_56 = (((((((_zz_add_oh_shift_1[32] || _zz_add_oh_shift_28) || _zz_add_oh_shift_29) || _zz_add_oh_shift_30) || _zz_add_oh_shift_31) || _zz_add_oh_shift_32) || _zz_add_oh_shift_33) || _zz_add_oh_shift_34);
  assign _zz_roundFront_exactMask = 6'h30;
  assign _zz_roundFront_exactMask_1 = (6'h2f < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_2 = (6'h2e < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_3 = {(6'h2d < roundFront_discardCountTrunk),{(6'h2c < roundFront_discardCountTrunk),{(6'h2b < roundFront_discardCountTrunk),{(6'h2a < roundFront_discardCountTrunk),{(6'h29 < roundFront_discardCountTrunk),{(_zz_roundFront_exactMask_4 < roundFront_discardCountTrunk),{_zz_roundFront_exactMask_5,{_zz_roundFront_exactMask_6,_zz_roundFront_exactMask_7}}}}}}}};
  assign _zz_roundFront_exactMask_4 = 6'h28;
  assign _zz_roundFront_exactMask_5 = (6'h27 < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_6 = (6'h26 < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_7 = {(6'h25 < roundFront_discardCountTrunk),{(6'h24 < roundFront_discardCountTrunk),{(6'h23 < roundFront_discardCountTrunk),{(6'h22 < roundFront_discardCountTrunk),{(6'h21 < roundFront_discardCountTrunk),{(_zz_roundFront_exactMask_8 < roundFront_discardCountTrunk),{_zz_roundFront_exactMask_9,{_zz_roundFront_exactMask_10,_zz_roundFront_exactMask_11}}}}}}}};
  assign _zz_roundFront_exactMask_8 = 6'h20;
  assign _zz_roundFront_exactMask_9 = (6'h1f < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_10 = (6'h1e < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_11 = {(6'h1d < roundFront_discardCountTrunk),{(6'h1c < roundFront_discardCountTrunk),{(6'h1b < roundFront_discardCountTrunk),{(6'h1a < roundFront_discardCountTrunk),{(6'h19 < roundFront_discardCountTrunk),{(_zz_roundFront_exactMask_12 < roundFront_discardCountTrunk),{_zz_roundFront_exactMask_13,{_zz_roundFront_exactMask_14,_zz_roundFront_exactMask_15}}}}}}}};
  assign _zz_roundFront_exactMask_12 = 6'h18;
  assign _zz_roundFront_exactMask_13 = (6'h17 < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_14 = (6'h16 < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_15 = {(6'h15 < roundFront_discardCountTrunk),{(6'h14 < roundFront_discardCountTrunk),{(6'h13 < roundFront_discardCountTrunk),{(6'h12 < roundFront_discardCountTrunk),{(6'h11 < roundFront_discardCountTrunk),{(_zz_roundFront_exactMask_16 < roundFront_discardCountTrunk),{_zz_roundFront_exactMask_17,{_zz_roundFront_exactMask_18,_zz_roundFront_exactMask_19}}}}}}}};
  assign _zz_roundFront_exactMask_16 = 6'h10;
  assign _zz_roundFront_exactMask_17 = (6'h0f < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_18 = (6'h0e < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_19 = {(6'h0d < roundFront_discardCountTrunk),{(6'h0c < roundFront_discardCountTrunk),{(6'h0b < roundFront_discardCountTrunk),{(6'h0a < roundFront_discardCountTrunk),{(6'h09 < roundFront_discardCountTrunk),{(_zz_roundFront_exactMask_20 < roundFront_discardCountTrunk),{_zz_roundFront_exactMask_21,{_zz_roundFront_exactMask_22,_zz_roundFront_exactMask_23}}}}}}}};
  assign _zz_roundFront_exactMask_20 = 6'h08;
  assign _zz_roundFront_exactMask_21 = (6'h07 < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_22 = (6'h06 < roundFront_discardCountTrunk);
  assign _zz_roundFront_exactMask_23 = {(6'h05 < roundFront_discardCountTrunk),{(6'h04 < roundFront_discardCountTrunk),{(6'h03 < roundFront_discardCountTrunk),{(6'h02 < roundFront_discardCountTrunk),{(6'h01 < roundFront_discardCountTrunk),{(6'h0 < roundFront_discardCountTrunk),1'b1}}}}}};
  always @(posedge io_systemClk) begin
    if(_zz_read_rs_0_boxed_1) begin
      rf_ram_spinal_port0 <= rf_ram[_zz_read_rs_0_boxed];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_read_rs_1_boxed_1) begin
      rf_ram_spinal_port1 <= rf_ram[_zz_read_rs_1_boxed];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_read_rs_2_boxed_1) begin
      rf_ram_spinal_port2 <= rf_ram[_zz_read_rs_2_boxed];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      rf_ram[writeback_port_payload_address] <= _zz_rf_ram_port;
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_7) begin
      rf_scoreboards_0_target[rf_scoreboards_0_targetWrite_payload_address] <= _zz_rf_scoreboards_0_target_port;
    end
  end

  assign rf_scoreboards_0_target_spinal_port1 = rf_scoreboards_0_target[scheduler_0_input_payload_rs1];
  assign rf_scoreboards_0_target_spinal_port2 = rf_scoreboards_0_target[scheduler_0_input_payload_rs2];
  assign rf_scoreboards_0_target_spinal_port3 = rf_scoreboards_0_target[scheduler_0_input_payload_rs3];
  assign rf_scoreboards_0_target_spinal_port4 = rf_scoreboards_0_target[scheduler_0_input_payload_rd];
  always @(posedge io_systemClk) begin
    if(_zz_6) begin
      rf_scoreboards_0_hit[rf_scoreboards_0_hitWrite_payload_address] <= _zz_rf_scoreboards_0_hit_port;
    end
  end

  assign rf_scoreboards_0_hit_spinal_port1 = rf_scoreboards_0_hit[scheduler_0_input_payload_rs1];
  assign rf_scoreboards_0_hit_spinal_port2 = rf_scoreboards_0_hit[scheduler_0_input_payload_rs2];
  assign rf_scoreboards_0_hit_spinal_port3 = rf_scoreboards_0_hit[scheduler_0_input_payload_rs3];
  assign rf_scoreboards_0_hit_spinal_port4 = rf_scoreboards_0_hit[scheduler_0_input_payload_rd];
  assign rf_scoreboards_0_hit_spinal_port5 = rf_scoreboards_0_hit[writeback_input_payload_rd];
  always @(posedge io_systemClk) begin
    if(_zz_3) begin
      rf_scoreboards_0_writes[commitLogic_0_input_payload_rd] <= _zz_rf_scoreboards_0_writes_port;
    end
  end

  assign rf_scoreboards_0_writes_spinal_port1 = rf_scoreboards_0_writes[roundBack_input_payload_rd];
  always @(posedge io_systemClk) begin
    if(_zz_5) begin
      rf_scoreboards_1_target[rf_scoreboards_1_targetWrite_payload_address] <= _zz_rf_scoreboards_1_target_port;
    end
  end

  assign rf_scoreboards_1_target_spinal_port1 = rf_scoreboards_1_target[scheduler_1_input_payload_rs1];
  assign rf_scoreboards_1_target_spinal_port2 = rf_scoreboards_1_target[scheduler_1_input_payload_rs2];
  assign rf_scoreboards_1_target_spinal_port3 = rf_scoreboards_1_target[scheduler_1_input_payload_rs3];
  assign rf_scoreboards_1_target_spinal_port4 = rf_scoreboards_1_target[scheduler_1_input_payload_rd];
  always @(posedge io_systemClk) begin
    if(_zz_4) begin
      rf_scoreboards_1_hit[rf_scoreboards_1_hitWrite_payload_address] <= _zz_rf_scoreboards_1_hit_port;
    end
  end

  assign rf_scoreboards_1_hit_spinal_port1 = rf_scoreboards_1_hit[scheduler_1_input_payload_rs1];
  assign rf_scoreboards_1_hit_spinal_port2 = rf_scoreboards_1_hit[scheduler_1_input_payload_rs2];
  assign rf_scoreboards_1_hit_spinal_port3 = rf_scoreboards_1_hit[scheduler_1_input_payload_rs3];
  assign rf_scoreboards_1_hit_spinal_port4 = rf_scoreboards_1_hit[scheduler_1_input_payload_rd];
  assign rf_scoreboards_1_hit_spinal_port5 = rf_scoreboards_1_hit[writeback_input_payload_rd];
  always @(posedge io_systemClk) begin
    if(_zz_2) begin
      rf_scoreboards_1_writes[commitLogic_1_input_payload_rd] <= _zz_rf_scoreboards_1_writes_port;
    end
  end

  assign rf_scoreboards_1_writes_spinal_port1 = rf_scoreboards_1_writes[roundBack_input_payload_rd];
  StreamFork streamFork_3 (
    .io_input_valid              (io_port_0_commit_valid                       ), //i
    .io_input_ready              (streamFork_3_io_input_ready                  ), //o
    .io_input_payload_opcode     (io_port_0_commit_payload_opcode[3:0]         ), //i
    .io_input_payload_rd         (io_port_0_commit_payload_rd[4:0]             ), //i
    .io_input_payload_write      (io_port_0_commit_payload_write               ), //i
    .io_input_payload_value      (io_port_0_commit_payload_value[63:0]         ), //i
    .io_outputs_0_valid          (streamFork_3_io_outputs_0_valid              ), //o
    .io_outputs_0_ready          (commitFork_load_0_ready                      ), //i
    .io_outputs_0_payload_opcode (streamFork_3_io_outputs_0_payload_opcode[3:0]), //o
    .io_outputs_0_payload_rd     (streamFork_3_io_outputs_0_payload_rd[4:0]    ), //o
    .io_outputs_0_payload_write  (streamFork_3_io_outputs_0_payload_write      ), //o
    .io_outputs_0_payload_value  (streamFork_3_io_outputs_0_payload_value[63:0]), //o
    .io_outputs_1_valid          (streamFork_3_io_outputs_1_valid              ), //o
    .io_outputs_1_ready          (streamFork_3_io_outputs_1_rValidN            ), //i
    .io_outputs_1_payload_opcode (streamFork_3_io_outputs_1_payload_opcode[3:0]), //o
    .io_outputs_1_payload_rd     (streamFork_3_io_outputs_1_payload_rd[4:0]    ), //o
    .io_outputs_1_payload_write  (streamFork_3_io_outputs_1_payload_write      ), //o
    .io_outputs_1_payload_value  (streamFork_3_io_outputs_1_payload_value[63:0])  //o
  );
  StreamFork streamFork_4 (
    .io_input_valid              (io_port_1_commit_valid                       ), //i
    .io_input_ready              (streamFork_4_io_input_ready                  ), //o
    .io_input_payload_opcode     (io_port_1_commit_payload_opcode[3:0]         ), //i
    .io_input_payload_rd         (io_port_1_commit_payload_rd[4:0]             ), //i
    .io_input_payload_write      (io_port_1_commit_payload_write               ), //i
    .io_input_payload_value      (io_port_1_commit_payload_value[63:0]         ), //i
    .io_outputs_0_valid          (streamFork_4_io_outputs_0_valid              ), //o
    .io_outputs_0_ready          (commitFork_load_1_ready                      ), //i
    .io_outputs_0_payload_opcode (streamFork_4_io_outputs_0_payload_opcode[3:0]), //o
    .io_outputs_0_payload_rd     (streamFork_4_io_outputs_0_payload_rd[4:0]    ), //o
    .io_outputs_0_payload_write  (streamFork_4_io_outputs_0_payload_write      ), //o
    .io_outputs_0_payload_value  (streamFork_4_io_outputs_0_payload_value[63:0]), //o
    .io_outputs_1_valid          (streamFork_4_io_outputs_1_valid              ), //o
    .io_outputs_1_ready          (streamFork_4_io_outputs_1_rValidN            ), //i
    .io_outputs_1_payload_opcode (streamFork_4_io_outputs_1_payload_opcode[3:0]), //o
    .io_outputs_1_payload_rd     (streamFork_4_io_outputs_1_payload_rd[4:0]    ), //o
    .io_outputs_1_payload_write  (streamFork_4_io_outputs_1_payload_write      ), //o
    .io_outputs_1_payload_value  (streamFork_4_io_outputs_1_payload_value[63:0])  //o
  );
  StreamArbiter cmdArbiter_arbiter (
    .io_inputs_0_valid             (scheduler_0_output_m2sPipe_valid                   ), //i
    .io_inputs_0_ready             (cmdArbiter_arbiter_io_inputs_0_ready               ), //o
    .io_inputs_0_payload_opcode    (scheduler_0_output_m2sPipe_payload_opcode[3:0]     ), //i
    .io_inputs_0_payload_arg       (scheduler_0_output_m2sPipe_payload_arg[1:0]        ), //i
    .io_inputs_0_payload_rs1       (scheduler_0_output_m2sPipe_payload_rs1[4:0]        ), //i
    .io_inputs_0_payload_rs2       (scheduler_0_output_m2sPipe_payload_rs2[4:0]        ), //i
    .io_inputs_0_payload_rs3       (scheduler_0_output_m2sPipe_payload_rs3[4:0]        ), //i
    .io_inputs_0_payload_rd        (scheduler_0_output_m2sPipe_payload_rd[4:0]         ), //i
    .io_inputs_0_payload_format    (scheduler_0_output_m2sPipe_payload_format          ), //i
    .io_inputs_0_payload_roundMode (scheduler_0_output_m2sPipe_payload_roundMode[2:0]  ), //i
    .io_inputs_1_valid             (scheduler_1_output_m2sPipe_valid                   ), //i
    .io_inputs_1_ready             (cmdArbiter_arbiter_io_inputs_1_ready               ), //o
    .io_inputs_1_payload_opcode    (scheduler_1_output_m2sPipe_payload_opcode[3:0]     ), //i
    .io_inputs_1_payload_arg       (scheduler_1_output_m2sPipe_payload_arg[1:0]        ), //i
    .io_inputs_1_payload_rs1       (scheduler_1_output_m2sPipe_payload_rs1[4:0]        ), //i
    .io_inputs_1_payload_rs2       (scheduler_1_output_m2sPipe_payload_rs2[4:0]        ), //i
    .io_inputs_1_payload_rs3       (scheduler_1_output_m2sPipe_payload_rs3[4:0]        ), //i
    .io_inputs_1_payload_rd        (scheduler_1_output_m2sPipe_payload_rd[4:0]         ), //i
    .io_inputs_1_payload_format    (scheduler_1_output_m2sPipe_payload_format          ), //i
    .io_inputs_1_payload_roundMode (scheduler_1_output_m2sPipe_payload_roundMode[2:0]  ), //i
    .io_output_valid               (cmdArbiter_arbiter_io_output_valid                 ), //o
    .io_output_ready               (cmdArbiter_output_ready                            ), //i
    .io_output_payload_opcode      (cmdArbiter_arbiter_io_output_payload_opcode[3:0]   ), //o
    .io_output_payload_arg         (cmdArbiter_arbiter_io_output_payload_arg[1:0]      ), //o
    .io_output_payload_rs1         (cmdArbiter_arbiter_io_output_payload_rs1[4:0]      ), //o
    .io_output_payload_rs2         (cmdArbiter_arbiter_io_output_payload_rs2[4:0]      ), //o
    .io_output_payload_rs3         (cmdArbiter_arbiter_io_output_payload_rs3[4:0]      ), //o
    .io_output_payload_rd          (cmdArbiter_arbiter_io_output_payload_rd[4:0]       ), //o
    .io_output_payload_format      (cmdArbiter_arbiter_io_output_payload_format        ), //o
    .io_output_payload_roundMode   (cmdArbiter_arbiter_io_output_payload_roundMode[2:0]), //o
    .io_chosen                     (cmdArbiter_arbiter_io_chosen                       ), //o
    .io_chosenOH                   (cmdArbiter_arbiter_io_chosenOH[1:0]                ), //o
    .io_systemClk                  (io_systemClk                                       ), //i
    .systemCd_logic_outputReset    (systemCd_logic_outputReset                         )  //i
  );
  FpuDiv div_divider (
    .io_input_valid             (div_divider_io_input_valid                ), //i
    .io_input_ready             (div_divider_io_input_ready                ), //o
    .io_input_payload_a         (div_input_payload_rs1_mantissa[51:0]      ), //i
    .io_input_payload_b         (div_input_payload_rs2_mantissa[51:0]      ), //i
    .io_output_valid            (div_divider_io_output_valid               ), //o
    .io_output_ready            (div_input_ready                           ), //i
    .io_output_payload_result   (div_divider_io_output_payload_result[54:0]), //o
    .io_output_payload_remain   (div_divider_io_output_payload_remain[52:0]), //o
    .io_systemClk               (io_systemClk                              ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                )  //i
  );
  FpuSqrt sqrt_sqrt (
    .io_input_valid             (sqrt_sqrt_io_input_valid                ), //i
    .io_input_ready             (sqrt_sqrt_io_input_ready                ), //o
    .io_input_payload_a         (sqrt_sqrt_io_input_payload_a[53:0]      ), //i
    .io_output_valid            (sqrt_sqrt_io_output_valid               ), //o
    .io_output_ready            (sqrt_input_ready                        ), //i
    .io_output_payload_result   (sqrt_sqrt_io_output_payload_result[52:0]), //o
    .io_output_payload_remain   (sqrt_sqrt_io_output_payload_remain[56:0]), //o
    .io_systemClk               (io_systemClk                            ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset              )  //i
  );
  StreamArbiter_1 streamArbiter_10 (
    .io_inputs_0_valid                  (load_s1_output_m2sPipe_valid                           ), //i
    .io_inputs_0_ready                  (streamArbiter_10_io_inputs_0_ready                     ), //o
    .io_inputs_0_payload_source         (load_s1_output_m2sPipe_payload_source                  ), //i
    .io_inputs_0_payload_rd             (load_s1_output_m2sPipe_payload_rd[4:0]                 ), //i
    .io_inputs_0_payload_value_mantissa (load_s1_output_m2sPipe_payload_value_mantissa[52:0]    ), //i
    .io_inputs_0_payload_value_exponent (load_s1_output_m2sPipe_payload_value_exponent[11:0]    ), //i
    .io_inputs_0_payload_value_sign     (load_s1_output_m2sPipe_payload_value_sign              ), //i
    .io_inputs_0_payload_value_special  (load_s1_output_m2sPipe_payload_value_special           ), //i
    .io_inputs_0_payload_scrap          (load_s1_output_m2sPipe_payload_scrap                   ), //i
    .io_inputs_0_payload_roundMode      (load_s1_output_m2sPipe_payload_roundMode[2:0]          ), //i
    .io_inputs_0_payload_format         (load_s1_output_m2sPipe_payload_format                  ), //i
    .io_inputs_0_payload_NV             (load_s1_output_m2sPipe_payload_NV                      ), //i
    .io_inputs_0_payload_DZ             (load_s1_output_m2sPipe_payload_DZ                      ), //i
    .io_inputs_1_valid                  (sqrt_output_valid                                      ), //i
    .io_inputs_1_ready                  (streamArbiter_10_io_inputs_1_ready                     ), //o
    .io_inputs_1_payload_source         (sqrt_output_payload_source                             ), //i
    .io_inputs_1_payload_rd             (sqrt_output_payload_rd[4:0]                            ), //i
    .io_inputs_1_payload_value_mantissa (sqrt_output_payload_value_mantissa[52:0]               ), //i
    .io_inputs_1_payload_value_exponent (sqrt_output_payload_value_exponent[11:0]               ), //i
    .io_inputs_1_payload_value_sign     (sqrt_output_payload_value_sign                         ), //i
    .io_inputs_1_payload_value_special  (sqrt_output_payload_value_special                      ), //i
    .io_inputs_1_payload_scrap          (sqrt_output_payload_scrap                              ), //i
    .io_inputs_1_payload_roundMode      (sqrt_output_payload_roundMode[2:0]                     ), //i
    .io_inputs_1_payload_format         (sqrt_output_payload_format                             ), //i
    .io_inputs_1_payload_NV             (sqrt_output_payload_NV                                 ), //i
    .io_inputs_1_payload_DZ             (sqrt_output_payload_DZ                                 ), //i
    .io_inputs_2_valid                  (div_output_valid                                       ), //i
    .io_inputs_2_ready                  (streamArbiter_10_io_inputs_2_ready                     ), //o
    .io_inputs_2_payload_source         (div_output_payload_source                              ), //i
    .io_inputs_2_payload_rd             (div_output_payload_rd[4:0]                             ), //i
    .io_inputs_2_payload_value_mantissa (div_output_payload_value_mantissa[52:0]                ), //i
    .io_inputs_2_payload_value_exponent (div_output_payload_value_exponent[11:0]                ), //i
    .io_inputs_2_payload_value_sign     (div_output_payload_value_sign                          ), //i
    .io_inputs_2_payload_value_special  (div_output_payload_value_special                       ), //i
    .io_inputs_2_payload_scrap          (div_output_payload_scrap                               ), //i
    .io_inputs_2_payload_roundMode      (div_output_payload_roundMode[2:0]                      ), //i
    .io_inputs_2_payload_format         (div_output_payload_format                              ), //i
    .io_inputs_2_payload_NV             (div_output_payload_NV                                  ), //i
    .io_inputs_2_payload_DZ             (div_output_payload_DZ                                  ), //i
    .io_inputs_3_valid                  (add_result_output_valid                                ), //i
    .io_inputs_3_ready                  (streamArbiter_10_io_inputs_3_ready                     ), //o
    .io_inputs_3_payload_source         (add_result_output_payload_source                       ), //i
    .io_inputs_3_payload_rd             (add_result_output_payload_rd[4:0]                      ), //i
    .io_inputs_3_payload_value_mantissa (add_result_output_payload_value_mantissa[52:0]         ), //i
    .io_inputs_3_payload_value_exponent (add_result_output_payload_value_exponent[11:0]         ), //i
    .io_inputs_3_payload_value_sign     (add_result_output_payload_value_sign                   ), //i
    .io_inputs_3_payload_value_special  (add_result_output_payload_value_special                ), //i
    .io_inputs_3_payload_scrap          (add_result_output_payload_scrap                        ), //i
    .io_inputs_3_payload_roundMode      (add_result_output_payload_roundMode[2:0]               ), //i
    .io_inputs_3_payload_format         (add_result_output_payload_format                       ), //i
    .io_inputs_3_payload_NV             (add_result_output_payload_NV                           ), //i
    .io_inputs_3_payload_DZ             (add_result_output_payload_DZ                           ), //i
    .io_inputs_4_valid                  (mul_result_output_valid                                ), //i
    .io_inputs_4_ready                  (streamArbiter_10_io_inputs_4_ready                     ), //o
    .io_inputs_4_payload_source         (mul_result_output_payload_source                       ), //i
    .io_inputs_4_payload_rd             (mul_result_output_payload_rd[4:0]                      ), //i
    .io_inputs_4_payload_value_mantissa (mul_result_output_payload_value_mantissa[52:0]         ), //i
    .io_inputs_4_payload_value_exponent (mul_result_output_payload_value_exponent[11:0]         ), //i
    .io_inputs_4_payload_value_sign     (mul_result_output_payload_value_sign                   ), //i
    .io_inputs_4_payload_value_special  (mul_result_output_payload_value_special                ), //i
    .io_inputs_4_payload_scrap          (mul_result_output_payload_scrap                        ), //i
    .io_inputs_4_payload_roundMode      (mul_result_output_payload_roundMode[2:0]               ), //i
    .io_inputs_4_payload_format         (mul_result_output_payload_format                       ), //i
    .io_inputs_4_payload_NV             (mul_result_output_payload_NV                           ), //i
    .io_inputs_4_payload_DZ             (mul_result_output_payload_DZ                           ), //i
    .io_inputs_5_valid                  (shortPip_output_m2sPipe_valid                          ), //i
    .io_inputs_5_ready                  (streamArbiter_10_io_inputs_5_ready                     ), //o
    .io_inputs_5_payload_source         (shortPip_output_m2sPipe_payload_source                 ), //i
    .io_inputs_5_payload_rd             (shortPip_output_m2sPipe_payload_rd[4:0]                ), //i
    .io_inputs_5_payload_value_mantissa (shortPip_output_m2sPipe_payload_value_mantissa[52:0]   ), //i
    .io_inputs_5_payload_value_exponent (shortPip_output_m2sPipe_payload_value_exponent[11:0]   ), //i
    .io_inputs_5_payload_value_sign     (shortPip_output_m2sPipe_payload_value_sign             ), //i
    .io_inputs_5_payload_value_special  (shortPip_output_m2sPipe_payload_value_special          ), //i
    .io_inputs_5_payload_scrap          (shortPip_output_m2sPipe_payload_scrap                  ), //i
    .io_inputs_5_payload_roundMode      (shortPip_output_m2sPipe_payload_roundMode[2:0]         ), //i
    .io_inputs_5_payload_format         (shortPip_output_m2sPipe_payload_format                 ), //i
    .io_inputs_5_payload_NV             (shortPip_output_m2sPipe_payload_NV                     ), //i
    .io_inputs_5_payload_DZ             (shortPip_output_m2sPipe_payload_DZ                     ), //i
    .io_output_valid                    (streamArbiter_10_io_output_valid                       ), //o
    .io_output_ready                    (streamArbiter_10_io_output_combStage_ready             ), //i
    .io_output_payload_source           (streamArbiter_10_io_output_payload_source              ), //o
    .io_output_payload_rd               (streamArbiter_10_io_output_payload_rd[4:0]             ), //o
    .io_output_payload_value_mantissa   (streamArbiter_10_io_output_payload_value_mantissa[52:0]), //o
    .io_output_payload_value_exponent   (streamArbiter_10_io_output_payload_value_exponent[11:0]), //o
    .io_output_payload_value_sign       (streamArbiter_10_io_output_payload_value_sign          ), //o
    .io_output_payload_value_special    (streamArbiter_10_io_output_payload_value_special       ), //o
    .io_output_payload_scrap            (streamArbiter_10_io_output_payload_scrap               ), //o
    .io_output_payload_roundMode        (streamArbiter_10_io_output_payload_roundMode[2:0]      ), //o
    .io_output_payload_format           (streamArbiter_10_io_output_payload_format              ), //o
    .io_output_payload_NV               (streamArbiter_10_io_output_payload_NV                  ), //o
    .io_output_payload_DZ               (streamArbiter_10_io_output_payload_DZ                  ), //o
    .io_chosen                          (streamArbiter_10_io_chosen[2:0]                        ), //o
    .io_chosenOH                        (streamArbiter_10_io_chosenOH[5:0]                      ), //o
    .io_systemClk                       (io_systemClk                                           ), //i
    .systemCd_logic_outputReset         (systemCd_logic_outputReset                             )  //i
  );
  always @(*) begin
    case(load_s0_input_payload_source)
      1'b0 : begin
        _zz_load_s0_hazard = load_s0_filtred_0_valid;
        _zz_load_s0_output_payload_value = load_s0_filtred_0_payload_value;
      end
      default : begin
        _zz_load_s0_hazard = load_s0_filtred_1_valid;
        _zz_load_s0_output_payload_value = load_s0_filtred_1_payload_value;
      end
    endcase
  end

  always @(*) begin
    case(shortPip_input_payload_source)
      1'b0 : begin
        _zz_shortPip_isCommited = commitLogic_0_short_notEmpty;
        _zz_shortPip_input_ready = shortPip_rspStreams_0_ready;
      end
      default : begin
        _zz_shortPip_isCommited = commitLogic_1_short_notEmpty;
        _zz_shortPip_input_ready = shortPip_rspStreams_1_ready;
      end
    endcase
  end

  always @(*) begin
    case(mul_sum2_input_payload_source)
      1'b0 : _zz_mul_sum2_isCommited = commitLogic_0_mul_notEmpty;
      default : _zz_mul_sum2_isCommited = commitLogic_1_mul_notEmpty;
    endcase
  end

  always @(*) begin
    case(div_input_payload_source)
      1'b0 : _zz_div_isCommited = commitLogic_0_div_notEmpty;
      default : _zz_div_isCommited = commitLogic_1_div_notEmpty;
    endcase
  end

  always @(*) begin
    case(sqrt_input_payload_source)
      1'b0 : _zz_sqrt_isCommited = commitLogic_0_sqrt_notEmpty;
      default : _zz_sqrt_isCommited = commitLogic_1_sqrt_notEmpty;
    endcase
  end

  always @(*) begin
    case(add_oh_input_payload_source)
      1'b0 : _zz_add_oh_isCommited = commitLogic_0_add_notEmpty;
      default : _zz_add_oh_isCommited = commitLogic_1_add_notEmpty;
    endcase
  end

  always @(*) begin
    case(roundBack_input_payload_source)
      1'b0 : _zz_roundBack_write = roundBack_writes_0;
      default : _zz_roundBack_write = roundBack_writes_1;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_port_0_cmd_payload_opcode)
      FpuOpcode_LOAD : io_port_0_cmd_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_port_0_cmd_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_port_0_cmd_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_port_0_cmd_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_port_0_cmd_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_port_0_cmd_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_port_0_cmd_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_port_0_cmd_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_port_0_cmd_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_port_0_cmd_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_port_0_cmd_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_port_0_cmd_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_port_0_cmd_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_port_0_cmd_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_port_0_cmd_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_port_0_cmd_payload_opcode_string = "FCVT_X_X";
      default : io_port_0_cmd_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_port_0_cmd_payload_format)
      FpuFormat_FLOAT : io_port_0_cmd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_port_0_cmd_payload_format_string = "DOUBLE";
      default : io_port_0_cmd_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_port_0_cmd_payload_roundMode)
      FpuRoundMode_RNE : io_port_0_cmd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_port_0_cmd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_port_0_cmd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_port_0_cmd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_port_0_cmd_payload_roundMode_string = "RMM";
      default : io_port_0_cmd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_port_0_commit_payload_opcode)
      FpuOpcode_LOAD : io_port_0_commit_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_port_0_commit_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_port_0_commit_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_port_0_commit_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_port_0_commit_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_port_0_commit_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_port_0_commit_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_port_0_commit_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_port_0_commit_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_port_0_commit_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_port_0_commit_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_port_0_commit_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_port_0_commit_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_port_0_commit_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_port_0_commit_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_port_0_commit_payload_opcode_string = "FCVT_X_X";
      default : io_port_0_commit_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_port_1_cmd_payload_opcode)
      FpuOpcode_LOAD : io_port_1_cmd_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_port_1_cmd_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_port_1_cmd_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_port_1_cmd_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_port_1_cmd_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_port_1_cmd_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_port_1_cmd_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_port_1_cmd_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_port_1_cmd_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_port_1_cmd_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_port_1_cmd_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_port_1_cmd_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_port_1_cmd_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_port_1_cmd_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_port_1_cmd_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_port_1_cmd_payload_opcode_string = "FCVT_X_X";
      default : io_port_1_cmd_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_port_1_cmd_payload_format)
      FpuFormat_FLOAT : io_port_1_cmd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_port_1_cmd_payload_format_string = "DOUBLE";
      default : io_port_1_cmd_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_port_1_cmd_payload_roundMode)
      FpuRoundMode_RNE : io_port_1_cmd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_port_1_cmd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_port_1_cmd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_port_1_cmd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_port_1_cmd_payload_roundMode_string = "RMM";
      default : io_port_1_cmd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_port_1_commit_payload_opcode)
      FpuOpcode_LOAD : io_port_1_commit_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_port_1_commit_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_port_1_commit_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_port_1_commit_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_port_1_commit_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_port_1_commit_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_port_1_commit_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_port_1_commit_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_port_1_commit_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_port_1_commit_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_port_1_commit_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_port_1_commit_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_port_1_commit_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_port_1_commit_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_port_1_commit_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_port_1_commit_payload_opcode_string = "FCVT_X_X";
      default : io_port_1_commit_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(commitFork_load_0_payload_opcode)
      FpuOpcode_LOAD : commitFork_load_0_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : commitFork_load_0_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : commitFork_load_0_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : commitFork_load_0_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : commitFork_load_0_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : commitFork_load_0_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : commitFork_load_0_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : commitFork_load_0_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : commitFork_load_0_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : commitFork_load_0_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : commitFork_load_0_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : commitFork_load_0_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : commitFork_load_0_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : commitFork_load_0_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : commitFork_load_0_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : commitFork_load_0_payload_opcode_string = "FCVT_X_X";
      default : commitFork_load_0_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(commitFork_load_1_payload_opcode)
      FpuOpcode_LOAD : commitFork_load_1_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : commitFork_load_1_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : commitFork_load_1_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : commitFork_load_1_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : commitFork_load_1_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : commitFork_load_1_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : commitFork_load_1_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : commitFork_load_1_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : commitFork_load_1_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : commitFork_load_1_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : commitFork_load_1_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : commitFork_load_1_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : commitFork_load_1_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : commitFork_load_1_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : commitFork_load_1_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : commitFork_load_1_payload_opcode_string = "FCVT_X_X";
      default : commitFork_load_1_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(commitFork_commit_0_payload_opcode)
      FpuOpcode_LOAD : commitFork_commit_0_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : commitFork_commit_0_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : commitFork_commit_0_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : commitFork_commit_0_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : commitFork_commit_0_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : commitFork_commit_0_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : commitFork_commit_0_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : commitFork_commit_0_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : commitFork_commit_0_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : commitFork_commit_0_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : commitFork_commit_0_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : commitFork_commit_0_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : commitFork_commit_0_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : commitFork_commit_0_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : commitFork_commit_0_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : commitFork_commit_0_payload_opcode_string = "FCVT_X_X";
      default : commitFork_commit_0_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(commitFork_commit_1_payload_opcode)
      FpuOpcode_LOAD : commitFork_commit_1_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : commitFork_commit_1_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : commitFork_commit_1_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : commitFork_commit_1_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : commitFork_commit_1_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : commitFork_commit_1_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : commitFork_commit_1_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : commitFork_commit_1_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : commitFork_commit_1_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : commitFork_commit_1_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : commitFork_commit_1_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : commitFork_commit_1_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : commitFork_commit_1_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : commitFork_commit_1_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : commitFork_commit_1_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : commitFork_commit_1_payload_opcode_string = "FCVT_X_X";
      default : commitFork_commit_1_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(streamFork_3_io_outputs_1_s2mPipe_payload_opcode)
      FpuOpcode_LOAD : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "FCVT_X_X";
      default : streamFork_3_io_outputs_1_s2mPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(streamFork_3_io_outputs_1_rData_opcode)
      FpuOpcode_LOAD : streamFork_3_io_outputs_1_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : streamFork_3_io_outputs_1_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : streamFork_3_io_outputs_1_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : streamFork_3_io_outputs_1_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : streamFork_3_io_outputs_1_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : streamFork_3_io_outputs_1_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : streamFork_3_io_outputs_1_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : streamFork_3_io_outputs_1_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : streamFork_3_io_outputs_1_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : streamFork_3_io_outputs_1_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : streamFork_3_io_outputs_1_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : streamFork_3_io_outputs_1_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : streamFork_3_io_outputs_1_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : streamFork_3_io_outputs_1_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : streamFork_3_io_outputs_1_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : streamFork_3_io_outputs_1_rData_opcode_string = "FCVT_X_X";
      default : streamFork_3_io_outputs_1_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_opcode)
      FpuOpcode_LOAD : _zz_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_payload_opcode_string = "FCVT_X_X";
      default : _zz_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(streamFork_4_io_outputs_1_s2mPipe_payload_opcode)
      FpuOpcode_LOAD : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "FCVT_X_X";
      default : streamFork_4_io_outputs_1_s2mPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(streamFork_4_io_outputs_1_rData_opcode)
      FpuOpcode_LOAD : streamFork_4_io_outputs_1_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : streamFork_4_io_outputs_1_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : streamFork_4_io_outputs_1_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : streamFork_4_io_outputs_1_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : streamFork_4_io_outputs_1_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : streamFork_4_io_outputs_1_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : streamFork_4_io_outputs_1_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : streamFork_4_io_outputs_1_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : streamFork_4_io_outputs_1_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : streamFork_4_io_outputs_1_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : streamFork_4_io_outputs_1_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : streamFork_4_io_outputs_1_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : streamFork_4_io_outputs_1_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : streamFork_4_io_outputs_1_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : streamFork_4_io_outputs_1_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : streamFork_4_io_outputs_1_rData_opcode_string = "FCVT_X_X";
      default : streamFork_4_io_outputs_1_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_payload_opcode_1)
      FpuOpcode_LOAD : _zz_payload_opcode_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_payload_opcode_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_payload_opcode_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_payload_opcode_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_payload_opcode_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_payload_opcode_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_payload_opcode_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_payload_opcode_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_payload_opcode_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_payload_opcode_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_payload_opcode_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_payload_opcode_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_payload_opcode_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_payload_opcode_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_payload_opcode_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_payload_opcode_1_string = "FCVT_X_X";
      default : _zz_payload_opcode_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_commitLogic_0_input_payload_opcode)
      FpuOpcode_LOAD : _zz_commitLogic_0_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_commitLogic_0_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_commitLogic_0_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_commitLogic_0_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_commitLogic_0_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_commitLogic_0_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_commitLogic_0_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_commitLogic_0_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_commitLogic_0_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_commitLogic_0_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_commitLogic_0_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_commitLogic_0_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_commitLogic_0_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_commitLogic_0_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_commitLogic_0_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_commitLogic_0_input_payload_opcode_string = "FCVT_X_X";
      default : _zz_commitLogic_0_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(commitLogic_0_input_payload_opcode)
      FpuOpcode_LOAD : commitLogic_0_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : commitLogic_0_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : commitLogic_0_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : commitLogic_0_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : commitLogic_0_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : commitLogic_0_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : commitLogic_0_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : commitLogic_0_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : commitLogic_0_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : commitLogic_0_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : commitLogic_0_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : commitLogic_0_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : commitLogic_0_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : commitLogic_0_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : commitLogic_0_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : commitLogic_0_input_payload_opcode_string = "FCVT_X_X";
      default : commitLogic_0_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_commitLogic_1_input_payload_opcode)
      FpuOpcode_LOAD : _zz_commitLogic_1_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_commitLogic_1_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_commitLogic_1_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_commitLogic_1_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_commitLogic_1_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_commitLogic_1_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_commitLogic_1_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_commitLogic_1_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_commitLogic_1_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_commitLogic_1_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_commitLogic_1_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_commitLogic_1_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_commitLogic_1_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_commitLogic_1_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_commitLogic_1_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_commitLogic_1_input_payload_opcode_string = "FCVT_X_X";
      default : _zz_commitLogic_1_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(commitLogic_1_input_payload_opcode)
      FpuOpcode_LOAD : commitLogic_1_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : commitLogic_1_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : commitLogic_1_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : commitLogic_1_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : commitLogic_1_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : commitLogic_1_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : commitLogic_1_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : commitLogic_1_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : commitLogic_1_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : commitLogic_1_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : commitLogic_1_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : commitLogic_1_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : commitLogic_1_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : commitLogic_1_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : commitLogic_1_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : commitLogic_1_input_payload_opcode_string = "FCVT_X_X";
      default : commitLogic_1_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_input_payload_opcode)
      FpuOpcode_LOAD : scheduler_0_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_0_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_0_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_0_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_0_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_0_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_0_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_0_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_0_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_0_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_0_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_0_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_0_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_0_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_0_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_0_input_payload_opcode_string = "FCVT_X_X";
      default : scheduler_0_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_input_payload_format)
      FpuFormat_FLOAT : scheduler_0_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_0_input_payload_format_string = "DOUBLE";
      default : scheduler_0_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_input_payload_roundMode)
      FpuRoundMode_RNE : scheduler_0_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_0_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_0_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_0_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_0_input_payload_roundMode_string = "RMM";
      default : scheduler_0_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_port_0_cmd_rData_opcode)
      FpuOpcode_LOAD : io_port_0_cmd_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_port_0_cmd_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_port_0_cmd_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_port_0_cmd_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_port_0_cmd_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_port_0_cmd_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_port_0_cmd_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_port_0_cmd_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_port_0_cmd_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_port_0_cmd_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_port_0_cmd_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_port_0_cmd_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_port_0_cmd_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_port_0_cmd_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_port_0_cmd_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_port_0_cmd_rData_opcode_string = "FCVT_X_X";
      default : io_port_0_cmd_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_port_0_cmd_rData_format)
      FpuFormat_FLOAT : io_port_0_cmd_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_port_0_cmd_rData_format_string = "DOUBLE";
      default : io_port_0_cmd_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_port_0_cmd_rData_roundMode)
      FpuRoundMode_RNE : io_port_0_cmd_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_port_0_cmd_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_port_0_cmd_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_port_0_cmd_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_port_0_cmd_rData_roundMode_string = "RMM";
      default : io_port_0_cmd_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_scheduler_0_input_payload_opcode)
      FpuOpcode_LOAD : _zz_scheduler_0_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_scheduler_0_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_scheduler_0_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_scheduler_0_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_scheduler_0_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_scheduler_0_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_scheduler_0_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_scheduler_0_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_scheduler_0_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_scheduler_0_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_scheduler_0_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_scheduler_0_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_scheduler_0_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_scheduler_0_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_scheduler_0_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_scheduler_0_input_payload_opcode_string = "FCVT_X_X";
      default : _zz_scheduler_0_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_scheduler_0_input_payload_format)
      FpuFormat_FLOAT : _zz_scheduler_0_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_scheduler_0_input_payload_format_string = "DOUBLE";
      default : _zz_scheduler_0_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_scheduler_0_input_payload_roundMode)
      FpuRoundMode_RNE : _zz_scheduler_0_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : _zz_scheduler_0_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : _zz_scheduler_0_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : _zz_scheduler_0_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : _zz_scheduler_0_input_payload_roundMode_string = "RMM";
      default : _zz_scheduler_0_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_payload_opcode)
      FpuOpcode_LOAD : scheduler_0_output_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_0_output_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_0_output_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_0_output_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_0_output_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_0_output_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_0_output_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_0_output_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_0_output_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_0_output_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_0_output_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_0_output_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_0_output_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_0_output_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_0_output_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_0_output_payload_opcode_string = "FCVT_X_X";
      default : scheduler_0_output_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_payload_format)
      FpuFormat_FLOAT : scheduler_0_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_0_output_payload_format_string = "DOUBLE";
      default : scheduler_0_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_payload_roundMode)
      FpuRoundMode_RNE : scheduler_0_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_0_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_0_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_0_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_0_output_payload_roundMode_string = "RMM";
      default : scheduler_0_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(scheduler_1_input_payload_opcode)
      FpuOpcode_LOAD : scheduler_1_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_1_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_1_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_1_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_1_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_1_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_1_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_1_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_1_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_1_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_1_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_1_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_1_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_1_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_1_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_1_input_payload_opcode_string = "FCVT_X_X";
      default : scheduler_1_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_input_payload_format)
      FpuFormat_FLOAT : scheduler_1_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_1_input_payload_format_string = "DOUBLE";
      default : scheduler_1_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_input_payload_roundMode)
      FpuRoundMode_RNE : scheduler_1_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_1_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_1_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_1_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_1_input_payload_roundMode_string = "RMM";
      default : scheduler_1_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_port_1_cmd_rData_opcode)
      FpuOpcode_LOAD : io_port_1_cmd_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_port_1_cmd_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_port_1_cmd_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_port_1_cmd_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_port_1_cmd_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_port_1_cmd_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_port_1_cmd_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_port_1_cmd_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_port_1_cmd_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_port_1_cmd_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_port_1_cmd_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_port_1_cmd_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_port_1_cmd_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_port_1_cmd_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_port_1_cmd_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_port_1_cmd_rData_opcode_string = "FCVT_X_X";
      default : io_port_1_cmd_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_port_1_cmd_rData_format)
      FpuFormat_FLOAT : io_port_1_cmd_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_port_1_cmd_rData_format_string = "DOUBLE";
      default : io_port_1_cmd_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_port_1_cmd_rData_roundMode)
      FpuRoundMode_RNE : io_port_1_cmd_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_port_1_cmd_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_port_1_cmd_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_port_1_cmd_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_port_1_cmd_rData_roundMode_string = "RMM";
      default : io_port_1_cmd_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_scheduler_1_input_payload_opcode)
      FpuOpcode_LOAD : _zz_scheduler_1_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_scheduler_1_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_scheduler_1_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_scheduler_1_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_scheduler_1_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_scheduler_1_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_scheduler_1_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_scheduler_1_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_scheduler_1_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_scheduler_1_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_scheduler_1_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_scheduler_1_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_scheduler_1_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_scheduler_1_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_scheduler_1_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_scheduler_1_input_payload_opcode_string = "FCVT_X_X";
      default : _zz_scheduler_1_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_scheduler_1_input_payload_format)
      FpuFormat_FLOAT : _zz_scheduler_1_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_scheduler_1_input_payload_format_string = "DOUBLE";
      default : _zz_scheduler_1_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_scheduler_1_input_payload_roundMode)
      FpuRoundMode_RNE : _zz_scheduler_1_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : _zz_scheduler_1_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : _zz_scheduler_1_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : _zz_scheduler_1_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : _zz_scheduler_1_input_payload_roundMode_string = "RMM";
      default : _zz_scheduler_1_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_payload_opcode)
      FpuOpcode_LOAD : scheduler_1_output_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_1_output_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_1_output_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_1_output_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_1_output_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_1_output_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_1_output_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_1_output_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_1_output_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_1_output_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_1_output_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_1_output_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_1_output_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_1_output_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_1_output_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_1_output_payload_opcode_string = "FCVT_X_X";
      default : scheduler_1_output_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_payload_format)
      FpuFormat_FLOAT : scheduler_1_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_1_output_payload_format_string = "DOUBLE";
      default : scheduler_1_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_payload_roundMode)
      FpuRoundMode_RNE : scheduler_1_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_1_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_1_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_1_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_1_output_payload_roundMode_string = "RMM";
      default : scheduler_1_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_m2sPipe_payload_opcode)
      FpuOpcode_LOAD : scheduler_0_output_m2sPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_0_output_m2sPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_0_output_m2sPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_0_output_m2sPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_0_output_m2sPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_0_output_m2sPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_0_output_m2sPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_0_output_m2sPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_0_output_m2sPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_0_output_m2sPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_0_output_m2sPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_0_output_m2sPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_0_output_m2sPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_0_output_m2sPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_0_output_m2sPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_0_output_m2sPipe_payload_opcode_string = "FCVT_X_X";
      default : scheduler_0_output_m2sPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_m2sPipe_payload_format)
      FpuFormat_FLOAT : scheduler_0_output_m2sPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_0_output_m2sPipe_payload_format_string = "DOUBLE";
      default : scheduler_0_output_m2sPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_m2sPipe_payload_roundMode)
      FpuRoundMode_RNE : scheduler_0_output_m2sPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_0_output_m2sPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_0_output_m2sPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_0_output_m2sPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_0_output_m2sPipe_payload_roundMode_string = "RMM";
      default : scheduler_0_output_m2sPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_rData_opcode)
      FpuOpcode_LOAD : scheduler_0_output_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_0_output_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_0_output_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_0_output_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_0_output_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_0_output_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_0_output_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_0_output_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_0_output_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_0_output_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_0_output_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_0_output_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_0_output_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_0_output_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_0_output_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_0_output_rData_opcode_string = "FCVT_X_X";
      default : scheduler_0_output_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_rData_format)
      FpuFormat_FLOAT : scheduler_0_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_0_output_rData_format_string = "DOUBLE";
      default : scheduler_0_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_0_output_rData_roundMode)
      FpuRoundMode_RNE : scheduler_0_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_0_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_0_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_0_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_0_output_rData_roundMode_string = "RMM";
      default : scheduler_0_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_m2sPipe_payload_opcode)
      FpuOpcode_LOAD : scheduler_1_output_m2sPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_1_output_m2sPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_1_output_m2sPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_1_output_m2sPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_1_output_m2sPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_1_output_m2sPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_1_output_m2sPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_1_output_m2sPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_1_output_m2sPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_1_output_m2sPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_1_output_m2sPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_1_output_m2sPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_1_output_m2sPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_1_output_m2sPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_1_output_m2sPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_1_output_m2sPipe_payload_opcode_string = "FCVT_X_X";
      default : scheduler_1_output_m2sPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_m2sPipe_payload_format)
      FpuFormat_FLOAT : scheduler_1_output_m2sPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_1_output_m2sPipe_payload_format_string = "DOUBLE";
      default : scheduler_1_output_m2sPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_m2sPipe_payload_roundMode)
      FpuRoundMode_RNE : scheduler_1_output_m2sPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_1_output_m2sPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_1_output_m2sPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_1_output_m2sPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_1_output_m2sPipe_payload_roundMode_string = "RMM";
      default : scheduler_1_output_m2sPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_rData_opcode)
      FpuOpcode_LOAD : scheduler_1_output_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : scheduler_1_output_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : scheduler_1_output_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : scheduler_1_output_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : scheduler_1_output_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : scheduler_1_output_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : scheduler_1_output_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : scheduler_1_output_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : scheduler_1_output_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : scheduler_1_output_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : scheduler_1_output_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : scheduler_1_output_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : scheduler_1_output_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : scheduler_1_output_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : scheduler_1_output_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : scheduler_1_output_rData_opcode_string = "FCVT_X_X";
      default : scheduler_1_output_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_rData_format)
      FpuFormat_FLOAT : scheduler_1_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : scheduler_1_output_rData_format_string = "DOUBLE";
      default : scheduler_1_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(scheduler_1_output_rData_roundMode)
      FpuRoundMode_RNE : scheduler_1_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : scheduler_1_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : scheduler_1_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : scheduler_1_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : scheduler_1_output_rData_roundMode_string = "RMM";
      default : scheduler_1_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(cmdArbiter_output_payload_opcode)
      FpuOpcode_LOAD : cmdArbiter_output_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : cmdArbiter_output_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : cmdArbiter_output_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : cmdArbiter_output_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : cmdArbiter_output_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : cmdArbiter_output_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : cmdArbiter_output_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : cmdArbiter_output_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : cmdArbiter_output_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : cmdArbiter_output_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : cmdArbiter_output_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : cmdArbiter_output_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : cmdArbiter_output_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : cmdArbiter_output_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : cmdArbiter_output_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : cmdArbiter_output_payload_opcode_string = "FCVT_X_X";
      default : cmdArbiter_output_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(cmdArbiter_output_payload_roundMode)
      FpuRoundMode_RNE : cmdArbiter_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : cmdArbiter_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : cmdArbiter_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : cmdArbiter_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : cmdArbiter_output_payload_roundMode_string = "RMM";
      default : cmdArbiter_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(cmdArbiter_output_payload_format)
      FpuFormat_FLOAT : cmdArbiter_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : cmdArbiter_output_payload_format_string = "DOUBLE";
      default : cmdArbiter_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(read_s0_payload_opcode)
      FpuOpcode_LOAD : read_s0_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : read_s0_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : read_s0_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : read_s0_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : read_s0_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : read_s0_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : read_s0_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : read_s0_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : read_s0_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : read_s0_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : read_s0_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : read_s0_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : read_s0_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : read_s0_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : read_s0_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : read_s0_payload_opcode_string = "FCVT_X_X";
      default : read_s0_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(read_s0_payload_roundMode)
      FpuRoundMode_RNE : read_s0_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : read_s0_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : read_s0_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : read_s0_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : read_s0_payload_roundMode_string = "RMM";
      default : read_s0_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(read_s0_payload_format)
      FpuFormat_FLOAT : read_s0_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : read_s0_payload_format_string = "DOUBLE";
      default : read_s0_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(read_s1_payload_opcode)
      FpuOpcode_LOAD : read_s1_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : read_s1_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : read_s1_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : read_s1_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : read_s1_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : read_s1_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : read_s1_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : read_s1_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : read_s1_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : read_s1_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : read_s1_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : read_s1_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : read_s1_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : read_s1_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : read_s1_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : read_s1_payload_opcode_string = "FCVT_X_X";
      default : read_s1_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(read_s1_payload_roundMode)
      FpuRoundMode_RNE : read_s1_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : read_s1_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : read_s1_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : read_s1_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : read_s1_payload_roundMode_string = "RMM";
      default : read_s1_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(read_s1_payload_format)
      FpuFormat_FLOAT : read_s1_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : read_s1_payload_format_string = "DOUBLE";
      default : read_s1_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(read_s0_rData_opcode)
      FpuOpcode_LOAD : read_s0_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : read_s0_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : read_s0_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : read_s0_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : read_s0_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : read_s0_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : read_s0_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : read_s0_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : read_s0_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : read_s0_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : read_s0_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : read_s0_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : read_s0_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : read_s0_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : read_s0_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : read_s0_rData_opcode_string = "FCVT_X_X";
      default : read_s0_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(read_s0_rData_roundMode)
      FpuRoundMode_RNE : read_s0_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : read_s0_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : read_s0_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : read_s0_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : read_s0_rData_roundMode_string = "RMM";
      default : read_s0_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(read_s0_rData_format)
      FpuFormat_FLOAT : read_s0_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : read_s0_rData_format_string = "DOUBLE";
      default : read_s0_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(read_output_payload_opcode)
      FpuOpcode_LOAD : read_output_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : read_output_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : read_output_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : read_output_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : read_output_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : read_output_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : read_output_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : read_output_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : read_output_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : read_output_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : read_output_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : read_output_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : read_output_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : read_output_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : read_output_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : read_output_payload_opcode_string = "FCVT_X_X";
      default : read_output_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(read_output_payload_roundMode)
      FpuRoundMode_RNE : read_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : read_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : read_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : read_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : read_output_payload_roundMode_string = "RMM";
      default : read_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(read_output_payload_format)
      FpuFormat_FLOAT : read_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : read_output_payload_format_string = "DOUBLE";
      default : read_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_read_output_payload_format)
      FpuFormat_FLOAT : _zz_read_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_read_output_payload_format_string = "DOUBLE";
      default : _zz_read_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_input_payload_opcode)
      FpuOpcode_LOAD : decode_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : decode_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : decode_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : decode_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : decode_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : decode_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : decode_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : decode_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : decode_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : decode_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : decode_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : decode_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : decode_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : decode_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : decode_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : decode_input_payload_opcode_string = "FCVT_X_X";
      default : decode_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_input_payload_roundMode)
      FpuRoundMode_RNE : decode_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_input_payload_roundMode_string = "RMM";
      default : decode_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_input_payload_format)
      FpuFormat_FLOAT : decode_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_input_payload_format_string = "DOUBLE";
      default : decode_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_load_payload_roundMode)
      FpuRoundMode_RNE : decode_load_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_load_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_load_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_load_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_load_payload_roundMode_string = "RMM";
      default : decode_load_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_load_payload_format)
      FpuFormat_FLOAT : decode_load_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_load_payload_format_string = "DOUBLE";
      default : decode_load_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_shortPip_payload_opcode)
      FpuOpcode_LOAD : decode_shortPip_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : decode_shortPip_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : decode_shortPip_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : decode_shortPip_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : decode_shortPip_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : decode_shortPip_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : decode_shortPip_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : decode_shortPip_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : decode_shortPip_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : decode_shortPip_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : decode_shortPip_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : decode_shortPip_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : decode_shortPip_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : decode_shortPip_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : decode_shortPip_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : decode_shortPip_payload_opcode_string = "FCVT_X_X";
      default : decode_shortPip_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_shortPip_payload_roundMode)
      FpuRoundMode_RNE : decode_shortPip_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_shortPip_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_shortPip_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_shortPip_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_shortPip_payload_roundMode_string = "RMM";
      default : decode_shortPip_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_shortPip_payload_format)
      FpuFormat_FLOAT : decode_shortPip_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_shortPip_payload_format_string = "DOUBLE";
      default : decode_shortPip_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_divSqrt_payload_roundMode)
      FpuRoundMode_RNE : decode_divSqrt_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_divSqrt_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_divSqrt_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_divSqrt_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_divSqrt_payload_roundMode_string = "RMM";
      default : decode_divSqrt_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_divSqrt_payload_format)
      FpuFormat_FLOAT : decode_divSqrt_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_divSqrt_payload_format_string = "DOUBLE";
      default : decode_divSqrt_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_div_payload_roundMode)
      FpuRoundMode_RNE : decode_div_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_div_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_div_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_div_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_div_payload_roundMode_string = "RMM";
      default : decode_div_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_div_payload_format)
      FpuFormat_FLOAT : decode_div_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_div_payload_format_string = "DOUBLE";
      default : decode_div_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_sqrt_payload_roundMode)
      FpuRoundMode_RNE : decode_sqrt_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_sqrt_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_sqrt_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_sqrt_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_sqrt_payload_roundMode_string = "RMM";
      default : decode_sqrt_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_sqrt_payload_format)
      FpuFormat_FLOAT : decode_sqrt_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_sqrt_payload_format_string = "DOUBLE";
      default : decode_sqrt_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_mul_payload_roundMode)
      FpuRoundMode_RNE : decode_mul_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_mul_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_mul_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_mul_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_mul_payload_roundMode_string = "RMM";
      default : decode_mul_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_mul_payload_format)
      FpuFormat_FLOAT : decode_mul_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_mul_payload_format_string = "DOUBLE";
      default : decode_mul_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_divSqrtToMul_payload_roundMode)
      FpuRoundMode_RNE : decode_divSqrtToMul_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_divSqrtToMul_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_divSqrtToMul_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_divSqrtToMul_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_divSqrtToMul_payload_roundMode_string = "RMM";
      default : decode_divSqrtToMul_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_divSqrtToMul_payload_format)
      FpuFormat_FLOAT : decode_divSqrtToMul_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_divSqrtToMul_payload_format_string = "DOUBLE";
      default : decode_divSqrtToMul_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_add_payload_roundMode)
      FpuRoundMode_RNE : decode_add_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_add_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_add_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_add_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_add_payload_roundMode_string = "RMM";
      default : decode_add_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_add_payload_format)
      FpuFormat_FLOAT : decode_add_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_add_payload_format_string = "DOUBLE";
      default : decode_add_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_mulToAdd_payload_roundMode)
      FpuRoundMode_RNE : decode_mulToAdd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_mulToAdd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_mulToAdd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_mulToAdd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_mulToAdd_payload_roundMode_string = "RMM";
      default : decode_mulToAdd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_mulToAdd_payload_format)
      FpuFormat_FLOAT : decode_mulToAdd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_mulToAdd_payload_format_string = "DOUBLE";
      default : decode_mulToAdd_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_payload_roundMode)
      FpuRoundMode_RNE : decode_load_s2mPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_load_s2mPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_load_s2mPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_load_s2mPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_load_s2mPipe_payload_roundMode_string = "RMM";
      default : decode_load_s2mPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_payload_format)
      FpuFormat_FLOAT : decode_load_s2mPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_load_s2mPipe_payload_format_string = "DOUBLE";
      default : decode_load_s2mPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_load_rData_roundMode)
      FpuRoundMode_RNE : decode_load_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_load_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_load_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_load_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_load_rData_roundMode_string = "RMM";
      default : decode_load_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_load_rData_format)
      FpuFormat_FLOAT : decode_load_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_load_rData_format_string = "DOUBLE";
      default : decode_load_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_load_s2mPipe_payload_roundMode)
      FpuRoundMode_RNE : _zz_decode_load_s2mPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : _zz_decode_load_s2mPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : _zz_decode_load_s2mPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : _zz_decode_load_s2mPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : _zz_decode_load_s2mPipe_payload_roundMode_string = "RMM";
      default : _zz_decode_load_s2mPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_load_s2mPipe_payload_format)
      FpuFormat_FLOAT : _zz_decode_load_s2mPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_decode_load_s2mPipe_payload_format_string = "DOUBLE";
      default : _zz_decode_load_s2mPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_m2sPipe_payload_roundMode)
      FpuRoundMode_RNE : decode_load_s2mPipe_m2sPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_load_s2mPipe_m2sPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_load_s2mPipe_m2sPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_load_s2mPipe_m2sPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_load_s2mPipe_m2sPipe_payload_roundMode_string = "RMM";
      default : decode_load_s2mPipe_m2sPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_m2sPipe_payload_format)
      FpuFormat_FLOAT : decode_load_s2mPipe_m2sPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_load_s2mPipe_m2sPipe_payload_format_string = "DOUBLE";
      default : decode_load_s2mPipe_m2sPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_rData_roundMode)
      FpuRoundMode_RNE : decode_load_s2mPipe_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_load_s2mPipe_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_load_s2mPipe_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_load_s2mPipe_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_load_s2mPipe_rData_roundMode_string = "RMM";
      default : decode_load_s2mPipe_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_rData_format)
      FpuFormat_FLOAT : decode_load_s2mPipe_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_load_s2mPipe_rData_format_string = "DOUBLE";
      default : decode_load_s2mPipe_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(load_s0_input_payload_roundMode)
      FpuRoundMode_RNE : load_s0_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : load_s0_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : load_s0_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : load_s0_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : load_s0_input_payload_roundMode_string = "RMM";
      default : load_s0_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(load_s0_input_payload_format)
      FpuFormat_FLOAT : load_s0_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : load_s0_input_payload_format_string = "DOUBLE";
      default : load_s0_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_m2sPipe_rData_roundMode)
      FpuRoundMode_RNE : decode_load_s2mPipe_m2sPipe_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_load_s2mPipe_m2sPipe_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_load_s2mPipe_m2sPipe_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_load_s2mPipe_m2sPipe_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_load_s2mPipe_m2sPipe_rData_roundMode_string = "RMM";
      default : decode_load_s2mPipe_m2sPipe_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_load_s2mPipe_m2sPipe_rData_format)
      FpuFormat_FLOAT : decode_load_s2mPipe_m2sPipe_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_load_s2mPipe_m2sPipe_rData_format_string = "DOUBLE";
      default : decode_load_s2mPipe_m2sPipe_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(load_s0_filtred_0_payload_opcode)
      FpuOpcode_LOAD : load_s0_filtred_0_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : load_s0_filtred_0_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : load_s0_filtred_0_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : load_s0_filtred_0_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : load_s0_filtred_0_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : load_s0_filtred_0_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : load_s0_filtred_0_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : load_s0_filtred_0_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : load_s0_filtred_0_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : load_s0_filtred_0_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : load_s0_filtred_0_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : load_s0_filtred_0_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : load_s0_filtred_0_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : load_s0_filtred_0_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : load_s0_filtred_0_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : load_s0_filtred_0_payload_opcode_string = "FCVT_X_X";
      default : load_s0_filtred_0_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(load_s0_filtred_1_payload_opcode)
      FpuOpcode_LOAD : load_s0_filtred_1_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : load_s0_filtred_1_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : load_s0_filtred_1_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : load_s0_filtred_1_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : load_s0_filtred_1_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : load_s0_filtred_1_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : load_s0_filtred_1_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : load_s0_filtred_1_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : load_s0_filtred_1_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : load_s0_filtred_1_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : load_s0_filtred_1_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : load_s0_filtred_1_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : load_s0_filtred_1_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : load_s0_filtred_1_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : load_s0_filtred_1_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : load_s0_filtred_1_payload_opcode_string = "FCVT_X_X";
      default : load_s0_filtred_1_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(load_s0_output_payload_roundMode)
      FpuRoundMode_RNE : load_s0_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : load_s0_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : load_s0_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : load_s0_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : load_s0_output_payload_roundMode_string = "RMM";
      default : load_s0_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(load_s0_output_payload_format)
      FpuFormat_FLOAT : load_s0_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : load_s0_output_payload_format_string = "DOUBLE";
      default : load_s0_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(load_s1_input_payload_roundMode)
      FpuRoundMode_RNE : load_s1_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : load_s1_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : load_s1_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : load_s1_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : load_s1_input_payload_roundMode_string = "RMM";
      default : load_s1_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(load_s1_input_payload_format)
      FpuFormat_FLOAT : load_s1_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : load_s1_input_payload_format_string = "DOUBLE";
      default : load_s1_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(load_s0_output_rData_roundMode)
      FpuRoundMode_RNE : load_s0_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : load_s0_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : load_s0_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : load_s0_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : load_s0_output_rData_roundMode_string = "RMM";
      default : load_s0_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(load_s0_output_rData_format)
      FpuFormat_FLOAT : load_s0_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : load_s0_output_rData_format_string = "DOUBLE";
      default : load_s0_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(load_s1_output_payload_roundMode)
      FpuRoundMode_RNE : load_s1_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : load_s1_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : load_s1_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : load_s1_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : load_s1_output_payload_roundMode_string = "RMM";
      default : load_s1_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(load_s1_output_payload_format)
      FpuFormat_FLOAT : load_s1_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : load_s1_output_payload_format_string = "DOUBLE";
      default : load_s1_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(shortPip_input_payload_opcode)
      FpuOpcode_LOAD : shortPip_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : shortPip_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : shortPip_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : shortPip_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : shortPip_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : shortPip_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : shortPip_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : shortPip_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : shortPip_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : shortPip_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : shortPip_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : shortPip_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : shortPip_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : shortPip_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : shortPip_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : shortPip_input_payload_opcode_string = "FCVT_X_X";
      default : shortPip_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(shortPip_input_payload_roundMode)
      FpuRoundMode_RNE : shortPip_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : shortPip_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : shortPip_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : shortPip_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : shortPip_input_payload_roundMode_string = "RMM";
      default : shortPip_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(shortPip_input_payload_format)
      FpuFormat_FLOAT : shortPip_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : shortPip_input_payload_format_string = "DOUBLE";
      default : shortPip_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_shortPip_rData_opcode)
      FpuOpcode_LOAD : decode_shortPip_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : decode_shortPip_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : decode_shortPip_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : decode_shortPip_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : decode_shortPip_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : decode_shortPip_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : decode_shortPip_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : decode_shortPip_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : decode_shortPip_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : decode_shortPip_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : decode_shortPip_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : decode_shortPip_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : decode_shortPip_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : decode_shortPip_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : decode_shortPip_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : decode_shortPip_rData_opcode_string = "FCVT_X_X";
      default : decode_shortPip_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_shortPip_rData_roundMode)
      FpuRoundMode_RNE : decode_shortPip_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_shortPip_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_shortPip_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_shortPip_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_shortPip_rData_roundMode_string = "RMM";
      default : decode_shortPip_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_shortPip_rData_format)
      FpuFormat_FLOAT : decode_shortPip_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_shortPip_rData_format_string = "DOUBLE";
      default : decode_shortPip_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(shortPip_rfOutput_payload_roundMode)
      FpuRoundMode_RNE : shortPip_rfOutput_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : shortPip_rfOutput_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : shortPip_rfOutput_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : shortPip_rfOutput_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : shortPip_rfOutput_payload_roundMode_string = "RMM";
      default : shortPip_rfOutput_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(shortPip_rfOutput_payload_format)
      FpuFormat_FLOAT : shortPip_rfOutput_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : shortPip_rfOutput_payload_format_string = "DOUBLE";
      default : shortPip_rfOutput_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(shortPip_output_payload_roundMode)
      FpuRoundMode_RNE : shortPip_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : shortPip_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : shortPip_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : shortPip_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : shortPip_output_payload_roundMode_string = "RMM";
      default : shortPip_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(shortPip_output_payload_format)
      FpuFormat_FLOAT : shortPip_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : shortPip_output_payload_format_string = "DOUBLE";
      default : shortPip_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_shortPip_rfOutput_payload_format)
      FpuFormat_FLOAT : _zz_shortPip_rfOutput_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_shortPip_rfOutput_payload_format_string = "DOUBLE";
      default : _zz_shortPip_rfOutput_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_preMul_input_payload_roundMode)
      FpuRoundMode_RNE : mul_preMul_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_preMul_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_preMul_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_preMul_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_preMul_input_payload_roundMode_string = "RMM";
      default : mul_preMul_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_preMul_input_payload_format)
      FpuFormat_FLOAT : mul_preMul_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_preMul_input_payload_format_string = "DOUBLE";
      default : mul_preMul_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_mul_rData_roundMode)
      FpuRoundMode_RNE : decode_mul_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_mul_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_mul_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_mul_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_mul_rData_roundMode_string = "RMM";
      default : decode_mul_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_mul_rData_format)
      FpuFormat_FLOAT : decode_mul_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_mul_rData_format_string = "DOUBLE";
      default : decode_mul_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_preMul_output_payload_roundMode)
      FpuRoundMode_RNE : mul_preMul_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_preMul_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_preMul_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_preMul_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_preMul_output_payload_roundMode_string = "RMM";
      default : mul_preMul_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_preMul_output_payload_format)
      FpuFormat_FLOAT : mul_preMul_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_preMul_output_payload_format_string = "DOUBLE";
      default : mul_preMul_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_mul_input_payload_roundMode)
      FpuRoundMode_RNE : mul_mul_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_mul_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_mul_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_mul_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_mul_input_payload_roundMode_string = "RMM";
      default : mul_mul_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_mul_input_payload_format)
      FpuFormat_FLOAT : mul_mul_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_mul_input_payload_format_string = "DOUBLE";
      default : mul_mul_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_preMul_output_rData_roundMode)
      FpuRoundMode_RNE : mul_preMul_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_preMul_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_preMul_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_preMul_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_preMul_output_rData_roundMode_string = "RMM";
      default : mul_preMul_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_preMul_output_rData_format)
      FpuFormat_FLOAT : mul_preMul_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_preMul_output_rData_format_string = "DOUBLE";
      default : mul_preMul_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_mul_output_payload_roundMode)
      FpuRoundMode_RNE : mul_mul_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_mul_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_mul_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_mul_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_mul_output_payload_roundMode_string = "RMM";
      default : mul_mul_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_mul_output_payload_format)
      FpuFormat_FLOAT : mul_mul_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_mul_output_payload_format_string = "DOUBLE";
      default : mul_mul_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_sum1_input_payload_roundMode)
      FpuRoundMode_RNE : mul_sum1_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_sum1_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_sum1_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_sum1_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_sum1_input_payload_roundMode_string = "RMM";
      default : mul_sum1_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_sum1_input_payload_format)
      FpuFormat_FLOAT : mul_sum1_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_sum1_input_payload_format_string = "DOUBLE";
      default : mul_sum1_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_mul_output_rData_roundMode)
      FpuRoundMode_RNE : mul_mul_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_mul_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_mul_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_mul_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_mul_output_rData_roundMode_string = "RMM";
      default : mul_mul_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_mul_output_rData_format)
      FpuFormat_FLOAT : mul_mul_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_mul_output_rData_format_string = "DOUBLE";
      default : mul_mul_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_sum1_output_payload_roundMode)
      FpuRoundMode_RNE : mul_sum1_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_sum1_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_sum1_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_sum1_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_sum1_output_payload_roundMode_string = "RMM";
      default : mul_sum1_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_sum1_output_payload_format)
      FpuFormat_FLOAT : mul_sum1_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_sum1_output_payload_format_string = "DOUBLE";
      default : mul_sum1_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_sum2_input_payload_roundMode)
      FpuRoundMode_RNE : mul_sum2_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_sum2_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_sum2_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_sum2_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_sum2_input_payload_roundMode_string = "RMM";
      default : mul_sum2_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_sum2_input_payload_format)
      FpuFormat_FLOAT : mul_sum2_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_sum2_input_payload_format_string = "DOUBLE";
      default : mul_sum2_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_sum1_output_rData_roundMode)
      FpuRoundMode_RNE : mul_sum1_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_sum1_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_sum1_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_sum1_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_sum1_output_rData_roundMode_string = "RMM";
      default : mul_sum1_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_sum1_output_rData_format)
      FpuFormat_FLOAT : mul_sum1_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_sum1_output_rData_format_string = "DOUBLE";
      default : mul_sum1_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_sum2_output_payload_roundMode)
      FpuRoundMode_RNE : mul_sum2_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_sum2_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_sum2_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_sum2_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_sum2_output_payload_roundMode_string = "RMM";
      default : mul_sum2_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_sum2_output_payload_format)
      FpuFormat_FLOAT : mul_sum2_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_sum2_output_payload_format_string = "DOUBLE";
      default : mul_sum2_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_norm_input_payload_roundMode)
      FpuRoundMode_RNE : mul_norm_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_norm_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_norm_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_norm_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_norm_input_payload_roundMode_string = "RMM";
      default : mul_norm_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_norm_input_payload_format)
      FpuFormat_FLOAT : mul_norm_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_norm_input_payload_format_string = "DOUBLE";
      default : mul_norm_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_sum2_output_rData_roundMode)
      FpuRoundMode_RNE : mul_sum2_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_sum2_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_sum2_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_sum2_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_sum2_output_rData_roundMode_string = "RMM";
      default : mul_sum2_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_sum2_output_rData_format)
      FpuFormat_FLOAT : mul_sum2_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_sum2_output_rData_format_string = "DOUBLE";
      default : mul_sum2_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_result_output_payload_roundMode)
      FpuRoundMode_RNE : mul_result_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_result_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_result_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_result_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_result_output_payload_roundMode_string = "RMM";
      default : mul_result_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_result_output_payload_format)
      FpuFormat_FLOAT : mul_result_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_result_output_payload_format_string = "DOUBLE";
      default : mul_result_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_result_mulToAdd_payload_roundMode)
      FpuRoundMode_RNE : mul_result_mulToAdd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_result_mulToAdd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_result_mulToAdd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_result_mulToAdd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_result_mulToAdd_payload_roundMode_string = "RMM";
      default : mul_result_mulToAdd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_result_mulToAdd_payload_format)
      FpuFormat_FLOAT : mul_result_mulToAdd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_result_mulToAdd_payload_format_string = "DOUBLE";
      default : mul_result_mulToAdd_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_result_mulToAdd_m2sPipe_payload_roundMode)
      FpuRoundMode_RNE : mul_result_mulToAdd_m2sPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_result_mulToAdd_m2sPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_result_mulToAdd_m2sPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_result_mulToAdd_m2sPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_result_mulToAdd_m2sPipe_payload_roundMode_string = "RMM";
      default : mul_result_mulToAdd_m2sPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_result_mulToAdd_m2sPipe_payload_format)
      FpuFormat_FLOAT : mul_result_mulToAdd_m2sPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_result_mulToAdd_m2sPipe_payload_format_string = "DOUBLE";
      default : mul_result_mulToAdd_m2sPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(mul_result_mulToAdd_rData_roundMode)
      FpuRoundMode_RNE : mul_result_mulToAdd_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : mul_result_mulToAdd_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : mul_result_mulToAdd_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : mul_result_mulToAdd_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : mul_result_mulToAdd_rData_roundMode_string = "RMM";
      default : mul_result_mulToAdd_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(mul_result_mulToAdd_rData_format)
      FpuFormat_FLOAT : mul_result_mulToAdd_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : mul_result_mulToAdd_rData_format_string = "DOUBLE";
      default : mul_result_mulToAdd_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(div_input_payload_roundMode)
      FpuRoundMode_RNE : div_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : div_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : div_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : div_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : div_input_payload_roundMode_string = "RMM";
      default : div_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(div_input_payload_format)
      FpuFormat_FLOAT : div_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : div_input_payload_format_string = "DOUBLE";
      default : div_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_div_rData_roundMode)
      FpuRoundMode_RNE : decode_div_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_div_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_div_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_div_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_div_rData_roundMode_string = "RMM";
      default : decode_div_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_div_rData_format)
      FpuFormat_FLOAT : decode_div_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_div_rData_format_string = "DOUBLE";
      default : decode_div_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(div_output_payload_roundMode)
      FpuRoundMode_RNE : div_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : div_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : div_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : div_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : div_output_payload_roundMode_string = "RMM";
      default : div_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(div_output_payload_format)
      FpuFormat_FLOAT : div_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : div_output_payload_format_string = "DOUBLE";
      default : div_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(sqrt_input_payload_roundMode)
      FpuRoundMode_RNE : sqrt_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : sqrt_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : sqrt_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : sqrt_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : sqrt_input_payload_roundMode_string = "RMM";
      default : sqrt_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(sqrt_input_payload_format)
      FpuFormat_FLOAT : sqrt_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : sqrt_input_payload_format_string = "DOUBLE";
      default : sqrt_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_sqrt_rData_roundMode)
      FpuRoundMode_RNE : decode_sqrt_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : decode_sqrt_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : decode_sqrt_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : decode_sqrt_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : decode_sqrt_rData_roundMode_string = "RMM";
      default : decode_sqrt_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_sqrt_rData_format)
      FpuFormat_FLOAT : decode_sqrt_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_sqrt_rData_format_string = "DOUBLE";
      default : decode_sqrt_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(sqrt_output_payload_roundMode)
      FpuRoundMode_RNE : sqrt_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : sqrt_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : sqrt_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : sqrt_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : sqrt_output_payload_roundMode_string = "RMM";
      default : sqrt_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(sqrt_output_payload_format)
      FpuFormat_FLOAT : sqrt_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : sqrt_output_payload_format_string = "DOUBLE";
      default : sqrt_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_preShifter_input_payload_roundMode)
      FpuRoundMode_RNE : add_preShifter_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_preShifter_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_preShifter_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_preShifter_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_preShifter_input_payload_roundMode_string = "RMM";
      default : add_preShifter_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_preShifter_input_payload_format)
      FpuFormat_FLOAT : add_preShifter_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_preShifter_input_payload_format_string = "DOUBLE";
      default : add_preShifter_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_preShifter_output_payload_roundMode)
      FpuRoundMode_RNE : add_preShifter_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_preShifter_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_preShifter_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_preShifter_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_preShifter_output_payload_roundMode_string = "RMM";
      default : add_preShifter_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_preShifter_output_payload_format)
      FpuFormat_FLOAT : add_preShifter_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_preShifter_output_payload_format_string = "DOUBLE";
      default : add_preShifter_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_shifter_input_payload_roundMode)
      FpuRoundMode_RNE : add_shifter_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_shifter_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_shifter_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_shifter_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_shifter_input_payload_roundMode_string = "RMM";
      default : add_shifter_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_shifter_input_payload_format)
      FpuFormat_FLOAT : add_shifter_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_shifter_input_payload_format_string = "DOUBLE";
      default : add_shifter_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_preShifter_output_rData_roundMode)
      FpuRoundMode_RNE : add_preShifter_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_preShifter_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_preShifter_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_preShifter_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_preShifter_output_rData_roundMode_string = "RMM";
      default : add_preShifter_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_preShifter_output_rData_format)
      FpuFormat_FLOAT : add_preShifter_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_preShifter_output_rData_format_string = "DOUBLE";
      default : add_preShifter_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_shifter_output_payload_roundMode)
      FpuRoundMode_RNE : add_shifter_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_shifter_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_shifter_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_shifter_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_shifter_output_payload_roundMode_string = "RMM";
      default : add_shifter_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_shifter_output_payload_format)
      FpuFormat_FLOAT : add_shifter_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_shifter_output_payload_format_string = "DOUBLE";
      default : add_shifter_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_math_input_payload_roundMode)
      FpuRoundMode_RNE : add_math_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_math_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_math_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_math_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_math_input_payload_roundMode_string = "RMM";
      default : add_math_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_math_input_payload_format)
      FpuFormat_FLOAT : add_math_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_math_input_payload_format_string = "DOUBLE";
      default : add_math_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_shifter_output_rData_roundMode)
      FpuRoundMode_RNE : add_shifter_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_shifter_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_shifter_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_shifter_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_shifter_output_rData_roundMode_string = "RMM";
      default : add_shifter_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_shifter_output_rData_format)
      FpuFormat_FLOAT : add_shifter_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_shifter_output_rData_format_string = "DOUBLE";
      default : add_shifter_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_math_output_payload_roundMode)
      FpuRoundMode_RNE : add_math_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_math_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_math_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_math_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_math_output_payload_roundMode_string = "RMM";
      default : add_math_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_math_output_payload_format)
      FpuFormat_FLOAT : add_math_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_math_output_payload_format_string = "DOUBLE";
      default : add_math_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_oh_input_payload_roundMode)
      FpuRoundMode_RNE : add_oh_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_oh_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_oh_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_oh_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_oh_input_payload_roundMode_string = "RMM";
      default : add_oh_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_oh_input_payload_format)
      FpuFormat_FLOAT : add_oh_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_oh_input_payload_format_string = "DOUBLE";
      default : add_oh_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_math_output_rData_roundMode)
      FpuRoundMode_RNE : add_math_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_math_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_math_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_math_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_math_output_rData_roundMode_string = "RMM";
      default : add_math_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_math_output_rData_format)
      FpuFormat_FLOAT : add_math_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_math_output_rData_format_string = "DOUBLE";
      default : add_math_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_oh_output_payload_roundMode)
      FpuRoundMode_RNE : add_oh_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_oh_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_oh_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_oh_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_oh_output_payload_roundMode_string = "RMM";
      default : add_oh_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_oh_output_payload_format)
      FpuFormat_FLOAT : add_oh_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_oh_output_payload_format_string = "DOUBLE";
      default : add_oh_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_norm_input_payload_roundMode)
      FpuRoundMode_RNE : add_norm_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_norm_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_norm_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_norm_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_norm_input_payload_roundMode_string = "RMM";
      default : add_norm_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_norm_input_payload_format)
      FpuFormat_FLOAT : add_norm_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_norm_input_payload_format_string = "DOUBLE";
      default : add_norm_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_oh_output_rData_roundMode)
      FpuRoundMode_RNE : add_oh_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_oh_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_oh_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_oh_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_oh_output_rData_roundMode_string = "RMM";
      default : add_oh_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_oh_output_rData_format)
      FpuFormat_FLOAT : add_oh_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_oh_output_rData_format_string = "DOUBLE";
      default : add_oh_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_norm_output_payload_roundMode)
      FpuRoundMode_RNE : add_norm_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_norm_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_norm_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_norm_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_norm_output_payload_roundMode_string = "RMM";
      default : add_norm_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_norm_output_payload_format)
      FpuFormat_FLOAT : add_norm_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_norm_output_payload_format_string = "DOUBLE";
      default : add_norm_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_result_input_payload_roundMode)
      FpuRoundMode_RNE : add_result_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_result_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_result_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_result_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_result_input_payload_roundMode_string = "RMM";
      default : add_result_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_result_input_payload_format)
      FpuFormat_FLOAT : add_result_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_result_input_payload_format_string = "DOUBLE";
      default : add_result_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(add_result_output_payload_roundMode)
      FpuRoundMode_RNE : add_result_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : add_result_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : add_result_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : add_result_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : add_result_output_payload_roundMode_string = "RMM";
      default : add_result_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(add_result_output_payload_format)
      FpuFormat_FLOAT : add_result_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : add_result_output_payload_format_string = "DOUBLE";
      default : add_result_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(load_s1_output_m2sPipe_payload_roundMode)
      FpuRoundMode_RNE : load_s1_output_m2sPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : load_s1_output_m2sPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : load_s1_output_m2sPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : load_s1_output_m2sPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : load_s1_output_m2sPipe_payload_roundMode_string = "RMM";
      default : load_s1_output_m2sPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(load_s1_output_m2sPipe_payload_format)
      FpuFormat_FLOAT : load_s1_output_m2sPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : load_s1_output_m2sPipe_payload_format_string = "DOUBLE";
      default : load_s1_output_m2sPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(load_s1_output_rData_roundMode)
      FpuRoundMode_RNE : load_s1_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : load_s1_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : load_s1_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : load_s1_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : load_s1_output_rData_roundMode_string = "RMM";
      default : load_s1_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(load_s1_output_rData_format)
      FpuFormat_FLOAT : load_s1_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : load_s1_output_rData_format_string = "DOUBLE";
      default : load_s1_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(shortPip_output_m2sPipe_payload_roundMode)
      FpuRoundMode_RNE : shortPip_output_m2sPipe_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : shortPip_output_m2sPipe_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : shortPip_output_m2sPipe_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : shortPip_output_m2sPipe_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : shortPip_output_m2sPipe_payload_roundMode_string = "RMM";
      default : shortPip_output_m2sPipe_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(shortPip_output_m2sPipe_payload_format)
      FpuFormat_FLOAT : shortPip_output_m2sPipe_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : shortPip_output_m2sPipe_payload_format_string = "DOUBLE";
      default : shortPip_output_m2sPipe_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(shortPip_output_rData_roundMode)
      FpuRoundMode_RNE : shortPip_output_rData_roundMode_string = "RNE";
      FpuRoundMode_RTZ : shortPip_output_rData_roundMode_string = "RTZ";
      FpuRoundMode_RDN : shortPip_output_rData_roundMode_string = "RDN";
      FpuRoundMode_RUP : shortPip_output_rData_roundMode_string = "RUP";
      FpuRoundMode_RMM : shortPip_output_rData_roundMode_string = "RMM";
      default : shortPip_output_rData_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(shortPip_output_rData_format)
      FpuFormat_FLOAT : shortPip_output_rData_format_string = "FLOAT ";
      FpuFormat_DOUBLE : shortPip_output_rData_format_string = "DOUBLE";
      default : shortPip_output_rData_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(streamArbiter_10_io_output_combStage_payload_roundMode)
      FpuRoundMode_RNE : streamArbiter_10_io_output_combStage_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : streamArbiter_10_io_output_combStage_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : streamArbiter_10_io_output_combStage_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : streamArbiter_10_io_output_combStage_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : streamArbiter_10_io_output_combStage_payload_roundMode_string = "RMM";
      default : streamArbiter_10_io_output_combStage_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(streamArbiter_10_io_output_combStage_payload_format)
      FpuFormat_FLOAT : streamArbiter_10_io_output_combStage_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : streamArbiter_10_io_output_combStage_payload_format_string = "DOUBLE";
      default : streamArbiter_10_io_output_combStage_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(merge_arbitrated_payload_roundMode)
      FpuRoundMode_RNE : merge_arbitrated_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : merge_arbitrated_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : merge_arbitrated_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : merge_arbitrated_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : merge_arbitrated_payload_roundMode_string = "RMM";
      default : merge_arbitrated_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(merge_arbitrated_payload_format)
      FpuFormat_FLOAT : merge_arbitrated_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : merge_arbitrated_payload_format_string = "DOUBLE";
      default : merge_arbitrated_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(roundFront_input_payload_roundMode)
      FpuRoundMode_RNE : roundFront_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : roundFront_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : roundFront_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : roundFront_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : roundFront_input_payload_roundMode_string = "RMM";
      default : roundFront_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(roundFront_input_payload_format)
      FpuFormat_FLOAT : roundFront_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : roundFront_input_payload_format_string = "DOUBLE";
      default : roundFront_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(roundFront_output_payload_roundMode)
      FpuRoundMode_RNE : roundFront_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : roundFront_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : roundFront_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : roundFront_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : roundFront_output_payload_roundMode_string = "RMM";
      default : roundFront_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(roundFront_output_payload_format)
      FpuFormat_FLOAT : roundFront_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : roundFront_output_payload_format_string = "DOUBLE";
      default : roundFront_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(roundBack_input_payload_roundMode)
      FpuRoundMode_RNE : roundBack_input_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : roundBack_input_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : roundBack_input_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : roundBack_input_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : roundBack_input_payload_roundMode_string = "RMM";
      default : roundBack_input_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(roundBack_input_payload_format)
      FpuFormat_FLOAT : roundBack_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : roundBack_input_payload_format_string = "DOUBLE";
      default : roundBack_input_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(roundBack_output_payload_format)
      FpuFormat_FLOAT : roundBack_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : roundBack_output_payload_format_string = "DOUBLE";
      default : roundBack_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(writeback_input_payload_format)
      FpuFormat_FLOAT : writeback_input_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : writeback_input_payload_format_string = "DOUBLE";
      default : writeback_input_payload_format_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    if(writeback_port_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    roundFront_discardCount_1 = roundFront_discardCount;
    if(when_FpuCore_l1551) begin
      roundFront_discardCount_1 = (roundFront_discardCount + 13'h001d);
    end
  end

  always @(*) begin
    add_shifter_yMantissa_6 = add_shifter_yMantissa_5;
    add_shifter_yMantissa_6 = (add_shifter_shiftBy[0] ? _zz_add_shifter_yMantissa_6 : add_shifter_yMantissa_5);
    if(add_shifter_passThrough) begin
      add_shifter_yMantissa_6 = 55'h0;
    end
  end

  always @(*) begin
    add_shifter_yMantissa_5 = add_shifter_yMantissa_4;
    add_shifter_yMantissa_5 = (add_shifter_shiftBy[1] ? _zz_add_shifter_yMantissa_5 : add_shifter_yMantissa_4);
  end

  always @(*) begin
    add_shifter_yMantissa_4 = add_shifter_yMantissa_3;
    add_shifter_yMantissa_4 = (add_shifter_shiftBy[2] ? _zz_add_shifter_yMantissa_4 : add_shifter_yMantissa_3);
  end

  always @(*) begin
    add_shifter_yMantissa_3 = add_shifter_yMantissa_2;
    add_shifter_yMantissa_3 = (add_shifter_shiftBy[3] ? _zz_add_shifter_yMantissa_3 : add_shifter_yMantissa_2);
  end

  always @(*) begin
    add_shifter_yMantissa_2 = add_shifter_yMantissa_1;
    add_shifter_yMantissa_2 = (add_shifter_shiftBy[4] ? _zz_add_shifter_yMantissa_2 : add_shifter_yMantissa_1);
  end

  always @(*) begin
    add_shifter_yMantissa_1 = add_shifter_yMantissa;
    add_shifter_yMantissa_1 = (add_shifter_shiftBy[5] ? _zz_add_shifter_yMantissa_1 : add_shifter_yMantissa);
  end

  always @(*) begin
    shortPip_fsm_shift_input_6 = shortPip_fsm_shift_input_5;
    shortPip_fsm_shift_input_6 = (shortPip_fsm_shift_by[0] ? _zz_shortPip_fsm_shift_input_6 : shortPip_fsm_shift_input_5);
  end

  always @(*) begin
    shortPip_fsm_shift_input_5 = shortPip_fsm_shift_input_4;
    shortPip_fsm_shift_input_5 = (shortPip_fsm_shift_by[1] ? _zz_shortPip_fsm_shift_input_5 : shortPip_fsm_shift_input_4);
  end

  always @(*) begin
    shortPip_fsm_shift_input_4 = shortPip_fsm_shift_input_3;
    shortPip_fsm_shift_input_4 = (shortPip_fsm_shift_by[2] ? _zz_shortPip_fsm_shift_input_4 : shortPip_fsm_shift_input_3);
  end

  always @(*) begin
    shortPip_fsm_shift_input_3 = shortPip_fsm_shift_input_2;
    shortPip_fsm_shift_input_3 = (shortPip_fsm_shift_by[3] ? _zz_shortPip_fsm_shift_input_3 : shortPip_fsm_shift_input_2);
  end

  always @(*) begin
    shortPip_fsm_shift_input_2 = shortPip_fsm_shift_input_1;
    shortPip_fsm_shift_input_2 = (shortPip_fsm_shift_by[4] ? _zz_shortPip_fsm_shift_input_2 : shortPip_fsm_shift_input_1);
  end

  always @(*) begin
    shortPip_fsm_shift_input_1 = shortPip_fsm_shift_input;
    shortPip_fsm_shift_input_1 = (shortPip_fsm_shift_by[5] ? _zz_shortPip_fsm_shift_input_1 : shortPip_fsm_shift_input);
  end

  always @(*) begin
    load_s1_fsm_shift_input_6 = load_s1_fsm_shift_input_5;
    load_s1_fsm_shift_input_6 = (load_s1_fsm_shift_by[5] ? _zz_load_s1_fsm_shift_input_6 : load_s1_fsm_shift_input_5);
  end

  always @(*) begin
    load_s1_fsm_shift_input_5 = load_s1_fsm_shift_input_4;
    load_s1_fsm_shift_input_5 = (load_s1_fsm_shift_by[4] ? _zz_load_s1_fsm_shift_input_5 : load_s1_fsm_shift_input_4);
  end

  always @(*) begin
    load_s1_fsm_shift_input_4 = load_s1_fsm_shift_input_3;
    load_s1_fsm_shift_input_4 = (load_s1_fsm_shift_by[3] ? _zz_load_s1_fsm_shift_input_4 : load_s1_fsm_shift_input_3);
  end

  always @(*) begin
    load_s1_fsm_shift_input_3 = load_s1_fsm_shift_input_2;
    load_s1_fsm_shift_input_3 = (load_s1_fsm_shift_by[2] ? _zz_load_s1_fsm_shift_input_3 : load_s1_fsm_shift_input_2);
  end

  always @(*) begin
    load_s1_fsm_shift_input_2 = load_s1_fsm_shift_input_1;
    load_s1_fsm_shift_input_2 = (load_s1_fsm_shift_by[1] ? _zz_load_s1_fsm_shift_input_2 : load_s1_fsm_shift_input_1);
  end

  always @(*) begin
    load_s1_fsm_shift_input_1 = load_s1_fsm_shift_input;
    load_s1_fsm_shift_input_1 = (load_s1_fsm_shift_by[0] ? _zz_load_s1_fsm_shift_input_1 : load_s1_fsm_shift_input);
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(commitLogic_1_input_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(commitLogic_0_input_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(rf_scoreboards_1_hitWrite_valid) begin
      _zz_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(rf_scoreboards_1_targetWrite_valid) begin
      _zz_5 = 1'b1;
    end
  end

  always @(*) begin
    _zz_6 = 1'b0;
    if(rf_scoreboards_0_hitWrite_valid) begin
      _zz_6 = 1'b1;
    end
  end

  always @(*) begin
    _zz_7 = 1'b0;
    if(rf_scoreboards_0_targetWrite_valid) begin
      _zz_7 = 1'b1;
    end
  end

  assign rf_init_done = rf_init_counter[5];
  assign when_FpuCore_l163 = (! rf_init_done);
  always @(*) begin
    rf_scoreboards_0_targetWrite_valid = (! rf_init_done);
    if(when_FpuCore_l265) begin
      rf_scoreboards_0_targetWrite_valid = 1'b1;
    end
  end

  always @(*) begin
    rf_scoreboards_0_targetWrite_payload_address = rf_init_counter[4:0];
    if(when_FpuCore_l261) begin
      rf_scoreboards_0_targetWrite_payload_address = scheduler_0_input_payload_rd;
    end
  end

  always @(*) begin
    rf_scoreboards_0_targetWrite_payload_data = 1'b0;
    if(when_FpuCore_l261) begin
      rf_scoreboards_0_targetWrite_payload_data = (! scheduler_0_rfTargets_3);
    end
  end

  always @(*) begin
    rf_scoreboards_0_hitWrite_valid = (! rf_init_done);
    if(writeback_input_valid) begin
      if(when_FpuCore_l1689) begin
        rf_scoreboards_0_hitWrite_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    rf_scoreboards_0_hitWrite_payload_address = rf_init_counter[4:0];
    if(writeback_input_valid) begin
      rf_scoreboards_0_hitWrite_payload_address = writeback_input_payload_rd;
    end
  end

  always @(*) begin
    rf_scoreboards_0_hitWrite_payload_data = 1'b0;
    if(writeback_input_valid) begin
      rf_scoreboards_0_hitWrite_payload_data = (! rf_scoreboards_0_hit_spinal_port5[0]);
    end
  end

  always @(*) begin
    rf_scoreboards_1_targetWrite_valid = (! rf_init_done);
    if(when_FpuCore_l265_1) begin
      rf_scoreboards_1_targetWrite_valid = 1'b1;
    end
  end

  always @(*) begin
    rf_scoreboards_1_targetWrite_payload_address = rf_init_counter[4:0];
    if(when_FpuCore_l261_1) begin
      rf_scoreboards_1_targetWrite_payload_address = scheduler_1_input_payload_rd;
    end
  end

  always @(*) begin
    rf_scoreboards_1_targetWrite_payload_data = 1'b0;
    if(when_FpuCore_l261_1) begin
      rf_scoreboards_1_targetWrite_payload_data = (! scheduler_1_rfTargets_3);
    end
  end

  always @(*) begin
    rf_scoreboards_1_hitWrite_valid = (! rf_init_done);
    if(writeback_input_valid) begin
      if(when_FpuCore_l1689_1) begin
        rf_scoreboards_1_hitWrite_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    rf_scoreboards_1_hitWrite_payload_address = rf_init_counter[4:0];
    if(writeback_input_valid) begin
      rf_scoreboards_1_hitWrite_payload_address = writeback_input_payload_rd;
    end
  end

  always @(*) begin
    rf_scoreboards_1_hitWrite_payload_data = 1'b0;
    if(writeback_input_valid) begin
      rf_scoreboards_1_hitWrite_payload_data = (! rf_scoreboards_1_hit_spinal_port5[0]);
    end
  end

  assign io_port_0_commit_ready = streamFork_3_io_input_ready;
  assign commitFork_load_0_valid = streamFork_3_io_outputs_0_valid;
  assign commitFork_load_0_payload_opcode = streamFork_3_io_outputs_0_payload_opcode;
  assign commitFork_load_0_payload_rd = streamFork_3_io_outputs_0_payload_rd;
  assign commitFork_load_0_payload_write = streamFork_3_io_outputs_0_payload_write;
  assign commitFork_load_0_payload_value = streamFork_3_io_outputs_0_payload_value;
  assign streamFork_3_io_outputs_1_s2mPipe_valid = (streamFork_3_io_outputs_1_valid || (! streamFork_3_io_outputs_1_rValidN));
  assign _zz_payload_opcode = (streamFork_3_io_outputs_1_rValidN ? streamFork_3_io_outputs_1_payload_opcode : streamFork_3_io_outputs_1_rData_opcode);
  assign streamFork_3_io_outputs_1_s2mPipe_payload_opcode = _zz_payload_opcode;
  assign streamFork_3_io_outputs_1_s2mPipe_payload_rd = (streamFork_3_io_outputs_1_rValidN ? streamFork_3_io_outputs_1_payload_rd : streamFork_3_io_outputs_1_rData_rd);
  assign streamFork_3_io_outputs_1_s2mPipe_payload_write = (streamFork_3_io_outputs_1_rValidN ? streamFork_3_io_outputs_1_payload_write : streamFork_3_io_outputs_1_rData_write);
  assign streamFork_3_io_outputs_1_s2mPipe_payload_value = (streamFork_3_io_outputs_1_rValidN ? streamFork_3_io_outputs_1_payload_value : streamFork_3_io_outputs_1_rData_value);
  assign commitFork_commit_0_valid = streamFork_3_io_outputs_1_s2mPipe_valid;
  assign streamFork_3_io_outputs_1_s2mPipe_ready = commitFork_commit_0_ready;
  assign commitFork_commit_0_payload_opcode = streamFork_3_io_outputs_1_s2mPipe_payload_opcode;
  assign commitFork_commit_0_payload_rd = streamFork_3_io_outputs_1_s2mPipe_payload_rd;
  assign commitFork_commit_0_payload_write = streamFork_3_io_outputs_1_s2mPipe_payload_write;
  assign commitFork_commit_0_payload_value = streamFork_3_io_outputs_1_s2mPipe_payload_value;
  assign io_port_1_commit_ready = streamFork_4_io_input_ready;
  assign commitFork_load_1_valid = streamFork_4_io_outputs_0_valid;
  assign commitFork_load_1_payload_opcode = streamFork_4_io_outputs_0_payload_opcode;
  assign commitFork_load_1_payload_rd = streamFork_4_io_outputs_0_payload_rd;
  assign commitFork_load_1_payload_write = streamFork_4_io_outputs_0_payload_write;
  assign commitFork_load_1_payload_value = streamFork_4_io_outputs_0_payload_value;
  assign streamFork_4_io_outputs_1_s2mPipe_valid = (streamFork_4_io_outputs_1_valid || (! streamFork_4_io_outputs_1_rValidN));
  assign _zz_payload_opcode_1 = (streamFork_4_io_outputs_1_rValidN ? streamFork_4_io_outputs_1_payload_opcode : streamFork_4_io_outputs_1_rData_opcode);
  assign streamFork_4_io_outputs_1_s2mPipe_payload_opcode = _zz_payload_opcode_1;
  assign streamFork_4_io_outputs_1_s2mPipe_payload_rd = (streamFork_4_io_outputs_1_rValidN ? streamFork_4_io_outputs_1_payload_rd : streamFork_4_io_outputs_1_rData_rd);
  assign streamFork_4_io_outputs_1_s2mPipe_payload_write = (streamFork_4_io_outputs_1_rValidN ? streamFork_4_io_outputs_1_payload_write : streamFork_4_io_outputs_1_rData_write);
  assign streamFork_4_io_outputs_1_s2mPipe_payload_value = (streamFork_4_io_outputs_1_rValidN ? streamFork_4_io_outputs_1_payload_value : streamFork_4_io_outputs_1_rData_value);
  assign commitFork_commit_1_valid = streamFork_4_io_outputs_1_s2mPipe_valid;
  assign streamFork_4_io_outputs_1_s2mPipe_ready = commitFork_commit_1_ready;
  assign commitFork_commit_1_payload_opcode = streamFork_4_io_outputs_1_s2mPipe_payload_opcode;
  assign commitFork_commit_1_payload_rd = streamFork_4_io_outputs_1_s2mPipe_payload_rd;
  assign commitFork_commit_1_payload_write = streamFork_4_io_outputs_1_s2mPipe_payload_write;
  assign commitFork_commit_1_payload_value = streamFork_4_io_outputs_1_s2mPipe_payload_value;
  assign commitLogic_0_pending_full = (&commitLogic_0_pending_counter);
  assign commitLogic_0_pending_notEmpty = (|commitLogic_0_pending_counter);
  always @(*) begin
    commitLogic_0_pending_inc = 1'b0;
    if(when_FpuCore_l265) begin
      commitLogic_0_pending_inc = 1'b1;
    end
  end

  always @(*) begin
    commitLogic_0_pending_dec = 1'b0;
    if(commitLogic_0_input_valid) begin
      commitLogic_0_pending_dec = 1'b1;
    end
  end

  assign commitLogic_0_add_full = (&commitLogic_0_add_counter);
  assign commitLogic_0_add_notEmpty = (|commitLogic_0_add_counter);
  always @(*) begin
    commitLogic_0_add_inc = 1'b0;
    if(commitLogic_0_input_valid) begin
      if(when_FpuCore_l208) begin
        commitLogic_0_add_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_0_add_dec = 1'b0;
    if(when_FpuCore_l221_8) begin
      commitLogic_0_add_dec = 1'b1;
    end
  end

  assign commitLogic_0_mul_full = (&commitLogic_0_mul_counter);
  assign commitLogic_0_mul_notEmpty = (|commitLogic_0_mul_counter);
  always @(*) begin
    commitLogic_0_mul_inc = 1'b0;
    if(commitLogic_0_input_valid) begin
      if(when_FpuCore_l209) begin
        commitLogic_0_mul_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_0_mul_dec = 1'b0;
    if(when_FpuCore_l221_2) begin
      commitLogic_0_mul_dec = 1'b1;
    end
  end

  assign commitLogic_0_div_full = (&commitLogic_0_div_counter);
  assign commitLogic_0_div_notEmpty = (|commitLogic_0_div_counter);
  always @(*) begin
    commitLogic_0_div_inc = 1'b0;
    if(commitLogic_0_input_valid) begin
      if(when_FpuCore_l210) begin
        commitLogic_0_div_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_0_div_dec = 1'b0;
    if(when_FpuCore_l221_4) begin
      commitLogic_0_div_dec = 1'b1;
    end
  end

  assign commitLogic_0_sqrt_full = (&commitLogic_0_sqrt_counter);
  assign commitLogic_0_sqrt_notEmpty = (|commitLogic_0_sqrt_counter);
  always @(*) begin
    commitLogic_0_sqrt_inc = 1'b0;
    if(commitLogic_0_input_valid) begin
      if(when_FpuCore_l211) begin
        commitLogic_0_sqrt_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_0_sqrt_dec = 1'b0;
    if(when_FpuCore_l221_6) begin
      commitLogic_0_sqrt_dec = 1'b1;
    end
  end

  assign commitLogic_0_short_full = (&commitLogic_0_short_counter);
  assign commitLogic_0_short_notEmpty = (|commitLogic_0_short_counter);
  always @(*) begin
    commitLogic_0_short_inc = 1'b0;
    if(commitLogic_0_input_valid) begin
      if(when_FpuCore_l212) begin
        commitLogic_0_short_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_0_short_dec = 1'b0;
    if(when_FpuCore_l221) begin
      commitLogic_0_short_dec = 1'b1;
    end
  end

  assign _zz_commitFork_commit_0_ready = (! ((|{commitLogic_0_short_full,{commitLogic_0_sqrt_full,{commitLogic_0_div_full,{commitLogic_0_mul_full,commitLogic_0_add_full}}}}) || (! commitLogic_0_pending_notEmpty)));
  assign commitFork_commit_0_ready = (1'b1 && _zz_commitFork_commit_0_ready);
  assign _zz_commitLogic_0_input_payload_opcode = commitFork_commit_0_payload_opcode;
  assign commitLogic_0_input_valid = (commitFork_commit_0_valid && _zz_commitFork_commit_0_ready);
  assign commitLogic_0_input_payload_opcode = _zz_commitLogic_0_input_payload_opcode;
  assign commitLogic_0_input_payload_rd = commitFork_commit_0_payload_rd;
  assign commitLogic_0_input_payload_write = commitFork_commit_0_payload_write;
  assign commitLogic_0_input_payload_value = commitFork_commit_0_payload_value;
  assign when_FpuCore_l208 = (|(commitLogic_0_input_payload_opcode == FpuOpcode_ADD));
  assign when_FpuCore_l209 = (|{(commitLogic_0_input_payload_opcode == FpuOpcode_FMA),(commitLogic_0_input_payload_opcode == FpuOpcode_MUL)});
  assign when_FpuCore_l210 = (|(commitLogic_0_input_payload_opcode == FpuOpcode_DIV));
  assign when_FpuCore_l211 = (|(commitLogic_0_input_payload_opcode == FpuOpcode_SQRT));
  assign when_FpuCore_l212 = (|{(commitLogic_0_input_payload_opcode == FpuOpcode_FCVT_X_X),{(commitLogic_0_input_payload_opcode == FpuOpcode_MIN_MAX),(commitLogic_0_input_payload_opcode == FpuOpcode_SGNJ)}});
  assign commitLogic_1_pending_full = (&commitLogic_1_pending_counter);
  assign commitLogic_1_pending_notEmpty = (|commitLogic_1_pending_counter);
  always @(*) begin
    commitLogic_1_pending_inc = 1'b0;
    if(when_FpuCore_l265_1) begin
      commitLogic_1_pending_inc = 1'b1;
    end
  end

  always @(*) begin
    commitLogic_1_pending_dec = 1'b0;
    if(commitLogic_1_input_valid) begin
      commitLogic_1_pending_dec = 1'b1;
    end
  end

  assign commitLogic_1_add_full = (&commitLogic_1_add_counter);
  assign commitLogic_1_add_notEmpty = (|commitLogic_1_add_counter);
  always @(*) begin
    commitLogic_1_add_inc = 1'b0;
    if(commitLogic_1_input_valid) begin
      if(when_FpuCore_l208_1) begin
        commitLogic_1_add_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_1_add_dec = 1'b0;
    if(when_FpuCore_l221_9) begin
      commitLogic_1_add_dec = 1'b1;
    end
  end

  assign commitLogic_1_mul_full = (&commitLogic_1_mul_counter);
  assign commitLogic_1_mul_notEmpty = (|commitLogic_1_mul_counter);
  always @(*) begin
    commitLogic_1_mul_inc = 1'b0;
    if(commitLogic_1_input_valid) begin
      if(when_FpuCore_l209_1) begin
        commitLogic_1_mul_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_1_mul_dec = 1'b0;
    if(when_FpuCore_l221_3) begin
      commitLogic_1_mul_dec = 1'b1;
    end
  end

  assign commitLogic_1_div_full = (&commitLogic_1_div_counter);
  assign commitLogic_1_div_notEmpty = (|commitLogic_1_div_counter);
  always @(*) begin
    commitLogic_1_div_inc = 1'b0;
    if(commitLogic_1_input_valid) begin
      if(when_FpuCore_l210_1) begin
        commitLogic_1_div_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_1_div_dec = 1'b0;
    if(when_FpuCore_l221_5) begin
      commitLogic_1_div_dec = 1'b1;
    end
  end

  assign commitLogic_1_sqrt_full = (&commitLogic_1_sqrt_counter);
  assign commitLogic_1_sqrt_notEmpty = (|commitLogic_1_sqrt_counter);
  always @(*) begin
    commitLogic_1_sqrt_inc = 1'b0;
    if(commitLogic_1_input_valid) begin
      if(when_FpuCore_l211_1) begin
        commitLogic_1_sqrt_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_1_sqrt_dec = 1'b0;
    if(when_FpuCore_l221_7) begin
      commitLogic_1_sqrt_dec = 1'b1;
    end
  end

  assign commitLogic_1_short_full = (&commitLogic_1_short_counter);
  assign commitLogic_1_short_notEmpty = (|commitLogic_1_short_counter);
  always @(*) begin
    commitLogic_1_short_inc = 1'b0;
    if(commitLogic_1_input_valid) begin
      if(when_FpuCore_l212_1) begin
        commitLogic_1_short_inc = 1'b1;
      end
    end
  end

  always @(*) begin
    commitLogic_1_short_dec = 1'b0;
    if(when_FpuCore_l221_1) begin
      commitLogic_1_short_dec = 1'b1;
    end
  end

  assign _zz_commitFork_commit_1_ready = (! ((|{commitLogic_1_short_full,{commitLogic_1_sqrt_full,{commitLogic_1_div_full,{commitLogic_1_mul_full,commitLogic_1_add_full}}}}) || (! commitLogic_1_pending_notEmpty)));
  assign commitFork_commit_1_ready = (1'b1 && _zz_commitFork_commit_1_ready);
  assign _zz_commitLogic_1_input_payload_opcode = commitFork_commit_1_payload_opcode;
  assign commitLogic_1_input_valid = (commitFork_commit_1_valid && _zz_commitFork_commit_1_ready);
  assign commitLogic_1_input_payload_opcode = _zz_commitLogic_1_input_payload_opcode;
  assign commitLogic_1_input_payload_rd = commitFork_commit_1_payload_rd;
  assign commitLogic_1_input_payload_write = commitFork_commit_1_payload_write;
  assign commitLogic_1_input_payload_value = commitFork_commit_1_payload_value;
  assign when_FpuCore_l208_1 = (|(commitLogic_1_input_payload_opcode == FpuOpcode_ADD));
  assign when_FpuCore_l209_1 = (|{(commitLogic_1_input_payload_opcode == FpuOpcode_FMA),(commitLogic_1_input_payload_opcode == FpuOpcode_MUL)});
  assign when_FpuCore_l210_1 = (|(commitLogic_1_input_payload_opcode == FpuOpcode_DIV));
  assign when_FpuCore_l211_1 = (|(commitLogic_1_input_payload_opcode == FpuOpcode_SQRT));
  assign when_FpuCore_l212_1 = (|{(commitLogic_1_input_payload_opcode == FpuOpcode_FCVT_X_X),{(commitLogic_1_input_payload_opcode == FpuOpcode_MIN_MAX),(commitLogic_1_input_payload_opcode == FpuOpcode_SGNJ)}});
  assign io_port_0_cmd_ready = io_port_0_cmd_rValidN;
  assign scheduler_0_input_valid = (io_port_0_cmd_valid || (! io_port_0_cmd_rValidN));
  assign _zz_scheduler_0_input_payload_opcode = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_opcode : io_port_0_cmd_rData_opcode);
  assign _zz_scheduler_0_input_payload_format = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_format : io_port_0_cmd_rData_format);
  assign _zz_scheduler_0_input_payload_roundMode = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_roundMode : io_port_0_cmd_rData_roundMode);
  assign scheduler_0_input_payload_opcode = _zz_scheduler_0_input_payload_opcode;
  assign scheduler_0_input_payload_arg = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_arg : io_port_0_cmd_rData_arg);
  assign scheduler_0_input_payload_rs1 = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_rs1 : io_port_0_cmd_rData_rs1);
  assign scheduler_0_input_payload_rs2 = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_rs2 : io_port_0_cmd_rData_rs2);
  assign scheduler_0_input_payload_rs3 = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_rs3 : io_port_0_cmd_rData_rs3);
  assign scheduler_0_input_payload_rd = (io_port_0_cmd_rValidN ? io_port_0_cmd_payload_rd : io_port_0_cmd_rData_rd);
  assign scheduler_0_input_payload_format = _zz_scheduler_0_input_payload_format;
  assign scheduler_0_input_payload_roundMode = _zz_scheduler_0_input_payload_roundMode;
  always @(*) begin
    scheduler_0_useRs1 = 1'b0;
    case(scheduler_0_input_payload_opcode)
      FpuOpcode_LOAD : begin
      end
      FpuOpcode_STORE : begin
      end
      FpuOpcode_ADD : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_MUL : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_DIV : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_SQRT : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_FMA : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_I2F : begin
      end
      FpuOpcode_F2I : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_MIN_MAX : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_CMP : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_SGNJ : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_FMV_X_W : begin
        scheduler_0_useRs1 = 1'b1;
      end
      FpuOpcode_FMV_W_X : begin
      end
      FpuOpcode_FCLASS : begin
        scheduler_0_useRs1 = 1'b1;
      end
      default : begin
        scheduler_0_useRs1 = 1'b1;
      end
    endcase
  end

  always @(*) begin
    scheduler_0_useRs2 = 1'b0;
    case(scheduler_0_input_payload_opcode)
      FpuOpcode_LOAD : begin
      end
      FpuOpcode_STORE : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_ADD : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_MUL : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_DIV : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_SQRT : begin
      end
      FpuOpcode_FMA : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_I2F : begin
      end
      FpuOpcode_F2I : begin
      end
      FpuOpcode_MIN_MAX : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_CMP : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_SGNJ : begin
        scheduler_0_useRs2 = 1'b1;
      end
      FpuOpcode_FMV_X_W : begin
      end
      FpuOpcode_FMV_W_X : begin
      end
      FpuOpcode_FCLASS : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    scheduler_0_useRs3 = 1'b0;
    case(scheduler_0_input_payload_opcode)
      FpuOpcode_LOAD : begin
      end
      FpuOpcode_STORE : begin
      end
      FpuOpcode_ADD : begin
      end
      FpuOpcode_MUL : begin
      end
      FpuOpcode_DIV : begin
      end
      FpuOpcode_SQRT : begin
      end
      FpuOpcode_FMA : begin
        scheduler_0_useRs3 = 1'b1;
      end
      FpuOpcode_I2F : begin
      end
      FpuOpcode_F2I : begin
      end
      FpuOpcode_MIN_MAX : begin
      end
      FpuOpcode_CMP : begin
      end
      FpuOpcode_SGNJ : begin
      end
      FpuOpcode_FMV_X_W : begin
      end
      FpuOpcode_FMV_W_X : begin
      end
      FpuOpcode_FCLASS : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    scheduler_0_useRd = 1'b0;
    case(scheduler_0_input_payload_opcode)
      FpuOpcode_LOAD : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_STORE : begin
      end
      FpuOpcode_ADD : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_MUL : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_DIV : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_SQRT : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_FMA : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_I2F : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_F2I : begin
      end
      FpuOpcode_MIN_MAX : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_CMP : begin
      end
      FpuOpcode_SGNJ : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_FMV_X_W : begin
      end
      FpuOpcode_FMV_W_X : begin
        scheduler_0_useRd = 1'b1;
      end
      FpuOpcode_FCLASS : begin
      end
      default : begin
        scheduler_0_useRd = 1'b1;
      end
    endcase
  end

  assign scheduler_0_rfHits_0 = rf_scoreboards_0_hit_spinal_port1[0];
  assign scheduler_0_rfHits_1 = rf_scoreboards_0_hit_spinal_port2[0];
  assign scheduler_0_rfHits_2 = rf_scoreboards_0_hit_spinal_port3[0];
  assign scheduler_0_rfHits_3 = rf_scoreboards_0_hit_spinal_port4[0];
  assign scheduler_0_rfTargets_0 = rf_scoreboards_0_target_spinal_port1[0];
  assign scheduler_0_rfTargets_1 = rf_scoreboards_0_target_spinal_port2[0];
  assign scheduler_0_rfTargets_2 = rf_scoreboards_0_target_spinal_port3[0];
  assign scheduler_0_rfTargets_3 = rf_scoreboards_0_target_spinal_port4[0];
  assign scheduler_0_rfBusy_0 = (scheduler_0_rfHits_0 ^ scheduler_0_rfTargets_0);
  assign scheduler_0_rfBusy_1 = (scheduler_0_rfHits_1 ^ scheduler_0_rfTargets_1);
  assign scheduler_0_rfBusy_2 = (scheduler_0_rfHits_2 ^ scheduler_0_rfTargets_2);
  assign scheduler_0_rfBusy_3 = (scheduler_0_rfHits_3 ^ scheduler_0_rfTargets_3);
  assign scheduler_0_hits_0 = (scheduler_0_useRs1 && scheduler_0_rfBusy_0);
  assign scheduler_0_hits_1 = (scheduler_0_useRs2 && scheduler_0_rfBusy_1);
  assign scheduler_0_hits_2 = (scheduler_0_useRs3 && scheduler_0_rfBusy_2);
  assign scheduler_0_hits_3 = (scheduler_0_useRd && scheduler_0_rfBusy_3);
  assign scheduler_0_hazard = (((|{scheduler_0_hits_3,{scheduler_0_hits_2,{scheduler_0_hits_1,scheduler_0_hits_0}}}) || (! rf_init_done)) || commitLogic_0_pending_full);
  assign _zz_scheduler_0_input_ready = (! scheduler_0_hazard);
  assign scheduler_0_output_valid = (scheduler_0_input_valid && _zz_scheduler_0_input_ready);
  assign scheduler_0_input_ready = (scheduler_0_output_ready && _zz_scheduler_0_input_ready);
  assign scheduler_0_output_payload_opcode = scheduler_0_input_payload_opcode;
  assign scheduler_0_output_payload_arg = scheduler_0_input_payload_arg;
  always @(*) begin
    scheduler_0_output_payload_rs1 = scheduler_0_input_payload_rs1;
    if(when_FpuCore_l258) begin
      scheduler_0_output_payload_rs1 = scheduler_0_input_payload_rs2;
    end
  end

  assign scheduler_0_output_payload_rs2 = scheduler_0_input_payload_rs2;
  assign scheduler_0_output_payload_rs3 = scheduler_0_input_payload_rs3;
  assign scheduler_0_output_payload_rd = scheduler_0_input_payload_rd;
  assign scheduler_0_output_payload_format = scheduler_0_input_payload_format;
  assign scheduler_0_output_payload_roundMode = scheduler_0_input_payload_roundMode;
  assign when_FpuCore_l258 = (scheduler_0_input_payload_opcode == FpuOpcode_STORE);
  assign when_FpuCore_l261 = (scheduler_0_input_valid && rf_init_done);
  assign scheduler_0_output_fire = (scheduler_0_output_valid && scheduler_0_output_ready);
  assign when_FpuCore_l265 = (scheduler_0_output_fire && scheduler_0_useRd);
  assign io_port_1_cmd_ready = io_port_1_cmd_rValidN;
  assign scheduler_1_input_valid = (io_port_1_cmd_valid || (! io_port_1_cmd_rValidN));
  assign _zz_scheduler_1_input_payload_opcode = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_opcode : io_port_1_cmd_rData_opcode);
  assign _zz_scheduler_1_input_payload_format = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_format : io_port_1_cmd_rData_format);
  assign _zz_scheduler_1_input_payload_roundMode = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_roundMode : io_port_1_cmd_rData_roundMode);
  assign scheduler_1_input_payload_opcode = _zz_scheduler_1_input_payload_opcode;
  assign scheduler_1_input_payload_arg = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_arg : io_port_1_cmd_rData_arg);
  assign scheduler_1_input_payload_rs1 = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_rs1 : io_port_1_cmd_rData_rs1);
  assign scheduler_1_input_payload_rs2 = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_rs2 : io_port_1_cmd_rData_rs2);
  assign scheduler_1_input_payload_rs3 = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_rs3 : io_port_1_cmd_rData_rs3);
  assign scheduler_1_input_payload_rd = (io_port_1_cmd_rValidN ? io_port_1_cmd_payload_rd : io_port_1_cmd_rData_rd);
  assign scheduler_1_input_payload_format = _zz_scheduler_1_input_payload_format;
  assign scheduler_1_input_payload_roundMode = _zz_scheduler_1_input_payload_roundMode;
  always @(*) begin
    scheduler_1_useRs1 = 1'b0;
    case(scheduler_1_input_payload_opcode)
      FpuOpcode_LOAD : begin
      end
      FpuOpcode_STORE : begin
      end
      FpuOpcode_ADD : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_MUL : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_DIV : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_SQRT : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_FMA : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_I2F : begin
      end
      FpuOpcode_F2I : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_MIN_MAX : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_CMP : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_SGNJ : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_FMV_X_W : begin
        scheduler_1_useRs1 = 1'b1;
      end
      FpuOpcode_FMV_W_X : begin
      end
      FpuOpcode_FCLASS : begin
        scheduler_1_useRs1 = 1'b1;
      end
      default : begin
        scheduler_1_useRs1 = 1'b1;
      end
    endcase
  end

  always @(*) begin
    scheduler_1_useRs2 = 1'b0;
    case(scheduler_1_input_payload_opcode)
      FpuOpcode_LOAD : begin
      end
      FpuOpcode_STORE : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_ADD : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_MUL : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_DIV : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_SQRT : begin
      end
      FpuOpcode_FMA : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_I2F : begin
      end
      FpuOpcode_F2I : begin
      end
      FpuOpcode_MIN_MAX : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_CMP : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_SGNJ : begin
        scheduler_1_useRs2 = 1'b1;
      end
      FpuOpcode_FMV_X_W : begin
      end
      FpuOpcode_FMV_W_X : begin
      end
      FpuOpcode_FCLASS : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    scheduler_1_useRs3 = 1'b0;
    case(scheduler_1_input_payload_opcode)
      FpuOpcode_LOAD : begin
      end
      FpuOpcode_STORE : begin
      end
      FpuOpcode_ADD : begin
      end
      FpuOpcode_MUL : begin
      end
      FpuOpcode_DIV : begin
      end
      FpuOpcode_SQRT : begin
      end
      FpuOpcode_FMA : begin
        scheduler_1_useRs3 = 1'b1;
      end
      FpuOpcode_I2F : begin
      end
      FpuOpcode_F2I : begin
      end
      FpuOpcode_MIN_MAX : begin
      end
      FpuOpcode_CMP : begin
      end
      FpuOpcode_SGNJ : begin
      end
      FpuOpcode_FMV_X_W : begin
      end
      FpuOpcode_FMV_W_X : begin
      end
      FpuOpcode_FCLASS : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    scheduler_1_useRd = 1'b0;
    case(scheduler_1_input_payload_opcode)
      FpuOpcode_LOAD : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_STORE : begin
      end
      FpuOpcode_ADD : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_MUL : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_DIV : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_SQRT : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_FMA : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_I2F : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_F2I : begin
      end
      FpuOpcode_MIN_MAX : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_CMP : begin
      end
      FpuOpcode_SGNJ : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_FMV_X_W : begin
      end
      FpuOpcode_FMV_W_X : begin
        scheduler_1_useRd = 1'b1;
      end
      FpuOpcode_FCLASS : begin
      end
      default : begin
        scheduler_1_useRd = 1'b1;
      end
    endcase
  end

  assign scheduler_1_rfHits_0 = rf_scoreboards_1_hit_spinal_port1[0];
  assign scheduler_1_rfHits_1 = rf_scoreboards_1_hit_spinal_port2[0];
  assign scheduler_1_rfHits_2 = rf_scoreboards_1_hit_spinal_port3[0];
  assign scheduler_1_rfHits_3 = rf_scoreboards_1_hit_spinal_port4[0];
  assign scheduler_1_rfTargets_0 = rf_scoreboards_1_target_spinal_port1[0];
  assign scheduler_1_rfTargets_1 = rf_scoreboards_1_target_spinal_port2[0];
  assign scheduler_1_rfTargets_2 = rf_scoreboards_1_target_spinal_port3[0];
  assign scheduler_1_rfTargets_3 = rf_scoreboards_1_target_spinal_port4[0];
  assign scheduler_1_rfBusy_0 = (scheduler_1_rfHits_0 ^ scheduler_1_rfTargets_0);
  assign scheduler_1_rfBusy_1 = (scheduler_1_rfHits_1 ^ scheduler_1_rfTargets_1);
  assign scheduler_1_rfBusy_2 = (scheduler_1_rfHits_2 ^ scheduler_1_rfTargets_2);
  assign scheduler_1_rfBusy_3 = (scheduler_1_rfHits_3 ^ scheduler_1_rfTargets_3);
  assign scheduler_1_hits_0 = (scheduler_1_useRs1 && scheduler_1_rfBusy_0);
  assign scheduler_1_hits_1 = (scheduler_1_useRs2 && scheduler_1_rfBusy_1);
  assign scheduler_1_hits_2 = (scheduler_1_useRs3 && scheduler_1_rfBusy_2);
  assign scheduler_1_hits_3 = (scheduler_1_useRd && scheduler_1_rfBusy_3);
  assign scheduler_1_hazard = (((|{scheduler_1_hits_3,{scheduler_1_hits_2,{scheduler_1_hits_1,scheduler_1_hits_0}}}) || (! rf_init_done)) || commitLogic_1_pending_full);
  assign _zz_scheduler_1_input_ready = (! scheduler_1_hazard);
  assign scheduler_1_output_valid = (scheduler_1_input_valid && _zz_scheduler_1_input_ready);
  assign scheduler_1_input_ready = (scheduler_1_output_ready && _zz_scheduler_1_input_ready);
  assign scheduler_1_output_payload_opcode = scheduler_1_input_payload_opcode;
  assign scheduler_1_output_payload_arg = scheduler_1_input_payload_arg;
  always @(*) begin
    scheduler_1_output_payload_rs1 = scheduler_1_input_payload_rs1;
    if(when_FpuCore_l258_1) begin
      scheduler_1_output_payload_rs1 = scheduler_1_input_payload_rs2;
    end
  end

  assign scheduler_1_output_payload_rs2 = scheduler_1_input_payload_rs2;
  assign scheduler_1_output_payload_rs3 = scheduler_1_input_payload_rs3;
  assign scheduler_1_output_payload_rd = scheduler_1_input_payload_rd;
  assign scheduler_1_output_payload_format = scheduler_1_input_payload_format;
  assign scheduler_1_output_payload_roundMode = scheduler_1_input_payload_roundMode;
  assign when_FpuCore_l258_1 = (scheduler_1_input_payload_opcode == FpuOpcode_STORE);
  assign when_FpuCore_l261_1 = (scheduler_1_input_valid && rf_init_done);
  assign scheduler_1_output_fire = (scheduler_1_output_valid && scheduler_1_output_ready);
  assign when_FpuCore_l265_1 = (scheduler_1_output_fire && scheduler_1_useRd);
  always @(*) begin
    scheduler_0_output_ready = scheduler_0_output_m2sPipe_ready;
    if(when_Stream_l375) begin
      scheduler_0_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! scheduler_0_output_m2sPipe_valid);
  assign scheduler_0_output_m2sPipe_valid = scheduler_0_output_rValid;
  assign scheduler_0_output_m2sPipe_payload_opcode = scheduler_0_output_rData_opcode;
  assign scheduler_0_output_m2sPipe_payload_arg = scheduler_0_output_rData_arg;
  assign scheduler_0_output_m2sPipe_payload_rs1 = scheduler_0_output_rData_rs1;
  assign scheduler_0_output_m2sPipe_payload_rs2 = scheduler_0_output_rData_rs2;
  assign scheduler_0_output_m2sPipe_payload_rs3 = scheduler_0_output_rData_rs3;
  assign scheduler_0_output_m2sPipe_payload_rd = scheduler_0_output_rData_rd;
  assign scheduler_0_output_m2sPipe_payload_format = scheduler_0_output_rData_format;
  assign scheduler_0_output_m2sPipe_payload_roundMode = scheduler_0_output_rData_roundMode;
  always @(*) begin
    scheduler_1_output_ready = scheduler_1_output_m2sPipe_ready;
    if(when_Stream_l375_1) begin
      scheduler_1_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! scheduler_1_output_m2sPipe_valid);
  assign scheduler_1_output_m2sPipe_valid = scheduler_1_output_rValid;
  assign scheduler_1_output_m2sPipe_payload_opcode = scheduler_1_output_rData_opcode;
  assign scheduler_1_output_m2sPipe_payload_arg = scheduler_1_output_rData_arg;
  assign scheduler_1_output_m2sPipe_payload_rs1 = scheduler_1_output_rData_rs1;
  assign scheduler_1_output_m2sPipe_payload_rs2 = scheduler_1_output_rData_rs2;
  assign scheduler_1_output_m2sPipe_payload_rs3 = scheduler_1_output_rData_rs3;
  assign scheduler_1_output_m2sPipe_payload_rd = scheduler_1_output_rData_rd;
  assign scheduler_1_output_m2sPipe_payload_format = scheduler_1_output_rData_format;
  assign scheduler_1_output_m2sPipe_payload_roundMode = scheduler_1_output_rData_roundMode;
  assign scheduler_0_output_m2sPipe_ready = cmdArbiter_arbiter_io_inputs_0_ready;
  assign scheduler_1_output_m2sPipe_ready = cmdArbiter_arbiter_io_inputs_1_ready;
  assign cmdArbiter_output_valid = cmdArbiter_arbiter_io_output_valid;
  assign cmdArbiter_output_payload_source = cmdArbiter_arbiter_io_chosen;
  assign cmdArbiter_output_payload_opcode = cmdArbiter_arbiter_io_output_payload_opcode;
  assign cmdArbiter_output_payload_rs1 = cmdArbiter_arbiter_io_output_payload_rs1;
  assign cmdArbiter_output_payload_rs2 = cmdArbiter_arbiter_io_output_payload_rs2;
  assign cmdArbiter_output_payload_rs3 = cmdArbiter_arbiter_io_output_payload_rs3;
  assign cmdArbiter_output_payload_rd = cmdArbiter_arbiter_io_output_payload_rd;
  assign cmdArbiter_output_payload_arg = cmdArbiter_arbiter_io_output_payload_arg;
  assign cmdArbiter_output_payload_roundMode = cmdArbiter_arbiter_io_output_payload_roundMode;
  assign cmdArbiter_output_payload_format = cmdArbiter_arbiter_io_output_payload_format;
  assign read_s0_valid = cmdArbiter_output_valid;
  assign cmdArbiter_output_ready = read_s0_ready;
  assign read_s0_payload_source = cmdArbiter_output_payload_source;
  assign read_s0_payload_opcode = cmdArbiter_output_payload_opcode;
  assign read_s0_payload_rs1 = cmdArbiter_output_payload_rs1;
  assign read_s0_payload_rs2 = cmdArbiter_output_payload_rs2;
  assign read_s0_payload_rs3 = cmdArbiter_output_payload_rs3;
  assign read_s0_payload_rd = cmdArbiter_output_payload_rd;
  assign read_s0_payload_arg = cmdArbiter_output_payload_arg;
  assign read_s0_payload_roundMode = cmdArbiter_output_payload_roundMode;
  assign read_s0_payload_format = cmdArbiter_output_payload_format;
  always @(*) begin
    read_s0_ready = read_s1_ready;
    if(when_Stream_l375_2) begin
      read_s0_ready = 1'b1;
    end
  end

  assign when_Stream_l375_2 = (! read_s1_valid);
  assign read_s1_valid = read_s0_rValid;
  assign read_s1_payload_source = read_s0_rData_source;
  assign read_s1_payload_opcode = read_s0_rData_opcode;
  assign read_s1_payload_rs1 = read_s0_rData_rs1;
  assign read_s1_payload_rs2 = read_s0_rData_rs2;
  assign read_s1_payload_rs3 = read_s0_rData_rs3;
  assign read_s1_payload_rd = read_s0_rData_rd;
  assign read_s1_payload_arg = read_s0_rData_arg;
  assign read_s1_payload_roundMode = read_s0_rData_roundMode;
  assign read_s1_payload_format = read_s0_rData_format;
  assign read_output_valid = read_s1_valid;
  assign read_s1_ready = read_output_ready;
  assign _zz_read_rs_0_boxed = {read_s0_payload_source,read_s0_payload_rs1};
  assign read_output_isStall = (read_output_valid && (! read_output_ready));
  assign _zz_read_rs_0_boxed_1 = (! read_output_isStall);
  assign _zz_read_rs_0_boxed_2 = rf_ram_spinal_port0;
  assign _zz_read_rs_0_value_mantissa = _zz_read_rs_0_boxed_2[65 : 0];
  assign read_rs_0_value_mantissa = _zz_read_rs_0_value_mantissa[51 : 0];
  assign read_rs_0_value_exponent = _zz_read_rs_0_value_mantissa[63 : 52];
  assign read_rs_0_value_sign = _zz_read_rs_0_value_mantissa[64];
  assign read_rs_0_value_special = _zz_read_rs_0_value_mantissa[65];
  assign read_rs_0_boxed = _zz_read_rs_0_boxed_2[66];
  assign _zz_read_rs_1_boxed = {read_s0_payload_source,read_s0_payload_rs2};
  assign _zz_read_rs_1_boxed_1 = (! read_output_isStall);
  assign _zz_read_rs_1_boxed_2 = rf_ram_spinal_port1;
  assign _zz_read_rs_1_value_mantissa = _zz_read_rs_1_boxed_2[65 : 0];
  assign read_rs_1_value_mantissa = _zz_read_rs_1_value_mantissa[51 : 0];
  assign read_rs_1_value_exponent = _zz_read_rs_1_value_mantissa[63 : 52];
  assign read_rs_1_value_sign = _zz_read_rs_1_value_mantissa[64];
  assign read_rs_1_value_special = _zz_read_rs_1_value_mantissa[65];
  assign read_rs_1_boxed = _zz_read_rs_1_boxed_2[66];
  assign _zz_read_rs_2_boxed = {read_s0_payload_source,read_s0_payload_rs3};
  assign _zz_read_rs_2_boxed_1 = (! read_output_isStall);
  assign _zz_read_rs_2_boxed_2 = rf_ram_spinal_port2;
  assign _zz_read_rs_2_value_mantissa = _zz_read_rs_2_boxed_2[65 : 0];
  assign read_rs_2_value_mantissa = _zz_read_rs_2_value_mantissa[51 : 0];
  assign read_rs_2_value_exponent = _zz_read_rs_2_value_mantissa[63 : 52];
  assign read_rs_2_value_sign = _zz_read_rs_2_value_mantissa[64];
  assign read_rs_2_value_special = _zz_read_rs_2_value_mantissa[65];
  assign read_rs_2_boxed = _zz_read_rs_2_boxed_2[66];
  assign read_output_payload_source = read_s1_payload_source;
  assign read_output_payload_opcode = read_s1_payload_opcode;
  assign read_output_payload_arg = read_s1_payload_arg;
  assign read_output_payload_roundMode = read_s1_payload_roundMode;
  assign read_output_payload_rd = read_s1_payload_rd;
  always @(*) begin
    read_output_payload_rs1_mantissa = read_rs_0_value_mantissa;
    if(when_FpuCore_l304) begin
      if(!when_FpuCore_l305) begin
        if(when_FpuCore_l307) begin
          read_output_payload_rs1_mantissa[51] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    read_output_payload_rs1_exponent = read_rs_0_value_exponent;
    if(when_FpuCore_l304) begin
      if(!when_FpuCore_l305) begin
        if(when_FpuCore_l307) begin
          read_output_payload_rs1_exponent[1 : 0] = 2'b10;
          read_output_payload_rs1_exponent[2] = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    read_output_payload_rs1_sign = read_rs_0_value_sign;
    if(when_FpuCore_l304) begin
      if(!when_FpuCore_l305) begin
        if(when_FpuCore_l307) begin
          read_output_payload_rs1_sign = 1'b0;
        end
      end
    end
  end

  always @(*) begin
    read_output_payload_rs1_special = read_rs_0_value_special;
    if(when_FpuCore_l304) begin
      if(!when_FpuCore_l305) begin
        if(when_FpuCore_l307) begin
          read_output_payload_rs1_special = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    read_output_payload_rs2_mantissa = read_rs_1_value_mantissa;
    if(when_FpuCore_l312) begin
      read_output_payload_rs2_mantissa[51] = 1'b1;
    end
  end

  always @(*) begin
    read_output_payload_rs2_exponent = read_rs_1_value_exponent;
    if(when_FpuCore_l312) begin
      read_output_payload_rs2_exponent[1 : 0] = 2'b10;
      read_output_payload_rs2_exponent[2] = 1'b1;
    end
  end

  always @(*) begin
    read_output_payload_rs2_sign = read_rs_1_value_sign;
    if(when_FpuCore_l312) begin
      read_output_payload_rs2_sign = 1'b0;
    end
  end

  always @(*) begin
    read_output_payload_rs2_special = read_rs_1_value_special;
    if(when_FpuCore_l312) begin
      read_output_payload_rs2_special = 1'b1;
    end
  end

  always @(*) begin
    read_output_payload_rs3_mantissa = read_rs_2_value_mantissa;
    if(when_FpuCore_l316) begin
      read_output_payload_rs3_mantissa[51] = 1'b1;
    end
  end

  always @(*) begin
    read_output_payload_rs3_exponent = read_rs_2_value_exponent;
    if(when_FpuCore_l316) begin
      read_output_payload_rs3_exponent[1 : 0] = 2'b10;
      read_output_payload_rs3_exponent[2] = 1'b1;
    end
  end

  assign read_output_payload_rs3_sign = read_rs_2_value_sign;
  always @(*) begin
    read_output_payload_rs3_special = read_rs_2_value_special;
    if(when_FpuCore_l316) begin
      read_output_payload_rs3_special = 1'b1;
    end
  end

  assign read_output_payload_rs1Boxed = read_rs_0_boxed;
  assign read_output_payload_rs2Boxed = read_rs_1_boxed;
  always @(*) begin
    read_output_payload_format = read_s1_payload_format;
    if(when_FpuCore_l304) begin
      if(when_FpuCore_l305) begin
        read_output_payload_format = _zz_read_output_payload_format;
      end
    end
  end

  assign when_FpuCore_l305 = ((read_s1_payload_opcode == FpuOpcode_STORE) || (read_s1_payload_opcode == FpuOpcode_FMV_X_W));
  assign when_FpuCore_l304 = (! ((read_s1_payload_opcode == FpuOpcode_SGNJ) && (read_s1_payload_format == FpuFormat_DOUBLE)));
  assign _zz_read_output_payload_format = (read_rs_0_boxed ? FpuFormat_FLOAT : FpuFormat_DOUBLE);
  assign when_FpuCore_l307 = ((read_s1_payload_format == FpuFormat_FLOAT) != read_rs_0_boxed);
  assign when_FpuCore_l312 = ((read_s1_payload_format == FpuFormat_FLOAT) != read_rs_1_boxed);
  assign when_FpuCore_l316 = ((read_s1_payload_format == FpuFormat_FLOAT) != read_rs_2_boxed);
  assign decode_input_valid = read_output_valid;
  assign read_output_ready = decode_input_ready;
  assign decode_input_payload_source = read_output_payload_source;
  assign decode_input_payload_opcode = read_output_payload_opcode;
  assign decode_input_payload_rs1_mantissa = read_output_payload_rs1_mantissa;
  assign decode_input_payload_rs1_exponent = read_output_payload_rs1_exponent;
  assign decode_input_payload_rs1_sign = read_output_payload_rs1_sign;
  assign decode_input_payload_rs1_special = read_output_payload_rs1_special;
  assign decode_input_payload_rs2_mantissa = read_output_payload_rs2_mantissa;
  assign decode_input_payload_rs2_exponent = read_output_payload_rs2_exponent;
  assign decode_input_payload_rs2_sign = read_output_payload_rs2_sign;
  assign decode_input_payload_rs2_special = read_output_payload_rs2_special;
  assign decode_input_payload_rs3_mantissa = read_output_payload_rs3_mantissa;
  assign decode_input_payload_rs3_exponent = read_output_payload_rs3_exponent;
  assign decode_input_payload_rs3_sign = read_output_payload_rs3_sign;
  assign decode_input_payload_rs3_special = read_output_payload_rs3_special;
  assign decode_input_payload_rd = read_output_payload_rd;
  assign decode_input_payload_arg = read_output_payload_arg;
  assign decode_input_payload_roundMode = read_output_payload_roundMode;
  assign decode_input_payload_format = read_output_payload_format;
  assign decode_input_payload_rs1Boxed = read_output_payload_rs1Boxed;
  assign decode_input_payload_rs2Boxed = read_output_payload_rs2Boxed;
  always @(*) begin
    decode_input_ready = 1'b0;
    if(when_FpuCore_l329) begin
      decode_input_ready = 1'b1;
    end
    if(when_FpuCore_l335) begin
      decode_input_ready = 1'b1;
    end
    if(when_FpuCore_l351) begin
      decode_input_ready = 1'b1;
    end
    if(when_FpuCore_l359) begin
      decode_input_ready = 1'b1;
    end
    if(when_FpuCore_l375) begin
      decode_input_ready = 1'b1;
    end
    if(when_FpuCore_l399) begin
      decode_input_ready = 1'b1;
    end
  end

  assign decode_loadHit = (|{(decode_input_payload_opcode == FpuOpcode_I2F),{(decode_input_payload_opcode == FpuOpcode_FMV_W_X),(decode_input_payload_opcode == FpuOpcode_LOAD)}});
  assign decode_load_valid = (decode_input_valid && decode_loadHit);
  assign when_FpuCore_l329 = (decode_loadHit && decode_load_ready);
  assign decode_load_payload_source = decode_input_payload_source;
  assign decode_load_payload_rd = decode_input_payload_rd;
  assign decode_load_payload_arg = decode_input_payload_arg;
  assign decode_load_payload_roundMode = decode_input_payload_roundMode;
  assign decode_load_payload_format = decode_input_payload_format;
  assign decode_load_payload_i2f = (decode_input_payload_opcode == FpuOpcode_I2F);
  assign decode_shortPipHit = (|{(decode_input_payload_opcode == FpuOpcode_FCVT_X_X),{(decode_input_payload_opcode == FpuOpcode_FCLASS),{(decode_input_payload_opcode == FpuOpcode_FMV_X_W),{(decode_input_payload_opcode == FpuOpcode_SGNJ),{(decode_input_payload_opcode == _zz_decode_shortPipHit),{_zz_decode_shortPipHit_1,{_zz_decode_shortPipHit_2,_zz_decode_shortPipHit_3}}}}}}});
  assign when_FpuCore_l335 = (decode_shortPipHit && decode_shortPip_ready);
  assign decode_shortPip_valid = (decode_input_valid && decode_shortPipHit);
  assign decode_shortPip_payload_source = decode_input_payload_source;
  assign decode_shortPip_payload_opcode = decode_input_payload_opcode;
  assign decode_shortPip_payload_rs1_mantissa = decode_input_payload_rs1_mantissa;
  assign decode_shortPip_payload_rs1_exponent = decode_input_payload_rs1_exponent;
  assign decode_shortPip_payload_rs1_sign = decode_input_payload_rs1_sign;
  assign decode_shortPip_payload_rs1_special = decode_input_payload_rs1_special;
  assign decode_shortPip_payload_rs2_mantissa = decode_input_payload_rs2_mantissa;
  assign decode_shortPip_payload_rs2_exponent = decode_input_payload_rs2_exponent;
  assign decode_shortPip_payload_rs2_sign = decode_input_payload_rs2_sign;
  assign decode_shortPip_payload_rs2_special = decode_input_payload_rs2_special;
  assign decode_shortPip_payload_rd = decode_input_payload_rd;
  assign decode_shortPip_payload_arg = decode_input_payload_arg;
  assign decode_shortPip_payload_roundMode = decode_input_payload_roundMode;
  assign decode_shortPip_payload_format = decode_input_payload_format;
  assign decode_shortPip_payload_rs1Boxed = decode_input_payload_rs1Boxed;
  assign decode_shortPip_payload_rs2Boxed = decode_input_payload_rs2Boxed;
  assign decode_divSqrtHit = ((decode_input_payload_opcode == FpuOpcode_DIV) || (decode_input_payload_opcode == FpuOpcode_SQRT));
  assign decode_divHit = (decode_input_payload_opcode == FpuOpcode_DIV);
  assign when_FpuCore_l351 = (decode_divHit && decode_div_ready);
  assign decode_div_valid = (decode_input_valid && decode_divHit);
  assign decode_div_payload_source = decode_input_payload_source;
  assign decode_div_payload_rs1_mantissa = decode_input_payload_rs1_mantissa;
  assign decode_div_payload_rs1_exponent = decode_input_payload_rs1_exponent;
  assign decode_div_payload_rs1_sign = decode_input_payload_rs1_sign;
  assign decode_div_payload_rs1_special = decode_input_payload_rs1_special;
  assign decode_div_payload_rs2_mantissa = decode_input_payload_rs2_mantissa;
  assign decode_div_payload_rs2_exponent = decode_input_payload_rs2_exponent;
  assign decode_div_payload_rs2_sign = decode_input_payload_rs2_sign;
  assign decode_div_payload_rs2_special = decode_input_payload_rs2_special;
  assign decode_div_payload_rd = decode_input_payload_rd;
  assign decode_div_payload_roundMode = decode_input_payload_roundMode;
  assign decode_div_payload_format = decode_input_payload_format;
  assign decode_sqrtHit = (decode_input_payload_opcode == FpuOpcode_SQRT);
  assign when_FpuCore_l359 = (decode_sqrtHit && decode_sqrt_ready);
  assign decode_sqrt_valid = (decode_input_valid && decode_sqrtHit);
  assign decode_sqrt_payload_source = decode_input_payload_source;
  assign decode_sqrt_payload_rs1_mantissa = decode_input_payload_rs1_mantissa;
  assign decode_sqrt_payload_rs1_exponent = decode_input_payload_rs1_exponent;
  assign decode_sqrt_payload_rs1_sign = decode_input_payload_rs1_sign;
  assign decode_sqrt_payload_rs1_special = decode_input_payload_rs1_special;
  assign decode_sqrt_payload_rd = decode_input_payload_rd;
  assign decode_sqrt_payload_roundMode = decode_input_payload_roundMode;
  assign decode_sqrt_payload_format = decode_input_payload_format;
  assign decode_fmaHit = (decode_input_payload_opcode == FpuOpcode_FMA);
  assign decode_mulHit = ((decode_input_payload_opcode == FpuOpcode_MUL) || decode_fmaHit);
  assign decode_divSqrtToMul_valid = 1'b0;
  assign decode_divSqrtToMul_payload_source = 1'bx;
  assign decode_divSqrtToMul_payload_rs1_mantissa = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign decode_divSqrtToMul_payload_rs1_exponent = 12'bxxxxxxxxxxxx;
  assign decode_divSqrtToMul_payload_rs1_sign = 1'bx;
  assign decode_divSqrtToMul_payload_rs1_special = 1'bx;
  assign decode_divSqrtToMul_payload_rs2_mantissa = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign decode_divSqrtToMul_payload_rs2_exponent = 12'bxxxxxxxxxxxx;
  assign decode_divSqrtToMul_payload_rs2_sign = 1'bx;
  assign decode_divSqrtToMul_payload_rs2_special = 1'bx;
  assign decode_divSqrtToMul_payload_rs3_mantissa = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign decode_divSqrtToMul_payload_rs3_exponent = 12'bxxxxxxxxxxxx;
  assign decode_divSqrtToMul_payload_rs3_sign = 1'bx;
  assign decode_divSqrtToMul_payload_rs3_special = 1'bx;
  assign decode_divSqrtToMul_payload_rd = 5'bxxxxx;
  assign decode_divSqrtToMul_payload_add = 1'bx;
  assign decode_divSqrtToMul_payload_divSqrt = 1'bx;
  assign decode_divSqrtToMul_payload_msb1 = 1'bx;
  assign decode_divSqrtToMul_payload_msb2 = 1'bx;
  assign decode_divSqrtToMul_payload_roundMode = (3'bxxx);
  assign decode_divSqrtToMul_payload_format = (1'bx);
  assign when_FpuCore_l375 = ((decode_mulHit && decode_mul_ready) && (! decode_divSqrtToMul_valid));
  assign decode_mul_valid = ((decode_input_valid && decode_mulHit) || decode_divSqrtToMul_valid);
  assign decode_divSqrtToMul_ready = decode_mul_ready;
  always @(*) begin
    decode_mul_payload_source = decode_divSqrtToMul_payload_source;
    if(when_FpuCore_l380) begin
      decode_mul_payload_source = decode_input_payload_source;
    end
  end

  always @(*) begin
    decode_mul_payload_rs1_mantissa = decode_divSqrtToMul_payload_rs1_mantissa;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs1_mantissa = decode_input_payload_rs1_mantissa;
    end
  end

  always @(*) begin
    decode_mul_payload_rs1_exponent = decode_divSqrtToMul_payload_rs1_exponent;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs1_exponent = decode_input_payload_rs1_exponent;
    end
  end

  always @(*) begin
    decode_mul_payload_rs1_sign = decode_divSqrtToMul_payload_rs1_sign;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs1_sign = decode_input_payload_rs1_sign;
    end
  end

  always @(*) begin
    decode_mul_payload_rs1_special = decode_divSqrtToMul_payload_rs1_special;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs1_special = decode_input_payload_rs1_special;
    end
  end

  always @(*) begin
    decode_mul_payload_rs2_mantissa = decode_divSqrtToMul_payload_rs2_mantissa;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs2_mantissa = decode_input_payload_rs2_mantissa;
    end
  end

  always @(*) begin
    decode_mul_payload_rs2_exponent = decode_divSqrtToMul_payload_rs2_exponent;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs2_exponent = decode_input_payload_rs2_exponent;
    end
  end

  always @(*) begin
    decode_mul_payload_rs2_sign = decode_divSqrtToMul_payload_rs2_sign;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs2_sign = decode_input_payload_rs2_sign;
      decode_mul_payload_rs2_sign = (decode_input_payload_rs2_sign ^ decode_input_payload_arg[0]);
    end
  end

  always @(*) begin
    decode_mul_payload_rs2_special = decode_divSqrtToMul_payload_rs2_special;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs2_special = decode_input_payload_rs2_special;
    end
  end

  always @(*) begin
    decode_mul_payload_rs3_mantissa = decode_divSqrtToMul_payload_rs3_mantissa;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs3_mantissa = decode_input_payload_rs3_mantissa;
    end
  end

  always @(*) begin
    decode_mul_payload_rs3_exponent = decode_divSqrtToMul_payload_rs3_exponent;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs3_exponent = decode_input_payload_rs3_exponent;
    end
  end

  always @(*) begin
    decode_mul_payload_rs3_sign = decode_divSqrtToMul_payload_rs3_sign;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs3_sign = decode_input_payload_rs3_sign;
      decode_mul_payload_rs3_sign = (decode_input_payload_rs3_sign ^ decode_input_payload_arg[1]);
    end
  end

  always @(*) begin
    decode_mul_payload_rs3_special = decode_divSqrtToMul_payload_rs3_special;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rs3_special = decode_input_payload_rs3_special;
    end
  end

  always @(*) begin
    decode_mul_payload_rd = decode_divSqrtToMul_payload_rd;
    if(when_FpuCore_l380) begin
      decode_mul_payload_rd = decode_input_payload_rd;
    end
  end

  always @(*) begin
    decode_mul_payload_add = decode_divSqrtToMul_payload_add;
    if(when_FpuCore_l380) begin
      decode_mul_payload_add = decode_fmaHit;
    end
  end

  always @(*) begin
    decode_mul_payload_divSqrt = decode_divSqrtToMul_payload_divSqrt;
    if(when_FpuCore_l380) begin
      decode_mul_payload_divSqrt = 1'b0;
    end
  end

  always @(*) begin
    decode_mul_payload_msb1 = decode_divSqrtToMul_payload_msb1;
    if(when_FpuCore_l380) begin
      decode_mul_payload_msb1 = 1'b1;
    end
  end

  always @(*) begin
    decode_mul_payload_msb2 = decode_divSqrtToMul_payload_msb2;
    if(when_FpuCore_l380) begin
      decode_mul_payload_msb2 = 1'b1;
    end
  end

  always @(*) begin
    decode_mul_payload_roundMode = decode_divSqrtToMul_payload_roundMode;
    if(when_FpuCore_l380) begin
      decode_mul_payload_roundMode = decode_input_payload_roundMode;
    end
  end

  always @(*) begin
    decode_mul_payload_format = decode_divSqrtToMul_payload_format;
    if(when_FpuCore_l380) begin
      decode_mul_payload_format = decode_input_payload_format;
    end
  end

  assign when_FpuCore_l380 = (! decode_divSqrtToMul_valid);
  assign decode_addHit = (decode_input_payload_opcode == FpuOpcode_ADD);
  assign when_FpuCore_l399 = ((decode_addHit && decode_add_ready) && (! decode_mulToAdd_valid));
  assign decode_add_valid = ((decode_input_valid && decode_addHit) || decode_mulToAdd_valid);
  assign decode_mulToAdd_ready = decode_add_ready;
  always @(*) begin
    decode_add_payload_source = decode_mulToAdd_payload_source;
    if(when_FpuCore_l404) begin
      decode_add_payload_source = decode_input_payload_source;
    end
  end

  always @(*) begin
    decode_add_payload_rs1_mantissa = decode_mulToAdd_payload_rs1_mantissa;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs1_mantissa = ({2'd0,decode_input_payload_rs1_mantissa} <<< 2'd2);
    end
  end

  always @(*) begin
    decode_add_payload_rs1_exponent = decode_mulToAdd_payload_rs1_exponent;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs1_exponent = decode_input_payload_rs1_exponent;
    end
  end

  always @(*) begin
    decode_add_payload_rs1_sign = decode_mulToAdd_payload_rs1_sign;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs1_sign = decode_input_payload_rs1_sign;
    end
  end

  always @(*) begin
    decode_add_payload_rs1_special = decode_mulToAdd_payload_rs1_special;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs1_special = decode_input_payload_rs1_special;
    end
  end

  always @(*) begin
    decode_add_payload_rs2_mantissa = decode_mulToAdd_payload_rs2_mantissa;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs2_mantissa = ({2'd0,decode_input_payload_rs2_mantissa} <<< 2'd2);
    end
  end

  always @(*) begin
    decode_add_payload_rs2_exponent = decode_mulToAdd_payload_rs2_exponent;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs2_exponent = decode_input_payload_rs2_exponent;
    end
  end

  always @(*) begin
    decode_add_payload_rs2_sign = decode_mulToAdd_payload_rs2_sign;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs2_sign = (decode_input_payload_rs2_sign ^ decode_input_payload_arg[0]);
    end
  end

  always @(*) begin
    decode_add_payload_rs2_special = decode_mulToAdd_payload_rs2_special;
    if(when_FpuCore_l404) begin
      decode_add_payload_rs2_special = decode_input_payload_rs2_special;
    end
  end

  always @(*) begin
    decode_add_payload_rd = decode_mulToAdd_payload_rd;
    if(when_FpuCore_l404) begin
      decode_add_payload_rd = decode_input_payload_rd;
    end
  end

  always @(*) begin
    decode_add_payload_roundMode = decode_mulToAdd_payload_roundMode;
    if(when_FpuCore_l404) begin
      decode_add_payload_roundMode = decode_input_payload_roundMode;
    end
  end

  always @(*) begin
    decode_add_payload_format = decode_mulToAdd_payload_format;
    if(when_FpuCore_l404) begin
      decode_add_payload_format = decode_input_payload_format;
    end
  end

  always @(*) begin
    decode_add_payload_needCommit = decode_mulToAdd_payload_needCommit;
    if(when_FpuCore_l404) begin
      decode_add_payload_needCommit = 1'b1;
    end
  end

  assign when_FpuCore_l404 = (! decode_mulToAdd_valid);
  assign decode_load_ready = decode_load_rValidN;
  assign decode_load_s2mPipe_valid = (decode_load_valid || (! decode_load_rValidN));
  assign _zz_decode_load_s2mPipe_payload_roundMode = (decode_load_rValidN ? decode_load_payload_roundMode : decode_load_rData_roundMode);
  assign _zz_decode_load_s2mPipe_payload_format = (decode_load_rValidN ? decode_load_payload_format : decode_load_rData_format);
  assign decode_load_s2mPipe_payload_source = (decode_load_rValidN ? decode_load_payload_source : decode_load_rData_source);
  assign decode_load_s2mPipe_payload_rd = (decode_load_rValidN ? decode_load_payload_rd : decode_load_rData_rd);
  assign decode_load_s2mPipe_payload_i2f = (decode_load_rValidN ? decode_load_payload_i2f : decode_load_rData_i2f);
  assign decode_load_s2mPipe_payload_arg = (decode_load_rValidN ? decode_load_payload_arg : decode_load_rData_arg);
  assign decode_load_s2mPipe_payload_roundMode = _zz_decode_load_s2mPipe_payload_roundMode;
  assign decode_load_s2mPipe_payload_format = _zz_decode_load_s2mPipe_payload_format;
  always @(*) begin
    decode_load_s2mPipe_ready = decode_load_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375_3) begin
      decode_load_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_3 = (! decode_load_s2mPipe_m2sPipe_valid);
  assign decode_load_s2mPipe_m2sPipe_valid = decode_load_s2mPipe_rValid;
  assign decode_load_s2mPipe_m2sPipe_payload_source = decode_load_s2mPipe_rData_source;
  assign decode_load_s2mPipe_m2sPipe_payload_rd = decode_load_s2mPipe_rData_rd;
  assign decode_load_s2mPipe_m2sPipe_payload_i2f = decode_load_s2mPipe_rData_i2f;
  assign decode_load_s2mPipe_m2sPipe_payload_arg = decode_load_s2mPipe_rData_arg;
  assign decode_load_s2mPipe_m2sPipe_payload_roundMode = decode_load_s2mPipe_rData_roundMode;
  assign decode_load_s2mPipe_m2sPipe_payload_format = decode_load_s2mPipe_rData_format;
  always @(*) begin
    decode_load_s2mPipe_m2sPipe_ready = load_s0_input_ready;
    if(when_Stream_l375_4) begin
      decode_load_s2mPipe_m2sPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375_4 = (! load_s0_input_valid);
  assign load_s0_input_valid = decode_load_s2mPipe_m2sPipe_rValid;
  assign load_s0_input_payload_source = decode_load_s2mPipe_m2sPipe_rData_source;
  assign load_s0_input_payload_rd = decode_load_s2mPipe_m2sPipe_rData_rd;
  assign load_s0_input_payload_i2f = decode_load_s2mPipe_m2sPipe_rData_i2f;
  assign load_s0_input_payload_arg = decode_load_s2mPipe_m2sPipe_rData_arg;
  assign load_s0_input_payload_roundMode = decode_load_s2mPipe_m2sPipe_rData_roundMode;
  assign load_s0_input_payload_format = decode_load_s2mPipe_m2sPipe_rData_format;
  assign when_Stream_l445 = (! (|{(commitFork_load_0_payload_opcode == FpuOpcode_I2F),{(commitFork_load_0_payload_opcode == FpuOpcode_FMV_W_X),(commitFork_load_0_payload_opcode == FpuOpcode_LOAD)}}));
  always @(*) begin
    load_s0_filtred_0_valid = commitFork_load_0_valid;
    if(when_Stream_l445) begin
      load_s0_filtred_0_valid = 1'b0;
    end
  end

  always @(*) begin
    commitFork_load_0_ready = load_s0_filtred_0_ready;
    if(when_Stream_l445) begin
      commitFork_load_0_ready = 1'b1;
    end
  end

  assign load_s0_filtred_0_payload_opcode = commitFork_load_0_payload_opcode;
  assign load_s0_filtred_0_payload_rd = commitFork_load_0_payload_rd;
  assign load_s0_filtred_0_payload_write = commitFork_load_0_payload_write;
  assign load_s0_filtred_0_payload_value = commitFork_load_0_payload_value;
  assign when_Stream_l445_1 = (! (|{(commitFork_load_1_payload_opcode == FpuOpcode_I2F),{(commitFork_load_1_payload_opcode == FpuOpcode_FMV_W_X),(commitFork_load_1_payload_opcode == FpuOpcode_LOAD)}}));
  always @(*) begin
    load_s0_filtred_1_valid = commitFork_load_1_valid;
    if(when_Stream_l445_1) begin
      load_s0_filtred_1_valid = 1'b0;
    end
  end

  always @(*) begin
    commitFork_load_1_ready = load_s0_filtred_1_ready;
    if(when_Stream_l445_1) begin
      commitFork_load_1_ready = 1'b1;
    end
  end

  assign load_s0_filtred_1_payload_opcode = commitFork_load_1_payload_opcode;
  assign load_s0_filtred_1_payload_rd = commitFork_load_1_payload_rd;
  assign load_s0_filtred_1_payload_write = commitFork_load_1_payload_write;
  assign load_s0_filtred_1_payload_value = commitFork_load_1_payload_value;
  assign load_s0_hazard = (! _zz_load_s0_hazard);
  assign _zz_load_s0_input_ready = (! load_s0_hazard);
  assign load_s0_input_ready = (load_s0_output_ready && _zz_load_s0_input_ready);
  assign load_s0_output_valid = (load_s0_input_valid && _zz_load_s0_input_ready);
  always @(*) begin
    load_s0_filtred_0_ready = 1'b0;
    if(_zz_33[0]) begin
      load_s0_filtred_0_ready = _zz_load_s0_filtred_0_ready;
    end
  end

  always @(*) begin
    load_s0_filtred_1_ready = 1'b0;
    if(_zz_33[1]) begin
      load_s0_filtred_1_ready = _zz_load_s0_filtred_0_ready;
    end
  end

  assign _zz_33 = ({1'd0,1'b1} <<< load_s0_input_payload_source);
  assign _zz_load_s0_filtred_0_ready = (load_s0_input_valid && load_s0_output_ready);
  assign load_s0_output_payload_source = load_s0_input_payload_source;
  assign load_s0_output_payload_rd = load_s0_input_payload_rd;
  assign load_s0_output_payload_value = _zz_load_s0_output_payload_value;
  assign load_s0_output_payload_i2f = load_s0_input_payload_i2f;
  assign load_s0_output_payload_arg = load_s0_input_payload_arg;
  assign load_s0_output_payload_roundMode = load_s0_input_payload_roundMode;
  always @(*) begin
    load_s0_output_payload_format = load_s0_input_payload_format;
    if(when_FpuCore_l452) begin
      load_s0_output_payload_format = FpuFormat_FLOAT;
    end
  end

  assign when_FpuCore_l452 = (((! load_s0_input_payload_i2f) && (load_s0_input_payload_format == FpuFormat_DOUBLE)) && (&load_s0_output_payload_value[63 : 32]));
  always @(*) begin
    load_s0_output_ready = load_s1_input_ready;
    if(when_Stream_l375_5) begin
      load_s0_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_5 = (! load_s1_input_valid);
  assign load_s1_input_valid = load_s0_output_rValid;
  assign load_s1_input_payload_source = load_s0_output_rData_source;
  assign load_s1_input_payload_rd = load_s0_output_rData_rd;
  assign load_s1_input_payload_value = load_s0_output_rData_value;
  assign load_s1_input_payload_i2f = load_s0_output_rData_i2f;
  assign load_s1_input_payload_arg = load_s0_output_rData_arg;
  assign load_s1_input_payload_roundMode = load_s0_output_rData_roundMode;
  assign load_s1_input_payload_format = load_s0_output_rData_format;
  always @(*) begin
    load_s1_busy = 1'b0;
    if(when_FpuCore_l529) begin
      load_s1_busy = 1'b1;
    end
  end

  assign load_s1_f32_mantissa = load_s1_input_payload_value[22 : 0];
  assign load_s1_f32_exponent = load_s1_input_payload_value[30 : 23];
  assign load_s1_f32_sign = load_s1_input_payload_value[31];
  assign load_s1_f64_mantissa = load_s1_input_payload_value[51 : 0];
  assign load_s1_f64_exponent = load_s1_input_payload_value[62 : 52];
  assign load_s1_f64_sign = load_s1_input_payload_value[63];
  assign load_s1_passThroughFloat_special = 1'b0;
  assign when_FpuCore_l31 = (load_s1_input_payload_format == FpuFormat_DOUBLE);
  always @(*) begin
    if(when_FpuCore_l31) begin
      load_s1_passThroughFloat_sign = load_s1_f64_sign;
    end else begin
      load_s1_passThroughFloat_sign = load_s1_f32_sign;
    end
  end

  always @(*) begin
    if(when_FpuCore_l31) begin
      load_s1_passThroughFloat_exponent = {1'd0, load_s1_f64_exponent};
    end else begin
      load_s1_passThroughFloat_exponent = {4'd0, load_s1_f32_exponent};
    end
  end

  always @(*) begin
    if(when_FpuCore_l31) begin
      load_s1_passThroughFloat_mantissa = load_s1_f64_mantissa;
    end else begin
      load_s1_passThroughFloat_mantissa = ({29'd0,load_s1_f32_mantissa} <<< 5'd29);
    end
  end

  always @(*) begin
    if(when_FpuCore_l31) begin
      load_s1_recodedExpOffset = 12'h400;
    end else begin
      load_s1_recodedExpOffset = 12'h780;
    end
  end

  assign load_s1_manZero = (load_s1_passThroughFloat_mantissa == 52'h0);
  always @(*) begin
    load_s1_expZero = (load_s1_passThroughFloat_exponent == 12'h0);
    if(when_FpuCore_l494) begin
      load_s1_expZero = 1'b0;
    end
  end

  always @(*) begin
    load_s1_expOne = (&load_s1_passThroughFloat_exponent[7 : 0]);
    if(when_FpuCore_l495) begin
      load_s1_expOne = 1'b0;
    end
  end

  assign when_FpuCore_l494 = ((load_s1_input_payload_format == FpuFormat_DOUBLE) && (load_s1_input_payload_value[62 : 60] != 3'b000));
  assign when_FpuCore_l495 = ((load_s1_input_payload_format == FpuFormat_DOUBLE) && (load_s1_input_payload_value[62 : 60] != 3'b111));
  assign load_s1_isZero = (load_s1_expZero && load_s1_manZero);
  assign load_s1_isSubnormal = (load_s1_expZero && (! load_s1_manZero));
  assign load_s1_isInfinity = (load_s1_expOne && load_s1_manZero);
  assign load_s1_isNan = (load_s1_expOne && (! load_s1_manZero));
  always @(*) begin
    load_s1_fsm_ohInput = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_FpuCore_l508) begin
      load_s1_fsm_ohInput = load_s1_passThroughFloat_mantissa;
    end else begin
      load_s1_fsm_ohInput[19 : 0] = 20'h0;
      load_s1_fsm_ohInput[51 : 20] = load_s1_input_payload_value[31 : 0];
    end
  end

  assign when_FpuCore_l508 = (! load_s1_input_payload_i2f);
  always @(*) begin
    load_s1_fsm_shift_input = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    load_s1_fsm_shift_input = (load_s1_fsm_ohInput <<< 1);
  end

  assign when_FpuCore_l525 = (! load_s1_fsm_done);
  assign when_FpuCore_l529 = ((load_s1_input_valid && (load_s1_input_payload_i2f || load_s1_isSubnormal)) && (! load_s1_fsm_done));
  assign when_FpuCore_l532 = (((load_s1_input_payload_i2f && (! load_s1_fsm_patched)) && load_s1_input_payload_value[31]) && load_s1_input_payload_arg[0]);
  assign _zz_load_s0_output_rData_value = load_s1_input_payload_value;
  assign _zz_load_s0_output_rData_value_1 = 1'b1;
  assign _zz_load_s1_fsm_shift_by = {load_s1_fsm_ohInput[0],{load_s1_fsm_ohInput[1],{load_s1_fsm_ohInput[2],{load_s1_fsm_ohInput[3],{load_s1_fsm_ohInput[4],{load_s1_fsm_ohInput[5],{load_s1_fsm_ohInput[6],{_zz__zz_load_s1_fsm_shift_by,{_zz__zz_load_s1_fsm_shift_by_1,_zz__zz_load_s1_fsm_shift_by_2}}}}}}}}};
  assign _zz_load_s1_fsm_shift_by_1 = (_zz_load_s1_fsm_shift_by & (~ _zz__zz_load_s1_fsm_shift_by_1_1));
  assign _zz_load_s1_fsm_shift_by_2 = _zz_load_s1_fsm_shift_by_1[3];
  assign _zz_load_s1_fsm_shift_by_3 = _zz_load_s1_fsm_shift_by_1[5];
  assign _zz_load_s1_fsm_shift_by_4 = _zz_load_s1_fsm_shift_by_1[6];
  assign _zz_load_s1_fsm_shift_by_5 = _zz_load_s1_fsm_shift_by_1[7];
  assign _zz_load_s1_fsm_shift_by_6 = _zz_load_s1_fsm_shift_by_1[9];
  assign _zz_load_s1_fsm_shift_by_7 = _zz_load_s1_fsm_shift_by_1[10];
  assign _zz_load_s1_fsm_shift_by_8 = _zz_load_s1_fsm_shift_by_1[11];
  assign _zz_load_s1_fsm_shift_by_9 = _zz_load_s1_fsm_shift_by_1[12];
  assign _zz_load_s1_fsm_shift_by_10 = _zz_load_s1_fsm_shift_by_1[13];
  assign _zz_load_s1_fsm_shift_by_11 = _zz_load_s1_fsm_shift_by_1[14];
  assign _zz_load_s1_fsm_shift_by_12 = _zz_load_s1_fsm_shift_by_1[15];
  assign _zz_load_s1_fsm_shift_by_13 = _zz_load_s1_fsm_shift_by_1[17];
  assign _zz_load_s1_fsm_shift_by_14 = _zz_load_s1_fsm_shift_by_1[18];
  assign _zz_load_s1_fsm_shift_by_15 = _zz_load_s1_fsm_shift_by_1[19];
  assign _zz_load_s1_fsm_shift_by_16 = _zz_load_s1_fsm_shift_by_1[20];
  assign _zz_load_s1_fsm_shift_by_17 = _zz_load_s1_fsm_shift_by_1[21];
  assign _zz_load_s1_fsm_shift_by_18 = _zz_load_s1_fsm_shift_by_1[22];
  assign _zz_load_s1_fsm_shift_by_19 = _zz_load_s1_fsm_shift_by_1[23];
  assign _zz_load_s1_fsm_shift_by_20 = _zz_load_s1_fsm_shift_by_1[24];
  assign _zz_load_s1_fsm_shift_by_21 = _zz_load_s1_fsm_shift_by_1[25];
  assign _zz_load_s1_fsm_shift_by_22 = _zz_load_s1_fsm_shift_by_1[26];
  assign _zz_load_s1_fsm_shift_by_23 = _zz_load_s1_fsm_shift_by_1[27];
  assign _zz_load_s1_fsm_shift_by_24 = _zz_load_s1_fsm_shift_by_1[28];
  assign _zz_load_s1_fsm_shift_by_25 = _zz_load_s1_fsm_shift_by_1[29];
  assign _zz_load_s1_fsm_shift_by_26 = _zz_load_s1_fsm_shift_by_1[30];
  assign _zz_load_s1_fsm_shift_by_27 = _zz_load_s1_fsm_shift_by_1[31];
  assign _zz_load_s1_fsm_shift_by_28 = _zz_load_s1_fsm_shift_by_1[33];
  assign _zz_load_s1_fsm_shift_by_29 = _zz_load_s1_fsm_shift_by_1[34];
  assign _zz_load_s1_fsm_shift_by_30 = _zz_load_s1_fsm_shift_by_1[35];
  assign _zz_load_s1_fsm_shift_by_31 = _zz_load_s1_fsm_shift_by_1[36];
  assign _zz_load_s1_fsm_shift_by_32 = _zz_load_s1_fsm_shift_by_1[37];
  assign _zz_load_s1_fsm_shift_by_33 = _zz_load_s1_fsm_shift_by_1[38];
  assign _zz_load_s1_fsm_shift_by_34 = _zz_load_s1_fsm_shift_by_1[39];
  assign _zz_load_s1_fsm_shift_by_35 = _zz_load_s1_fsm_shift_by_1[40];
  assign _zz_load_s1_fsm_shift_by_36 = _zz_load_s1_fsm_shift_by_1[41];
  assign _zz_load_s1_fsm_shift_by_37 = _zz_load_s1_fsm_shift_by_1[42];
  assign _zz_load_s1_fsm_shift_by_38 = _zz_load_s1_fsm_shift_by_1[43];
  assign _zz_load_s1_fsm_shift_by_39 = _zz_load_s1_fsm_shift_by_1[44];
  assign _zz_load_s1_fsm_shift_by_40 = _zz_load_s1_fsm_shift_by_1[45];
  assign _zz_load_s1_fsm_shift_by_41 = _zz_load_s1_fsm_shift_by_1[46];
  assign _zz_load_s1_fsm_shift_by_42 = _zz_load_s1_fsm_shift_by_1[47];
  assign _zz_load_s1_fsm_shift_by_43 = _zz_load_s1_fsm_shift_by_1[48];
  assign _zz_load_s1_fsm_shift_by_44 = _zz_load_s1_fsm_shift_by_1[49];
  assign _zz_load_s1_fsm_shift_by_45 = _zz_load_s1_fsm_shift_by_1[50];
  assign _zz_load_s1_fsm_shift_by_46 = _zz_load_s1_fsm_shift_by_1[51];
  assign _zz_load_s1_fsm_shift_by_47 = ((((((((((((((((_zz__zz_load_s1_fsm_shift_by_47 || _zz_load_s1_fsm_shift_by_17) || _zz_load_s1_fsm_shift_by_19) || _zz_load_s1_fsm_shift_by_21) || _zz_load_s1_fsm_shift_by_23) || _zz_load_s1_fsm_shift_by_25) || _zz_load_s1_fsm_shift_by_27) || _zz_load_s1_fsm_shift_by_28) || _zz_load_s1_fsm_shift_by_30) || _zz_load_s1_fsm_shift_by_32) || _zz_load_s1_fsm_shift_by_34) || _zz_load_s1_fsm_shift_by_36) || _zz_load_s1_fsm_shift_by_38) || _zz_load_s1_fsm_shift_by_40) || _zz_load_s1_fsm_shift_by_42) || _zz_load_s1_fsm_shift_by_44) || _zz_load_s1_fsm_shift_by_46);
  assign _zz_load_s1_fsm_shift_by_48 = ((((((((((((((((_zz__zz_load_s1_fsm_shift_by_48 || _zz_load_s1_fsm_shift_by_18) || _zz_load_s1_fsm_shift_by_19) || _zz_load_s1_fsm_shift_by_22) || _zz_load_s1_fsm_shift_by_23) || _zz_load_s1_fsm_shift_by_26) || _zz_load_s1_fsm_shift_by_27) || _zz_load_s1_fsm_shift_by_29) || _zz_load_s1_fsm_shift_by_30) || _zz_load_s1_fsm_shift_by_33) || _zz_load_s1_fsm_shift_by_34) || _zz_load_s1_fsm_shift_by_37) || _zz_load_s1_fsm_shift_by_38) || _zz_load_s1_fsm_shift_by_41) || _zz_load_s1_fsm_shift_by_42) || _zz_load_s1_fsm_shift_by_45) || _zz_load_s1_fsm_shift_by_46);
  assign _zz_load_s1_fsm_shift_by_49 = (((((((((((((((((_zz__zz_load_s1_fsm_shift_by_49 || _zz_load_s1_fsm_shift_by_12) || _zz_load_s1_fsm_shift_by_16) || _zz_load_s1_fsm_shift_by_17) || _zz_load_s1_fsm_shift_by_18) || _zz_load_s1_fsm_shift_by_19) || _zz_load_s1_fsm_shift_by_24) || _zz_load_s1_fsm_shift_by_25) || _zz_load_s1_fsm_shift_by_26) || _zz_load_s1_fsm_shift_by_27) || _zz_load_s1_fsm_shift_by_31) || _zz_load_s1_fsm_shift_by_32) || _zz_load_s1_fsm_shift_by_33) || _zz_load_s1_fsm_shift_by_34) || _zz_load_s1_fsm_shift_by_39) || _zz_load_s1_fsm_shift_by_40) || _zz_load_s1_fsm_shift_by_41) || _zz_load_s1_fsm_shift_by_42);
  assign _zz_load_s1_fsm_shift_by_50 = ((((((((((((((((_zz__zz_load_s1_fsm_shift_by_50 || _zz_load_s1_fsm_shift_by_20) || _zz_load_s1_fsm_shift_by_21) || _zz_load_s1_fsm_shift_by_22) || _zz_load_s1_fsm_shift_by_23) || _zz_load_s1_fsm_shift_by_24) || _zz_load_s1_fsm_shift_by_25) || _zz_load_s1_fsm_shift_by_26) || _zz_load_s1_fsm_shift_by_27) || _zz_load_s1_fsm_shift_by_35) || _zz_load_s1_fsm_shift_by_36) || _zz_load_s1_fsm_shift_by_37) || _zz_load_s1_fsm_shift_by_38) || _zz_load_s1_fsm_shift_by_39) || _zz_load_s1_fsm_shift_by_40) || _zz_load_s1_fsm_shift_by_41) || _zz_load_s1_fsm_shift_by_42);
  assign _zz_load_s1_fsm_shift_by_51 = (((((((((((((((((_zz__zz_load_s1_fsm_shift_by_51 || _zz_load_s1_fsm_shift_by_15) || _zz_load_s1_fsm_shift_by_16) || _zz_load_s1_fsm_shift_by_17) || _zz_load_s1_fsm_shift_by_18) || _zz_load_s1_fsm_shift_by_19) || _zz_load_s1_fsm_shift_by_20) || _zz_load_s1_fsm_shift_by_21) || _zz_load_s1_fsm_shift_by_22) || _zz_load_s1_fsm_shift_by_23) || _zz_load_s1_fsm_shift_by_24) || _zz_load_s1_fsm_shift_by_25) || _zz_load_s1_fsm_shift_by_26) || _zz_load_s1_fsm_shift_by_27) || _zz_load_s1_fsm_shift_by_43) || _zz_load_s1_fsm_shift_by_44) || _zz_load_s1_fsm_shift_by_45) || _zz_load_s1_fsm_shift_by_46);
  assign _zz_load_s1_fsm_shift_by_52 = ((((((((((((((((_zz__zz_load_s1_fsm_shift_by_52 || _zz_load_s1_fsm_shift_by_31) || _zz_load_s1_fsm_shift_by_32) || _zz_load_s1_fsm_shift_by_33) || _zz_load_s1_fsm_shift_by_34) || _zz_load_s1_fsm_shift_by_35) || _zz_load_s1_fsm_shift_by_36) || _zz_load_s1_fsm_shift_by_37) || _zz_load_s1_fsm_shift_by_38) || _zz_load_s1_fsm_shift_by_39) || _zz_load_s1_fsm_shift_by_40) || _zz_load_s1_fsm_shift_by_41) || _zz_load_s1_fsm_shift_by_42) || _zz_load_s1_fsm_shift_by_43) || _zz_load_s1_fsm_shift_by_44) || _zz_load_s1_fsm_shift_by_45) || _zz_load_s1_fsm_shift_by_46);
  always @(*) begin
    load_s1_fsm_expOffset = 12'h0;
    if(load_s1_isSubnormal) begin
      load_s1_fsm_expOffset = {6'd0, load_s1_fsm_shift_by};
    end
  end

  assign load_s1_input_isStall = (load_s1_input_valid && (! load_s1_input_ready));
  assign when_FpuCore_l551 = (! load_s1_input_isStall);
  assign load_s1_i2fHigh = load_s1_fsm_shift_output;
  assign load_s1_scrap = 1'b0;
  assign load_s1_recoded_mantissa = load_s1_passThroughFloat_mantissa;
  always @(*) begin
    load_s1_recoded_exponent = _zz_load_s1_recoded_exponent[11:0];
    if(load_s1_isZero) begin
      load_s1_recoded_exponent[1 : 0] = 2'b00;
    end
    if(load_s1_isInfinity) begin
      load_s1_recoded_exponent[1 : 0] = 2'b01;
    end
    if(load_s1_isNan) begin
      load_s1_recoded_exponent[1 : 0] = 2'b10;
      load_s1_recoded_exponent[2] = 1'b0;
    end
  end

  assign load_s1_recoded_sign = load_s1_passThroughFloat_sign;
  always @(*) begin
    load_s1_recoded_special = 1'b0;
    if(load_s1_isZero) begin
      load_s1_recoded_special = 1'b1;
    end
    if(load_s1_isInfinity) begin
      load_s1_recoded_special = 1'b1;
    end
    if(load_s1_isNan) begin
      load_s1_recoded_special = 1'b1;
    end
  end

  assign _zz_load_s1_input_ready = (! load_s1_busy);
  assign load_s1_input_ready = (load_s1_output_ready && _zz_load_s1_input_ready);
  assign load_s1_output_valid = (load_s1_input_valid && _zz_load_s1_input_ready);
  assign load_s1_output_payload_source = load_s1_input_payload_source;
  assign load_s1_output_payload_roundMode = load_s1_input_payload_roundMode;
  assign load_s1_output_payload_format = load_s1_input_payload_format;
  assign load_s1_output_payload_rd = load_s1_input_payload_rd;
  always @(*) begin
    load_s1_output_payload_value_sign = load_s1_recoded_sign;
    if(load_s1_input_payload_i2f) begin
      load_s1_output_payload_value_sign = load_s1_fsm_patched;
    end
  end

  always @(*) begin
    load_s1_output_payload_value_exponent = load_s1_recoded_exponent;
    if(load_s1_input_payload_i2f) begin
      load_s1_output_payload_value_exponent = (12'h81e - _zz_load_s1_output_payload_value_exponent);
      if(load_s1_fsm_i2fZero) begin
        load_s1_output_payload_value_exponent[1 : 0] = 2'b00;
      end
    end
  end

  always @(*) begin
    load_s1_output_payload_value_mantissa = {load_s1_recoded_mantissa,1'b0};
    if(when_FpuCore_l594) begin
      load_s1_output_payload_value_mantissa = {load_s1_i2fHigh,1'b0};
    end
  end

  always @(*) begin
    load_s1_output_payload_value_special = load_s1_recoded_special;
    if(load_s1_input_payload_i2f) begin
      load_s1_output_payload_value_special = 1'b0;
      if(load_s1_fsm_i2fZero) begin
        load_s1_output_payload_value_special = 1'b1;
      end
    end
  end

  always @(*) begin
    load_s1_output_payload_scrap = 1'b0;
    if(load_s1_input_payload_i2f) begin
      load_s1_output_payload_scrap = load_s1_scrap;
    end
  end

  assign load_s1_output_payload_NV = 1'b0;
  assign load_s1_output_payload_DZ = 1'b0;
  assign when_FpuCore_l594 = (load_s1_input_payload_i2f || load_s1_isSubnormal);
  always @(*) begin
    decode_shortPip_ready = shortPip_input_ready;
    if(when_Stream_l375_6) begin
      decode_shortPip_ready = 1'b1;
    end
  end

  assign when_Stream_l375_6 = (! shortPip_input_valid);
  assign shortPip_input_valid = decode_shortPip_rValid;
  assign shortPip_input_payload_source = decode_shortPip_rData_source;
  assign shortPip_input_payload_opcode = decode_shortPip_rData_opcode;
  assign shortPip_input_payload_rs1_mantissa = decode_shortPip_rData_rs1_mantissa;
  assign shortPip_input_payload_rs1_exponent = decode_shortPip_rData_rs1_exponent;
  assign shortPip_input_payload_rs1_sign = decode_shortPip_rData_rs1_sign;
  assign shortPip_input_payload_rs1_special = decode_shortPip_rData_rs1_special;
  assign shortPip_input_payload_rs2_mantissa = decode_shortPip_rData_rs2_mantissa;
  assign shortPip_input_payload_rs2_exponent = decode_shortPip_rData_rs2_exponent;
  assign shortPip_input_payload_rs2_sign = decode_shortPip_rData_rs2_sign;
  assign shortPip_input_payload_rs2_special = decode_shortPip_rData_rs2_special;
  assign shortPip_input_payload_rd = decode_shortPip_rData_rd;
  assign shortPip_input_payload_value = decode_shortPip_rData_value;
  assign shortPip_input_payload_arg = decode_shortPip_rData_arg;
  assign shortPip_input_payload_roundMode = decode_shortPip_rData_roundMode;
  assign shortPip_input_payload_format = decode_shortPip_rData_format;
  assign shortPip_input_payload_rs1Boxed = decode_shortPip_rData_rs1Boxed;
  assign shortPip_input_payload_rs2Boxed = decode_shortPip_rData_rs2Boxed;
  assign shortPip_toFpuRf = (|{(shortPip_input_payload_opcode == FpuOpcode_FCVT_X_X),{(shortPip_input_payload_opcode == FpuOpcode_SGNJ),(shortPip_input_payload_opcode == FpuOpcode_MIN_MAX)}});
  assign shortPip_input_fire = (shortPip_input_valid && shortPip_input_ready);
  assign _zz_when_FpuCore_l221 = (shortPip_input_fire && shortPip_toFpuRf);
  assign when_FpuCore_l221 = (_zz_when_FpuCore_l221 && (shortPip_input_payload_source == 1'b0));
  assign when_FpuCore_l221_1 = (_zz_when_FpuCore_l221 && (shortPip_input_payload_source == 1'b1));
  assign shortPip_isCommited = _zz_shortPip_isCommited;
  assign _zz_shortPip_rfOutput_ready = (! (! shortPip_isCommited));
  assign shortPip_output_valid = (shortPip_rfOutput_valid && _zz_shortPip_rfOutput_ready);
  assign shortPip_rfOutput_ready = (shortPip_output_ready && _zz_shortPip_rfOutput_ready);
  assign shortPip_output_payload_source = shortPip_rfOutput_payload_source;
  assign shortPip_output_payload_rd = shortPip_rfOutput_payload_rd;
  assign shortPip_output_payload_value_mantissa = shortPip_rfOutput_payload_value_mantissa;
  assign shortPip_output_payload_value_exponent = shortPip_rfOutput_payload_value_exponent;
  assign shortPip_output_payload_value_sign = shortPip_rfOutput_payload_value_sign;
  assign shortPip_output_payload_value_special = shortPip_rfOutput_payload_value_special;
  assign shortPip_output_payload_scrap = shortPip_rfOutput_payload_scrap;
  assign shortPip_output_payload_roundMode = shortPip_rfOutput_payload_roundMode;
  assign shortPip_output_payload_format = shortPip_rfOutput_payload_format;
  assign shortPip_output_payload_NV = shortPip_rfOutput_payload_NV;
  assign shortPip_output_payload_DZ = shortPip_rfOutput_payload_DZ;
  always @(*) begin
    shortPip_result = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(shortPip_input_payload_opcode)
      FpuOpcode_STORE : begin
        shortPip_result = shortPip_recodedResult;
      end
      FpuOpcode_FMV_X_W : begin
        shortPip_result = shortPip_recodedResult;
      end
      FpuOpcode_F2I : begin
        shortPip_result[31 : 0] = shortPip_f2i_result;
      end
      FpuOpcode_CMP : begin
        shortPip_result[31 : 0] = {31'd0, shortPip_cmpResult};
      end
      FpuOpcode_FCLASS : begin
        shortPip_result[31 : 0] = shortPip_fclassResult;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    shortPip_halt = 1'b0;
    if(when_FpuCore_l658) begin
      shortPip_halt = 1'b1;
    end
  end

  assign shortPip_f32_exp = _zz_shortPip_f32_exp[7:0];
  assign shortPip_f32_man = shortPip_input_payload_rs1_mantissa[51 : 29];
  assign shortPip_f64_exp = _zz_shortPip_f64_exp[10:0];
  assign shortPip_f64_man = shortPip_input_payload_rs1_mantissa;
  assign when_FpuCore_l31_1 = (shortPip_input_payload_format == FpuFormat_DOUBLE);
  always @(*) begin
    if(when_FpuCore_l31_1) begin
      shortPip_recodedResult = {{shortPip_input_payload_rs1_sign,shortPip_f64_exp},shortPip_f64_man};
    end else begin
      shortPip_recodedResult = {{{32'hffffffff,shortPip_input_payload_rs1_sign},shortPip_f32_exp},shortPip_f32_man};
    end
    if(shortPip_isSubnormal) begin
      shortPip_recodedResult[22 : 0] = shortPip_fsm_shift_output[22 : 0];
      if(when_FpuCore_l31_2) begin
        shortPip_recodedResult[51 : 23] = shortPip_fsm_shift_output[51 : 23];
      end
    end
    if(shortPip_mantissaForced) begin
      shortPip_recodedResult[22 : 0] = (shortPip_mantissaForcedValue ? 23'h7fffff : 23'h0);
      if(when_FpuCore_l31_3) begin
        shortPip_recodedResult[51 : 23] = (shortPip_mantissaForcedValue ? 29'h1fffffff : 29'h0);
      end
    end
    if(shortPip_exponentForced) begin
      if(when_FpuCore_l31_4) begin
        shortPip_recodedResult[62 : 52] = (shortPip_exponentForcedValue ? 11'h7ff : 11'h0);
      end else begin
        shortPip_recodedResult[30 : 23] = (shortPip_exponentForcedValue ? 8'hff : 8'h0);
      end
    end
    if(shortPip_cononicalForced) begin
      if(when_FpuCore_l31_5) begin
        shortPip_recodedResult[63] = 1'b0;
        shortPip_recodedResult[51] = 1'b1;
      end else begin
        shortPip_recodedResult[31] = 1'b0;
        shortPip_recodedResult[22] = 1'b1;
      end
    end
  end

  assign shortPip_expSubnormalThreshold = ((shortPip_input_payload_format == FpuFormat_DOUBLE) ? 11'h400 : 11'h780);
  assign shortPip_expInSubnormalRange = (shortPip_input_payload_rs1_exponent <= _zz_shortPip_expInSubnormalRange);
  assign shortPip_isSubnormal = ((! shortPip_input_payload_rs1_special) && shortPip_expInSubnormalRange);
  assign shortPip_isNormal = ((! shortPip_input_payload_rs1_special) && (! shortPip_expInSubnormalRange));
  assign shortPip_fsm_f2iShift = (shortPip_input_payload_rs1_exponent - 12'h7ff);
  assign shortPip_fsm_isF2i = (shortPip_input_payload_opcode == FpuOpcode_F2I);
  assign shortPip_fsm_needRecoding = ((|{(shortPip_input_payload_opcode == FpuOpcode_STORE),(shortPip_input_payload_opcode == FpuOpcode_FMV_X_W)}) && shortPip_isSubnormal);
  assign shortPip_fsm_isZero = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b00));
  always @(*) begin
    shortPip_fsm_shift_input = 53'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    shortPip_fsm_shift_input = {(! shortPip_fsm_isZero),shortPip_input_payload_rs1_mantissa};
  end

  assign when_FpuCore_l646 = (shortPip_fsm_shift_by[5] && (shortPip_fsm_shift_input[31 : 0] != 32'h0));
  assign when_FpuCore_l646_1 = (shortPip_fsm_shift_by[4] && (shortPip_fsm_shift_input_1[15 : 0] != 16'h0));
  assign when_FpuCore_l646_2 = (shortPip_fsm_shift_by[3] && (shortPip_fsm_shift_input_2[7 : 0] != 8'h0));
  assign when_FpuCore_l646_3 = (shortPip_fsm_shift_by[2] && (shortPip_fsm_shift_input_3[3 : 0] != 4'b0000));
  assign when_FpuCore_l646_4 = (shortPip_fsm_shift_by[1] && (shortPip_fsm_shift_input_4[1 : 0] != 2'b00));
  assign when_FpuCore_l646_5 = (shortPip_fsm_shift_by[0] && (shortPip_fsm_shift_input_5[0 : 0] != 1'b0));
  assign when_FpuCore_l652 = (! shortPip_fsm_done);
  assign shortPip_fsm_formatShiftOffset = ((shortPip_input_payload_format == FpuFormat_DOUBLE) ? 11'h401 : 11'h75e);
  assign when_FpuCore_l658 = ((shortPip_input_valid && (shortPip_fsm_needRecoding || shortPip_fsm_isF2i)) && (! shortPip_fsm_done));
  assign _zz_shortPip_fsm_shift_by = (12'h81e - shortPip_input_payload_rs1_exponent);
  assign _zz_shortPip_fsm_shift_by_1 = 6'h21;
  assign shortPip_input_isStall = (shortPip_input_valid && (! shortPip_input_ready));
  assign when_FpuCore_l672 = (! shortPip_input_isStall);
  always @(*) begin
    shortPip_mantissaForced = 1'b0;
    if(shortPip_input_payload_rs1_special) begin
      case(switch_FpuCore_l686)
        2'b00 : begin
          shortPip_mantissaForced = 1'b1;
        end
        2'b01 : begin
          shortPip_mantissaForced = 1'b1;
        end
        2'b10 : begin
          if(when_FpuCore_l702) begin
            shortPip_mantissaForced = 1'b1;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    shortPip_exponentForced = 1'b0;
    if(shortPip_input_payload_rs1_special) begin
      case(switch_FpuCore_l686)
        2'b00 : begin
          shortPip_exponentForced = 1'b1;
        end
        2'b01 : begin
          shortPip_exponentForced = 1'b1;
        end
        2'b10 : begin
          shortPip_exponentForced = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(shortPip_isSubnormal) begin
      shortPip_exponentForced = 1'b1;
    end
  end

  always @(*) begin
    shortPip_mantissaForcedValue = 1'bx;
    if(shortPip_input_payload_rs1_special) begin
      case(switch_FpuCore_l686)
        2'b00 : begin
          shortPip_mantissaForcedValue = 1'b0;
        end
        2'b01 : begin
          shortPip_mantissaForcedValue = 1'b0;
        end
        2'b10 : begin
          if(when_FpuCore_l702) begin
            shortPip_mantissaForcedValue = 1'b0;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    shortPip_exponentForcedValue = 1'bx;
    if(shortPip_input_payload_rs1_special) begin
      case(switch_FpuCore_l686)
        2'b00 : begin
          shortPip_exponentForcedValue = 1'b0;
        end
        2'b01 : begin
          shortPip_exponentForcedValue = 1'b1;
        end
        2'b10 : begin
          shortPip_exponentForcedValue = 1'b1;
        end
        default : begin
        end
      endcase
    end
    if(shortPip_isSubnormal) begin
      shortPip_exponentForcedValue = 1'b0;
    end
  end

  always @(*) begin
    shortPip_cononicalForced = 1'b0;
    if(shortPip_input_payload_rs1_special) begin
      case(switch_FpuCore_l686)
        2'b10 : begin
          if(when_FpuCore_l702) begin
            shortPip_cononicalForced = 1'b1;
          end
        end
        default : begin
        end
      endcase
    end
  end

  assign switch_FpuCore_l686 = shortPip_input_payload_rs1_exponent[1 : 0];
  assign when_FpuCore_l702 = shortPip_input_payload_rs1_exponent[2];
  assign when_FpuCore_l31_2 = (shortPip_input_payload_format == FpuFormat_DOUBLE);
  assign when_FpuCore_l31_3 = (shortPip_input_payload_format == FpuFormat_DOUBLE);
  assign when_FpuCore_l31_4 = (shortPip_input_payload_format == FpuFormat_DOUBLE);
  assign when_FpuCore_l31_5 = (shortPip_input_payload_format == FpuFormat_DOUBLE);
  always @(*) begin
    shortPip_rspNv = 1'b0;
    if(!shortPip_f2i_isZero) begin
      if(when_FpuCore_l767) begin
        shortPip_rspNv = (((shortPip_input_valid && (shortPip_input_payload_opcode == FpuOpcode_F2I)) && shortPip_fsm_done) && (! shortPip_f2i_isZero));
      end
    end
    if(shortPip_NV) begin
      shortPip_rspNv = 1'b1;
    end
  end

  always @(*) begin
    shortPip_rspNx = 1'b0;
    if(!shortPip_f2i_isZero) begin
      if(!when_FpuCore_l767) begin
        shortPip_rspNx = (((shortPip_input_valid && (shortPip_input_payload_opcode == FpuOpcode_F2I)) && shortPip_fsm_done) && (shortPip_f2i_round != 2'b00));
      end
    end
  end

  assign shortPip_f2i_unsigned = (shortPip_fsm_shift_output[32 : 0] >>> 1'd1);
  assign shortPip_f2i_resign = (shortPip_input_payload_arg[0] && shortPip_input_payload_rs1_sign);
  assign shortPip_f2i_round = {shortPip_fsm_shift_output[0],shortPip_fsm_shift_scrap};
  always @(*) begin
    case(shortPip_input_payload_roundMode)
      FpuRoundMode_RNE : begin
        shortPip_f2i_increment = (shortPip_f2i_round[1] && (shortPip_f2i_round[0] || shortPip_f2i_unsigned[0]));
      end
      FpuRoundMode_RTZ : begin
        shortPip_f2i_increment = 1'b0;
      end
      FpuRoundMode_RDN : begin
        shortPip_f2i_increment = ((shortPip_f2i_round != 2'b00) && shortPip_input_payload_rs1_sign);
      end
      FpuRoundMode_RUP : begin
        shortPip_f2i_increment = ((shortPip_f2i_round != 2'b00) && (! shortPip_input_payload_rs1_sign));
      end
      default : begin
        shortPip_f2i_increment = shortPip_f2i_round[1];
      end
    endcase
  end

  always @(*) begin
    shortPip_f2i_result = ((shortPip_f2i_resign ? (~ shortPip_f2i_unsigned) : shortPip_f2i_unsigned) + _zz_shortPip_f2i_result);
    if(shortPip_f2i_isZero) begin
      shortPip_f2i_result = 32'h0;
    end else begin
      if(when_FpuCore_l767) begin
        shortPip_f2i_result = (shortPip_f2i_overflow ? 32'hffffffff : 32'h0);
        shortPip_f2i_result[31] = (shortPip_input_payload_arg[0] ^ shortPip_f2i_overflow);
      end
    end
  end

  always @(*) begin
    shortPip_f2i_overflow = (((((shortPip_input_payload_arg[0] ? 12'h81d : 12'h81e) < shortPip_input_payload_rs1_exponent) || (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b01))) && (! shortPip_input_payload_rs1_sign)) || (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10)));
    if(when_FpuCore_l763) begin
      shortPip_f2i_overflow = 1'b1;
    end
  end

  assign shortPip_f2i_underflow = (((((12'h81e < shortPip_input_payload_rs1_exponent) || ((shortPip_input_payload_arg[0] && shortPip_f2i_unsigned[31]) && ((_zz_shortPip_f2i_underflow != _zz_shortPip_f2i_underflow_1) || shortPip_f2i_increment))) || ((! shortPip_input_payload_arg[0]) && ((shortPip_f2i_unsigned != 32'h0) || shortPip_f2i_increment))) || (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b01))) && shortPip_input_payload_rs1_sign);
  assign shortPip_f2i_isZero = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b00));
  assign when_FpuCore_l763 = ((((! shortPip_input_payload_rs1_sign) && shortPip_f2i_increment) && (&shortPip_f2i_unsigned[30 : 0])) && (shortPip_input_payload_arg[0] || shortPip_f2i_unsigned[31]));
  assign when_FpuCore_l767 = (shortPip_f2i_underflow || shortPip_f2i_overflow);
  assign shortPip_bothZero = ((shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b00)) && (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b00)));
  always @(*) begin
    shortPip_rs1Equal = ((((shortPip_input_payload_rs1_mantissa == shortPip_input_payload_rs2_mantissa) && (shortPip_input_payload_rs1_exponent == shortPip_input_payload_rs2_exponent)) && (shortPip_input_payload_rs1_sign == shortPip_input_payload_rs2_sign)) && (shortPip_input_payload_rs1_special == shortPip_input_payload_rs2_special));
    if(when_FpuCore_l784) begin
      shortPip_rs1Equal = 1'b1;
    end
  end

  always @(*) begin
    shortPip_rs1AbsSmaller = ({shortPip_input_payload_rs1_exponent,shortPip_input_payload_rs1_mantissa} < {shortPip_input_payload_rs2_exponent,shortPip_input_payload_rs2_mantissa});
    if(when_FpuCore_l780) begin
      shortPip_rs1AbsSmaller = 1'b1;
    end
    if(when_FpuCore_l781) begin
      shortPip_rs1AbsSmaller = 1'b1;
    end
    if(when_FpuCore_l782) begin
      shortPip_rs1AbsSmaller = 1'b0;
    end
    if(when_FpuCore_l783) begin
      shortPip_rs1AbsSmaller = 1'b0;
    end
  end

  assign when_FpuCore_l780 = (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b01));
  assign when_FpuCore_l781 = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b00));
  assign when_FpuCore_l782 = (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b00));
  assign when_FpuCore_l783 = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b01));
  assign when_FpuCore_l784 = (((shortPip_input_payload_rs1_sign == shortPip_input_payload_rs2_sign) && (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b01))) && (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b01)));
  assign switch_Misc_l241 = {shortPip_input_payload_rs1_sign,shortPip_input_payload_rs2_sign};
  always @(*) begin
    case(switch_Misc_l241)
      2'b00 : begin
        shortPip_rs1Smaller = shortPip_rs1AbsSmaller;
      end
      2'b01 : begin
        shortPip_rs1Smaller = 1'b0;
      end
      2'b10 : begin
        shortPip_rs1Smaller = 1'b1;
      end
      default : begin
        shortPip_rs1Smaller = ((! shortPip_rs1AbsSmaller) && (! shortPip_rs1Equal));
      end
    endcase
  end

  assign shortPip_minMaxSelectRs2 = (! (((shortPip_rs1Smaller ^ shortPip_input_payload_arg[0]) && (! (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10)))) || (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b10))));
  assign shortPip_minMaxSelectNanQuiet = ((shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10)) && (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b10)));
  always @(*) begin
    shortPip_cmpResult = (((shortPip_rs1Smaller && (! shortPip_bothZero)) && (! shortPip_input_payload_arg[1])) || ((shortPip_rs1Equal || shortPip_bothZero) && (! shortPip_input_payload_arg[0])));
    if(when_FpuCore_l796) begin
      shortPip_cmpResult = 1'b0;
    end
  end

  assign when_FpuCore_l796 = ((shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10)) || (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b10)));
  assign shortPip_sgnjRs1Sign = shortPip_input_payload_rs1_sign;
  always @(*) begin
    shortPip_sgnjRs2Sign = shortPip_input_payload_rs2_sign;
    if(when_FpuCore_l800) begin
      shortPip_sgnjRs2Sign = 1'b1;
    end
  end

  assign when_FpuCore_l800 = (shortPip_input_payload_rs2Boxed && (shortPip_input_payload_format == FpuFormat_DOUBLE));
  assign shortPip_sgnjResult = (((shortPip_sgnjRs1Sign && shortPip_input_payload_arg[1]) ^ shortPip_sgnjRs2Sign) ^ shortPip_input_payload_arg[0]);
  always @(*) begin
    shortPip_fclassResult = 32'h0;
    shortPip_fclassResult[0] = (shortPip_input_payload_rs1_sign && shortPip_decoded_isInfinity);
    shortPip_fclassResult[1] = (shortPip_input_payload_rs1_sign && shortPip_isNormal);
    shortPip_fclassResult[2] = (shortPip_input_payload_rs1_sign && shortPip_isSubnormal);
    shortPip_fclassResult[3] = (shortPip_input_payload_rs1_sign && shortPip_decoded_isZero);
    shortPip_fclassResult[4] = ((! shortPip_input_payload_rs1_sign) && shortPip_decoded_isZero);
    shortPip_fclassResult[5] = ((! shortPip_input_payload_rs1_sign) && shortPip_isSubnormal);
    shortPip_fclassResult[6] = ((! shortPip_input_payload_rs1_sign) && shortPip_isNormal);
    shortPip_fclassResult[7] = ((! shortPip_input_payload_rs1_sign) && shortPip_decoded_isInfinity);
    shortPip_fclassResult[8] = (shortPip_decoded_isNan && (! shortPip_decoded_isQuiet));
    shortPip_fclassResult[9] = (shortPip_decoded_isNan && shortPip_decoded_isQuiet);
  end

  assign shortPip_decoded_isZero = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b00));
  assign shortPip_decoded_isNormal = (! shortPip_input_payload_rs1_special);
  assign shortPip_decoded_isInfinity = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b01));
  assign shortPip_decoded_isNan = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10));
  assign shortPip_decoded_isQuiet = shortPip_input_payload_rs1_mantissa[51];
  assign shortPip_rfOutput_valid = ((shortPip_input_valid && shortPip_toFpuRf) && (! shortPip_halt));
  assign shortPip_rfOutput_payload_source = shortPip_input_payload_source;
  assign shortPip_rfOutput_payload_rd = shortPip_input_payload_rd;
  assign shortPip_rfOutput_payload_roundMode = shortPip_input_payload_roundMode;
  always @(*) begin
    shortPip_rfOutput_payload_format = shortPip_input_payload_format;
    case(shortPip_input_payload_opcode)
      FpuOpcode_SGNJ : begin
        if(when_FpuCore_l853) begin
          shortPip_rfOutput_payload_format = FpuFormat_FLOAT;
        end
      end
      FpuOpcode_FCVT_X_X : begin
        shortPip_rfOutput_payload_format = _zz_shortPip_rfOutput_payload_format;
      end
      default : begin
      end
    endcase
  end

  assign shortPip_rfOutput_payload_scrap = 1'b0;
  always @(*) begin
    shortPip_rfOutput_payload_value_sign = shortPip_input_payload_rs1_sign;
    case(shortPip_input_payload_opcode)
      FpuOpcode_MIN_MAX : begin
        if(shortPip_minMaxSelectRs2) begin
          shortPip_rfOutput_payload_value_sign = shortPip_input_payload_rs2_sign;
        end
      end
      FpuOpcode_SGNJ : begin
        if(when_FpuCore_l850) begin
          shortPip_rfOutput_payload_value_sign = shortPip_sgnjResult;
        end
        if(when_FpuCore_l853) begin
          shortPip_rfOutput_payload_value_sign = shortPip_input_payload_rs1_sign;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    shortPip_rfOutput_payload_value_exponent = shortPip_input_payload_rs1_exponent;
    case(shortPip_input_payload_opcode)
      FpuOpcode_MIN_MAX : begin
        if(shortPip_minMaxSelectRs2) begin
          shortPip_rfOutput_payload_value_exponent = shortPip_input_payload_rs2_exponent;
        end
        if(shortPip_minMaxSelectNanQuiet) begin
          shortPip_rfOutput_payload_value_exponent[1 : 0] = 2'b10;
          shortPip_rfOutput_payload_value_exponent[2] = 1'b1;
        end
      end
      FpuOpcode_FCVT_X_X : begin
        if(when_FpuCore_l860) begin
          shortPip_rfOutput_payload_value_exponent[1 : 0] = 2'b10;
          shortPip_rfOutput_payload_value_exponent[2] = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    shortPip_rfOutput_payload_value_mantissa = {shortPip_input_payload_rs1_mantissa,1'b0};
    case(shortPip_input_payload_opcode)
      FpuOpcode_MIN_MAX : begin
        if(shortPip_minMaxSelectRs2) begin
          shortPip_rfOutput_payload_value_mantissa = {shortPip_input_payload_rs2_mantissa,1'b0};
        end
        if(shortPip_minMaxSelectNanQuiet) begin
          shortPip_rfOutput_payload_value_mantissa[52] = 1'b1;
        end
      end
      FpuOpcode_FCVT_X_X : begin
        if(when_FpuCore_l860) begin
          shortPip_rfOutput_payload_value_mantissa[52] = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    shortPip_rfOutput_payload_value_special = shortPip_input_payload_rs1_special;
    case(shortPip_input_payload_opcode)
      FpuOpcode_MIN_MAX : begin
        if(shortPip_minMaxSelectRs2) begin
          shortPip_rfOutput_payload_value_special = shortPip_input_payload_rs2_special;
        end
        if(shortPip_minMaxSelectNanQuiet) begin
          shortPip_rfOutput_payload_value_special = 1'b1;
        end
      end
      FpuOpcode_FCVT_X_X : begin
        if(when_FpuCore_l860) begin
          shortPip_rfOutput_payload_value_special = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_FpuCore_l850 = (! (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10)));
  assign when_FpuCore_l853 = (shortPip_input_payload_rs1Boxed && (shortPip_input_payload_format == FpuFormat_DOUBLE));
  assign _zz_shortPip_rfOutput_payload_format = ((shortPip_input_payload_format == FpuFormat_FLOAT) ? FpuFormat_DOUBLE : FpuFormat_FLOAT);
  assign when_FpuCore_l860 = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10));
  assign shortPip_signalQuiet = ((shortPip_input_payload_opcode == FpuOpcode_CMP) && (shortPip_input_payload_arg != 2'b10));
  assign shortPip_rs1Nan = (shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10));
  assign shortPip_rs2Nan = (shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b10));
  assign shortPip_rs1NanNv = ((shortPip_input_payload_rs1_special && (shortPip_input_payload_rs1_exponent[1 : 0] == 2'b10)) && ((! shortPip_input_payload_rs1_mantissa[51]) || shortPip_signalQuiet));
  assign shortPip_rs2NanNv = ((shortPip_input_payload_rs2_special && (shortPip_input_payload_rs2_exponent[1 : 0] == 2'b10)) && ((! shortPip_input_payload_rs2_mantissa[51]) || shortPip_signalQuiet));
  assign shortPip_NV = (((|{(shortPip_input_payload_opcode == FpuOpcode_FCVT_X_X),{(shortPip_input_payload_opcode == FpuOpcode_MIN_MAX),(shortPip_input_payload_opcode == FpuOpcode_CMP)}}) && shortPip_rs1NanNv) || ((|{(shortPip_input_payload_opcode == FpuOpcode_MIN_MAX),(shortPip_input_payload_opcode == FpuOpcode_CMP)}) && shortPip_rs2NanNv));
  assign shortPip_input_ready = ((! shortPip_halt) && (shortPip_toFpuRf ? shortPip_rfOutput_ready : _zz_shortPip_input_ready));
  assign shortPip_rspStreams_0_valid = (((shortPip_input_valid && (shortPip_input_payload_source == 1'b0)) && (! shortPip_toFpuRf)) && (! shortPip_halt));
  assign shortPip_rspStreams_0_payload_value = shortPip_result;
  assign shortPip_rspStreams_0_payload_NV = shortPip_rspNv;
  assign shortPip_rspStreams_0_payload_NX = shortPip_rspNx;
  always @(*) begin
    shortPip_rspStreams_0_ready = shortPip_rspStreams_0_m2sPipe_ready;
    if(when_Stream_l375_7) begin
      shortPip_rspStreams_0_ready = 1'b1;
    end
  end

  assign when_Stream_l375_7 = (! shortPip_rspStreams_0_m2sPipe_valid);
  assign shortPip_rspStreams_0_m2sPipe_valid = shortPip_rspStreams_0_rValid;
  assign shortPip_rspStreams_0_m2sPipe_payload_value = shortPip_rspStreams_0_rData_value;
  assign shortPip_rspStreams_0_m2sPipe_payload_NV = shortPip_rspStreams_0_rData_NV;
  assign shortPip_rspStreams_0_m2sPipe_payload_NX = shortPip_rspStreams_0_rData_NX;
  assign io_port_0_rsp_valid = shortPip_rspStreams_0_m2sPipe_valid;
  assign shortPip_rspStreams_0_m2sPipe_ready = io_port_0_rsp_ready;
  assign io_port_0_rsp_payload_value = shortPip_rspStreams_0_m2sPipe_payload_value;
  assign io_port_0_rsp_payload_NV = shortPip_rspStreams_0_m2sPipe_payload_NV;
  assign io_port_0_rsp_payload_NX = shortPip_rspStreams_0_m2sPipe_payload_NX;
  assign shortPip_rspStreams_1_valid = (((shortPip_input_valid && (shortPip_input_payload_source == 1'b1)) && (! shortPip_toFpuRf)) && (! shortPip_halt));
  assign shortPip_rspStreams_1_payload_value = shortPip_result;
  assign shortPip_rspStreams_1_payload_NV = shortPip_rspNv;
  assign shortPip_rspStreams_1_payload_NX = shortPip_rspNx;
  always @(*) begin
    shortPip_rspStreams_1_ready = shortPip_rspStreams_1_m2sPipe_ready;
    if(when_Stream_l375_8) begin
      shortPip_rspStreams_1_ready = 1'b1;
    end
  end

  assign when_Stream_l375_8 = (! shortPip_rspStreams_1_m2sPipe_valid);
  assign shortPip_rspStreams_1_m2sPipe_valid = shortPip_rspStreams_1_rValid;
  assign shortPip_rspStreams_1_m2sPipe_payload_value = shortPip_rspStreams_1_rData_value;
  assign shortPip_rspStreams_1_m2sPipe_payload_NV = shortPip_rspStreams_1_rData_NV;
  assign shortPip_rspStreams_1_m2sPipe_payload_NX = shortPip_rspStreams_1_rData_NX;
  assign io_port_1_rsp_valid = shortPip_rspStreams_1_m2sPipe_valid;
  assign shortPip_rspStreams_1_m2sPipe_ready = io_port_1_rsp_ready;
  assign io_port_1_rsp_payload_value = shortPip_rspStreams_1_m2sPipe_payload_value;
  assign io_port_1_rsp_payload_NV = shortPip_rspStreams_1_m2sPipe_payload_NV;
  assign io_port_1_rsp_payload_NX = shortPip_rspStreams_1_m2sPipe_payload_NX;
  assign shortPip_rfOutput_payload_NV = shortPip_NV;
  assign shortPip_rfOutput_payload_DZ = 1'b0;
  always @(*) begin
    decode_mul_ready = mul_preMul_input_ready;
    if(when_Stream_l375_9) begin
      decode_mul_ready = 1'b1;
    end
  end

  assign when_Stream_l375_9 = (! mul_preMul_input_valid);
  assign mul_preMul_input_valid = decode_mul_rValid;
  assign mul_preMul_input_payload_source = decode_mul_rData_source;
  assign mul_preMul_input_payload_rs1_mantissa = decode_mul_rData_rs1_mantissa;
  assign mul_preMul_input_payload_rs1_exponent = decode_mul_rData_rs1_exponent;
  assign mul_preMul_input_payload_rs1_sign = decode_mul_rData_rs1_sign;
  assign mul_preMul_input_payload_rs1_special = decode_mul_rData_rs1_special;
  assign mul_preMul_input_payload_rs2_mantissa = decode_mul_rData_rs2_mantissa;
  assign mul_preMul_input_payload_rs2_exponent = decode_mul_rData_rs2_exponent;
  assign mul_preMul_input_payload_rs2_sign = decode_mul_rData_rs2_sign;
  assign mul_preMul_input_payload_rs2_special = decode_mul_rData_rs2_special;
  assign mul_preMul_input_payload_rs3_mantissa = decode_mul_rData_rs3_mantissa;
  assign mul_preMul_input_payload_rs3_exponent = decode_mul_rData_rs3_exponent;
  assign mul_preMul_input_payload_rs3_sign = decode_mul_rData_rs3_sign;
  assign mul_preMul_input_payload_rs3_special = decode_mul_rData_rs3_special;
  assign mul_preMul_input_payload_rd = decode_mul_rData_rd;
  assign mul_preMul_input_payload_add = decode_mul_rData_add;
  assign mul_preMul_input_payload_divSqrt = decode_mul_rData_divSqrt;
  assign mul_preMul_input_payload_msb1 = decode_mul_rData_msb1;
  assign mul_preMul_input_payload_msb2 = decode_mul_rData_msb2;
  assign mul_preMul_input_payload_roundMode = decode_mul_rData_roundMode;
  assign mul_preMul_input_payload_format = decode_mul_rData_format;
  assign mul_preMul_output_valid = mul_preMul_input_valid;
  assign mul_preMul_input_ready = mul_preMul_output_ready;
  assign mul_preMul_output_payload_source = mul_preMul_input_payload_source;
  assign mul_preMul_output_payload_rs1_mantissa = mul_preMul_input_payload_rs1_mantissa;
  assign mul_preMul_output_payload_rs1_exponent = mul_preMul_input_payload_rs1_exponent;
  assign mul_preMul_output_payload_rs1_sign = mul_preMul_input_payload_rs1_sign;
  assign mul_preMul_output_payload_rs1_special = mul_preMul_input_payload_rs1_special;
  assign mul_preMul_output_payload_rs2_mantissa = mul_preMul_input_payload_rs2_mantissa;
  assign mul_preMul_output_payload_rs2_exponent = mul_preMul_input_payload_rs2_exponent;
  assign mul_preMul_output_payload_rs2_sign = mul_preMul_input_payload_rs2_sign;
  assign mul_preMul_output_payload_rs2_special = mul_preMul_input_payload_rs2_special;
  assign mul_preMul_output_payload_rs3_mantissa = mul_preMul_input_payload_rs3_mantissa;
  assign mul_preMul_output_payload_rs3_exponent = mul_preMul_input_payload_rs3_exponent;
  assign mul_preMul_output_payload_rs3_sign = mul_preMul_input_payload_rs3_sign;
  assign mul_preMul_output_payload_rs3_special = mul_preMul_input_payload_rs3_special;
  assign mul_preMul_output_payload_rd = mul_preMul_input_payload_rd;
  assign mul_preMul_output_payload_add = mul_preMul_input_payload_add;
  assign mul_preMul_output_payload_divSqrt = mul_preMul_input_payload_divSqrt;
  assign mul_preMul_output_payload_msb1 = mul_preMul_input_payload_msb1;
  assign mul_preMul_output_payload_msb2 = mul_preMul_input_payload_msb2;
  assign mul_preMul_output_payload_roundMode = mul_preMul_input_payload_roundMode;
  assign mul_preMul_output_payload_format = mul_preMul_input_payload_format;
  assign mul_preMul_output_payload_exp = ({1'b0,mul_preMul_input_payload_rs1_exponent} + {1'b0,mul_preMul_input_payload_rs2_exponent});
  always @(*) begin
    mul_preMul_output_ready = mul_mul_input_ready;
    if(when_Stream_l375_10) begin
      mul_preMul_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_10 = (! mul_mul_input_valid);
  assign mul_mul_input_valid = mul_preMul_output_rValid;
  assign mul_mul_input_payload_source = mul_preMul_output_rData_source;
  assign mul_mul_input_payload_rs1_mantissa = mul_preMul_output_rData_rs1_mantissa;
  assign mul_mul_input_payload_rs1_exponent = mul_preMul_output_rData_rs1_exponent;
  assign mul_mul_input_payload_rs1_sign = mul_preMul_output_rData_rs1_sign;
  assign mul_mul_input_payload_rs1_special = mul_preMul_output_rData_rs1_special;
  assign mul_mul_input_payload_rs2_mantissa = mul_preMul_output_rData_rs2_mantissa;
  assign mul_mul_input_payload_rs2_exponent = mul_preMul_output_rData_rs2_exponent;
  assign mul_mul_input_payload_rs2_sign = mul_preMul_output_rData_rs2_sign;
  assign mul_mul_input_payload_rs2_special = mul_preMul_output_rData_rs2_special;
  assign mul_mul_input_payload_rs3_mantissa = mul_preMul_output_rData_rs3_mantissa;
  assign mul_mul_input_payload_rs3_exponent = mul_preMul_output_rData_rs3_exponent;
  assign mul_mul_input_payload_rs3_sign = mul_preMul_output_rData_rs3_sign;
  assign mul_mul_input_payload_rs3_special = mul_preMul_output_rData_rs3_special;
  assign mul_mul_input_payload_rd = mul_preMul_output_rData_rd;
  assign mul_mul_input_payload_add = mul_preMul_output_rData_add;
  assign mul_mul_input_payload_divSqrt = mul_preMul_output_rData_divSqrt;
  assign mul_mul_input_payload_msb1 = mul_preMul_output_rData_msb1;
  assign mul_mul_input_payload_msb2 = mul_preMul_output_rData_msb2;
  assign mul_mul_input_payload_roundMode = mul_preMul_output_rData_roundMode;
  assign mul_mul_input_payload_format = mul_preMul_output_rData_format;
  assign mul_mul_input_payload_exp = mul_preMul_output_rData_exp;
  assign mul_mul_output_valid = mul_mul_input_valid;
  assign mul_mul_input_ready = mul_mul_output_ready;
  assign mul_mul_mulA = {mul_mul_input_payload_msb1,mul_mul_input_payload_rs1_mantissa};
  assign mul_mul_mulB = {mul_mul_input_payload_msb2,mul_mul_input_payload_rs2_mantissa};
  assign mul_mul_output_payload_source = mul_mul_input_payload_source;
  assign mul_mul_output_payload_rs1_mantissa = mul_mul_input_payload_rs1_mantissa;
  assign mul_mul_output_payload_rs1_exponent = mul_mul_input_payload_rs1_exponent;
  assign mul_mul_output_payload_rs1_sign = mul_mul_input_payload_rs1_sign;
  assign mul_mul_output_payload_rs1_special = mul_mul_input_payload_rs1_special;
  assign mul_mul_output_payload_rs2_mantissa = mul_mul_input_payload_rs2_mantissa;
  assign mul_mul_output_payload_rs2_exponent = mul_mul_input_payload_rs2_exponent;
  assign mul_mul_output_payload_rs2_sign = mul_mul_input_payload_rs2_sign;
  assign mul_mul_output_payload_rs2_special = mul_mul_input_payload_rs2_special;
  assign mul_mul_output_payload_rs3_mantissa = mul_mul_input_payload_rs3_mantissa;
  assign mul_mul_output_payload_rs3_exponent = mul_mul_input_payload_rs3_exponent;
  assign mul_mul_output_payload_rs3_sign = mul_mul_input_payload_rs3_sign;
  assign mul_mul_output_payload_rs3_special = mul_mul_input_payload_rs3_special;
  assign mul_mul_output_payload_rd = mul_mul_input_payload_rd;
  assign mul_mul_output_payload_add = mul_mul_input_payload_add;
  assign mul_mul_output_payload_divSqrt = mul_mul_input_payload_divSqrt;
  assign mul_mul_output_payload_msb1 = mul_mul_input_payload_msb1;
  assign mul_mul_output_payload_msb2 = mul_mul_input_payload_msb2;
  assign mul_mul_output_payload_roundMode = mul_mul_input_payload_roundMode;
  assign mul_mul_output_payload_format = mul_mul_input_payload_format;
  assign mul_mul_output_payload_exp = mul_mul_input_payload_exp;
  assign mul_mul_output_payload_muls_0 = (mul_mul_mulA[17 : 0] * mul_mul_mulB[17 : 0]);
  assign mul_mul_output_payload_muls_1 = (mul_mul_mulA[17 : 0] * mul_mul_mulB[35 : 18]);
  assign mul_mul_output_payload_muls_2 = (mul_mul_mulA[35 : 18] * mul_mul_mulB[17 : 0]);
  assign mul_mul_output_payload_muls_3 = (mul_mul_mulA[17 : 0] * mul_mul_mulB[52 : 36]);
  assign mul_mul_output_payload_muls_4 = (mul_mul_mulA[52 : 36] * mul_mul_mulB[17 : 0]);
  assign mul_mul_output_payload_muls_5 = (mul_mul_mulA[35 : 18] * mul_mul_mulB[35 : 18]);
  assign mul_mul_output_payload_muls_6 = (mul_mul_mulA[35 : 18] * mul_mul_mulB[52 : 36]);
  assign mul_mul_output_payload_muls_7 = (mul_mul_mulA[52 : 36] * mul_mul_mulB[35 : 18]);
  assign mul_mul_output_payload_muls_8 = (mul_mul_mulA[52 : 36] * mul_mul_mulB[52 : 36]);
  always @(*) begin
    mul_mul_output_ready = mul_sum1_input_ready;
    if(when_Stream_l375_11) begin
      mul_mul_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_11 = (! mul_sum1_input_valid);
  assign mul_sum1_input_valid = mul_mul_output_rValid;
  assign mul_sum1_input_payload_source = mul_mul_output_rData_source;
  assign mul_sum1_input_payload_rs1_mantissa = mul_mul_output_rData_rs1_mantissa;
  assign mul_sum1_input_payload_rs1_exponent = mul_mul_output_rData_rs1_exponent;
  assign mul_sum1_input_payload_rs1_sign = mul_mul_output_rData_rs1_sign;
  assign mul_sum1_input_payload_rs1_special = mul_mul_output_rData_rs1_special;
  assign mul_sum1_input_payload_rs2_mantissa = mul_mul_output_rData_rs2_mantissa;
  assign mul_sum1_input_payload_rs2_exponent = mul_mul_output_rData_rs2_exponent;
  assign mul_sum1_input_payload_rs2_sign = mul_mul_output_rData_rs2_sign;
  assign mul_sum1_input_payload_rs2_special = mul_mul_output_rData_rs2_special;
  assign mul_sum1_input_payload_rs3_mantissa = mul_mul_output_rData_rs3_mantissa;
  assign mul_sum1_input_payload_rs3_exponent = mul_mul_output_rData_rs3_exponent;
  assign mul_sum1_input_payload_rs3_sign = mul_mul_output_rData_rs3_sign;
  assign mul_sum1_input_payload_rs3_special = mul_mul_output_rData_rs3_special;
  assign mul_sum1_input_payload_rd = mul_mul_output_rData_rd;
  assign mul_sum1_input_payload_add = mul_mul_output_rData_add;
  assign mul_sum1_input_payload_divSqrt = mul_mul_output_rData_divSqrt;
  assign mul_sum1_input_payload_msb1 = mul_mul_output_rData_msb1;
  assign mul_sum1_input_payload_msb2 = mul_mul_output_rData_msb2;
  assign mul_sum1_input_payload_roundMode = mul_mul_output_rData_roundMode;
  assign mul_sum1_input_payload_format = mul_mul_output_rData_format;
  assign mul_sum1_input_payload_exp = mul_mul_output_rData_exp;
  assign mul_sum1_input_payload_muls_0 = mul_mul_output_rData_muls_0;
  assign mul_sum1_input_payload_muls_1 = mul_mul_output_rData_muls_1;
  assign mul_sum1_input_payload_muls_2 = mul_mul_output_rData_muls_2;
  assign mul_sum1_input_payload_muls_3 = mul_mul_output_rData_muls_3;
  assign mul_sum1_input_payload_muls_4 = mul_mul_output_rData_muls_4;
  assign mul_sum1_input_payload_muls_5 = mul_mul_output_rData_muls_5;
  assign mul_sum1_input_payload_muls_6 = mul_mul_output_rData_muls_6;
  assign mul_sum1_input_payload_muls_7 = mul_mul_output_rData_muls_7;
  assign mul_sum1_input_payload_muls_8 = mul_mul_output_rData_muls_8;
  assign mul_sum1_sum = (_zz_mul_sum1_sum + _zz_mul_sum1_sum_4);
  assign mul_sum1_output_valid = mul_sum1_input_valid;
  assign mul_sum1_input_ready = mul_sum1_output_ready;
  assign mul_sum1_output_payload_source = mul_sum1_input_payload_source;
  assign mul_sum1_output_payload_rs1_mantissa = mul_sum1_input_payload_rs1_mantissa;
  assign mul_sum1_output_payload_rs1_exponent = mul_sum1_input_payload_rs1_exponent;
  assign mul_sum1_output_payload_rs1_sign = mul_sum1_input_payload_rs1_sign;
  assign mul_sum1_output_payload_rs1_special = mul_sum1_input_payload_rs1_special;
  assign mul_sum1_output_payload_rs2_mantissa = mul_sum1_input_payload_rs2_mantissa;
  assign mul_sum1_output_payload_rs2_exponent = mul_sum1_input_payload_rs2_exponent;
  assign mul_sum1_output_payload_rs2_sign = mul_sum1_input_payload_rs2_sign;
  assign mul_sum1_output_payload_rs2_special = mul_sum1_input_payload_rs2_special;
  assign mul_sum1_output_payload_rs3_mantissa = mul_sum1_input_payload_rs3_mantissa;
  assign mul_sum1_output_payload_rs3_exponent = mul_sum1_input_payload_rs3_exponent;
  assign mul_sum1_output_payload_rs3_sign = mul_sum1_input_payload_rs3_sign;
  assign mul_sum1_output_payload_rs3_special = mul_sum1_input_payload_rs3_special;
  assign mul_sum1_output_payload_rd = mul_sum1_input_payload_rd;
  assign mul_sum1_output_payload_add = mul_sum1_input_payload_add;
  assign mul_sum1_output_payload_divSqrt = mul_sum1_input_payload_divSqrt;
  assign mul_sum1_output_payload_msb1 = mul_sum1_input_payload_msb1;
  assign mul_sum1_output_payload_msb2 = mul_sum1_input_payload_msb2;
  assign mul_sum1_output_payload_roundMode = mul_sum1_input_payload_roundMode;
  assign mul_sum1_output_payload_format = mul_sum1_input_payload_format;
  assign mul_sum1_output_payload_exp = mul_sum1_input_payload_exp;
  assign mul_sum1_output_payload_mulC2 = mul_sum1_sum;
  assign mul_sum1_output_payload_muls2_0 = mul_sum1_input_payload_muls_4;
  assign mul_sum1_output_payload_muls2_1 = mul_sum1_input_payload_muls_5;
  assign mul_sum1_output_payload_muls2_2 = mul_sum1_input_payload_muls_6;
  assign mul_sum1_output_payload_muls2_3 = mul_sum1_input_payload_muls_7;
  assign mul_sum1_output_payload_muls2_4 = mul_sum1_input_payload_muls_8;
  always @(*) begin
    mul_sum1_output_ready = mul_sum2_input_ready;
    if(when_Stream_l375_12) begin
      mul_sum1_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_12 = (! mul_sum2_input_valid);
  assign mul_sum2_input_valid = mul_sum1_output_rValid;
  assign mul_sum2_input_payload_source = mul_sum1_output_rData_source;
  assign mul_sum2_input_payload_rs1_mantissa = mul_sum1_output_rData_rs1_mantissa;
  assign mul_sum2_input_payload_rs1_exponent = mul_sum1_output_rData_rs1_exponent;
  assign mul_sum2_input_payload_rs1_sign = mul_sum1_output_rData_rs1_sign;
  assign mul_sum2_input_payload_rs1_special = mul_sum1_output_rData_rs1_special;
  assign mul_sum2_input_payload_rs2_mantissa = mul_sum1_output_rData_rs2_mantissa;
  assign mul_sum2_input_payload_rs2_exponent = mul_sum1_output_rData_rs2_exponent;
  assign mul_sum2_input_payload_rs2_sign = mul_sum1_output_rData_rs2_sign;
  assign mul_sum2_input_payload_rs2_special = mul_sum1_output_rData_rs2_special;
  assign mul_sum2_input_payload_rs3_mantissa = mul_sum1_output_rData_rs3_mantissa;
  assign mul_sum2_input_payload_rs3_exponent = mul_sum1_output_rData_rs3_exponent;
  assign mul_sum2_input_payload_rs3_sign = mul_sum1_output_rData_rs3_sign;
  assign mul_sum2_input_payload_rs3_special = mul_sum1_output_rData_rs3_special;
  assign mul_sum2_input_payload_rd = mul_sum1_output_rData_rd;
  assign mul_sum2_input_payload_add = mul_sum1_output_rData_add;
  assign mul_sum2_input_payload_divSqrt = mul_sum1_output_rData_divSqrt;
  assign mul_sum2_input_payload_msb1 = mul_sum1_output_rData_msb1;
  assign mul_sum2_input_payload_msb2 = mul_sum1_output_rData_msb2;
  assign mul_sum2_input_payload_roundMode = mul_sum1_output_rData_roundMode;
  assign mul_sum2_input_payload_format = mul_sum1_output_rData_format;
  assign mul_sum2_input_payload_exp = mul_sum1_output_rData_exp;
  assign mul_sum2_input_payload_muls2_0 = mul_sum1_output_rData_muls2_0;
  assign mul_sum2_input_payload_muls2_1 = mul_sum1_output_rData_muls2_1;
  assign mul_sum2_input_payload_muls2_2 = mul_sum1_output_rData_muls2_2;
  assign mul_sum2_input_payload_muls2_3 = mul_sum1_output_rData_muls2_3;
  assign mul_sum2_input_payload_muls2_4 = mul_sum1_output_rData_muls2_4;
  assign mul_sum2_input_payload_mulC2 = mul_sum1_output_rData_mulC2;
  assign mul_sum2_sum = (mul_sum2_input_payload_mulC2 + _zz_mul_sum2_sum);
  assign mul_sum2_input_fire = (mul_sum2_input_valid && mul_sum2_input_ready);
  assign when_FpuCore_l221_2 = (mul_sum2_input_fire && (mul_sum2_input_payload_source == 1'b0));
  assign when_FpuCore_l221_3 = (mul_sum2_input_fire && (mul_sum2_input_payload_source == 1'b1));
  assign mul_sum2_isCommited = _zz_mul_sum2_isCommited;
  assign _zz_mul_sum2_input_ready = (! (! mul_sum2_isCommited));
  assign mul_sum2_input_ready = (mul_sum2_output_ready && _zz_mul_sum2_input_ready);
  assign mul_sum2_output_valid = (mul_sum2_input_valid && _zz_mul_sum2_input_ready);
  assign mul_sum2_output_payload_source = mul_sum2_input_payload_source;
  assign mul_sum2_output_payload_rs1_mantissa = mul_sum2_input_payload_rs1_mantissa;
  assign mul_sum2_output_payload_rs1_exponent = mul_sum2_input_payload_rs1_exponent;
  assign mul_sum2_output_payload_rs1_sign = mul_sum2_input_payload_rs1_sign;
  assign mul_sum2_output_payload_rs1_special = mul_sum2_input_payload_rs1_special;
  assign mul_sum2_output_payload_rs2_mantissa = mul_sum2_input_payload_rs2_mantissa;
  assign mul_sum2_output_payload_rs2_exponent = mul_sum2_input_payload_rs2_exponent;
  assign mul_sum2_output_payload_rs2_sign = mul_sum2_input_payload_rs2_sign;
  assign mul_sum2_output_payload_rs2_special = mul_sum2_input_payload_rs2_special;
  assign mul_sum2_output_payload_rs3_mantissa = mul_sum2_input_payload_rs3_mantissa;
  assign mul_sum2_output_payload_rs3_exponent = mul_sum2_input_payload_rs3_exponent;
  assign mul_sum2_output_payload_rs3_sign = mul_sum2_input_payload_rs3_sign;
  assign mul_sum2_output_payload_rs3_special = mul_sum2_input_payload_rs3_special;
  assign mul_sum2_output_payload_rd = mul_sum2_input_payload_rd;
  assign mul_sum2_output_payload_add = mul_sum2_input_payload_add;
  assign mul_sum2_output_payload_divSqrt = mul_sum2_input_payload_divSqrt;
  assign mul_sum2_output_payload_msb1 = mul_sum2_input_payload_msb1;
  assign mul_sum2_output_payload_msb2 = mul_sum2_input_payload_msb2;
  assign mul_sum2_output_payload_roundMode = mul_sum2_input_payload_roundMode;
  assign mul_sum2_output_payload_format = mul_sum2_input_payload_format;
  assign mul_sum2_output_payload_exp = mul_sum2_input_payload_exp;
  assign mul_sum2_output_payload_mulC = mul_sum2_sum;
  always @(*) begin
    mul_sum2_output_ready = mul_norm_input_ready;
    if(when_Stream_l375_13) begin
      mul_sum2_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_13 = (! mul_norm_input_valid);
  assign mul_norm_input_valid = mul_sum2_output_rValid;
  assign mul_norm_input_payload_source = mul_sum2_output_rData_source;
  assign mul_norm_input_payload_rs1_mantissa = mul_sum2_output_rData_rs1_mantissa;
  assign mul_norm_input_payload_rs1_exponent = mul_sum2_output_rData_rs1_exponent;
  assign mul_norm_input_payload_rs1_sign = mul_sum2_output_rData_rs1_sign;
  assign mul_norm_input_payload_rs1_special = mul_sum2_output_rData_rs1_special;
  assign mul_norm_input_payload_rs2_mantissa = mul_sum2_output_rData_rs2_mantissa;
  assign mul_norm_input_payload_rs2_exponent = mul_sum2_output_rData_rs2_exponent;
  assign mul_norm_input_payload_rs2_sign = mul_sum2_output_rData_rs2_sign;
  assign mul_norm_input_payload_rs2_special = mul_sum2_output_rData_rs2_special;
  assign mul_norm_input_payload_rs3_mantissa = mul_sum2_output_rData_rs3_mantissa;
  assign mul_norm_input_payload_rs3_exponent = mul_sum2_output_rData_rs3_exponent;
  assign mul_norm_input_payload_rs3_sign = mul_sum2_output_rData_rs3_sign;
  assign mul_norm_input_payload_rs3_special = mul_sum2_output_rData_rs3_special;
  assign mul_norm_input_payload_rd = mul_sum2_output_rData_rd;
  assign mul_norm_input_payload_add = mul_sum2_output_rData_add;
  assign mul_norm_input_payload_divSqrt = mul_sum2_output_rData_divSqrt;
  assign mul_norm_input_payload_msb1 = mul_sum2_output_rData_msb1;
  assign mul_norm_input_payload_msb2 = mul_sum2_output_rData_msb2;
  assign mul_norm_input_payload_roundMode = mul_sum2_output_rData_roundMode;
  assign mul_norm_input_payload_format = mul_sum2_output_rData_format;
  assign mul_norm_input_payload_exp = mul_sum2_output_rData_exp;
  assign mul_norm_input_payload_mulC = mul_sum2_output_rData_mulC;
  assign mul_norm_mulHigh = mul_norm_input_payload_mulC[105 : 51];
  assign mul_norm_mulLow = mul_norm_input_payload_mulC[50 : 0];
  always @(*) begin
    mul_norm_scrap = (mul_norm_mulLow != 51'h0);
    if(when_FpuCore_l967) begin
      mul_norm_scrap = 1'b1;
    end
  end

  assign mul_norm_needShift = mul_norm_mulHigh[54];
  assign mul_norm_exp = (mul_norm_input_payload_exp + _zz_mul_norm_exp);
  assign mul_norm_man = (mul_norm_needShift ? mul_norm_mulHigh[53 : 1] : mul_norm_mulHigh[52 : 0]);
  assign when_FpuCore_l967 = (mul_norm_needShift && mul_norm_mulHigh[0]);
  assign mul_norm_forceZero = ((mul_norm_input_payload_rs1_special && (mul_norm_input_payload_rs1_exponent[1 : 0] == 2'b00)) || (mul_norm_input_payload_rs2_special && (mul_norm_input_payload_rs2_exponent[1 : 0] == 2'b00)));
  assign mul_norm_underflowThreshold = ((mul_norm_input_payload_format == FpuFormat_DOUBLE) ? 12'hbca : 12'hf67);
  assign mul_norm_underflowExp = ((mul_norm_input_payload_format == FpuFormat_DOUBLE) ? 11'h3ca : 11'h767);
  assign mul_norm_forceUnderflow = (mul_norm_exp < _zz_mul_norm_forceUnderflow);
  assign mul_norm_forceOverflow = ((mul_norm_input_payload_rs1_special && (mul_norm_input_payload_rs1_exponent[1 : 0] == 2'b01)) || (mul_norm_input_payload_rs2_special && (mul_norm_input_payload_rs2_exponent[1 : 0] == 2'b01)));
  assign mul_norm_infinitynan = (((mul_norm_input_payload_rs1_special && (mul_norm_input_payload_rs1_exponent[1 : 0] == 2'b01)) || (mul_norm_input_payload_rs2_special && (mul_norm_input_payload_rs2_exponent[1 : 0] == 2'b01))) && ((mul_norm_input_payload_rs1_special && (mul_norm_input_payload_rs1_exponent[1 : 0] == 2'b00)) || (mul_norm_input_payload_rs2_special && (mul_norm_input_payload_rs2_exponent[1 : 0] == 2'b00))));
  assign mul_norm_forceNan = (((mul_norm_input_payload_rs1_special && (mul_norm_input_payload_rs1_exponent[1 : 0] == 2'b10)) || (mul_norm_input_payload_rs2_special && (mul_norm_input_payload_rs2_exponent[1 : 0] == 2'b10))) || mul_norm_infinitynan);
  assign mul_norm_output_sign = (mul_norm_input_payload_rs1_sign ^ mul_norm_input_payload_rs2_sign);
  always @(*) begin
    mul_norm_output_exponent = _zz_mul_norm_output_exponent[11:0];
    if(when_FpuCore_l983) begin
      mul_norm_output_exponent[11 : 10] = 2'b11;
    end
    if(mul_norm_forceNan) begin
      mul_norm_output_exponent[1 : 0] = 2'b10;
      mul_norm_output_exponent[2] = 1'b1;
    end else begin
      if(mul_norm_forceOverflow) begin
        mul_norm_output_exponent[1 : 0] = 2'b01;
      end else begin
        if(mul_norm_forceZero) begin
          mul_norm_output_exponent[1 : 0] = 2'b00;
        end else begin
          if(mul_norm_forceUnderflow) begin
            mul_norm_output_exponent = {1'd0, mul_norm_underflowExp};
          end
        end
      end
    end
  end

  always @(*) begin
    mul_norm_output_mantissa = mul_norm_man;
    if(mul_norm_forceNan) begin
      mul_norm_output_mantissa[52] = 1'b1;
    end
  end

  always @(*) begin
    mul_norm_output_special = 1'b0;
    if(mul_norm_forceNan) begin
      mul_norm_output_special = 1'b1;
    end else begin
      if(mul_norm_forceOverflow) begin
        mul_norm_output_special = 1'b1;
      end else begin
        if(mul_norm_forceZero) begin
          mul_norm_output_special = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    mul_norm_NV = 1'b0;
    if(mul_norm_forceNan) begin
      if(when_FpuCore_l987) begin
        mul_norm_NV = 1'b1;
      end
    end
  end

  assign when_FpuCore_l983 = (3'b101 <= mul_norm_exp[12 : 10]);
  assign when_FpuCore_l987 = ((mul_norm_infinitynan || ((mul_norm_input_payload_rs1_special && (mul_norm_input_payload_rs1_exponent[1 : 0] == 2'b10)) && (! mul_norm_input_payload_rs1_mantissa[51]))) || ((mul_norm_input_payload_rs2_special && (mul_norm_input_payload_rs2_exponent[1 : 0] == 2'b10)) && (! mul_norm_input_payload_rs2_mantissa[51])));
  assign mul_result_notMul_output_valid = (mul_norm_input_valid && mul_norm_input_payload_divSqrt);
  assign mul_result_notMul_output_payload = mul_norm_input_payload_mulC[104 : 52];
  assign mul_result_output_valid = ((mul_norm_input_valid && (! mul_norm_input_payload_add)) && (! mul_norm_input_payload_divSqrt));
  assign mul_result_output_payload_source = mul_norm_input_payload_source;
  assign mul_result_output_payload_rd = mul_norm_input_payload_rd;
  assign mul_result_output_payload_format = mul_norm_input_payload_format;
  assign mul_result_output_payload_roundMode = mul_norm_input_payload_roundMode;
  assign mul_result_output_payload_scrap = mul_norm_scrap;
  assign mul_result_output_payload_value_mantissa = mul_norm_output_mantissa;
  assign mul_result_output_payload_value_exponent = mul_norm_output_exponent;
  assign mul_result_output_payload_value_sign = mul_norm_output_sign;
  assign mul_result_output_payload_value_special = mul_norm_output_special;
  assign mul_result_output_payload_NV = mul_norm_NV;
  assign mul_result_output_payload_DZ = 1'b0;
  always @(*) begin
    mul_result_mulToAdd_ready = mul_result_mulToAdd_m2sPipe_ready;
    if(when_Stream_l375_14) begin
      mul_result_mulToAdd_ready = 1'b1;
    end
  end

  assign when_Stream_l375_14 = (! mul_result_mulToAdd_m2sPipe_valid);
  assign mul_result_mulToAdd_m2sPipe_valid = mul_result_mulToAdd_rValid;
  assign mul_result_mulToAdd_m2sPipe_payload_source = mul_result_mulToAdd_rData_source;
  assign mul_result_mulToAdd_m2sPipe_payload_rs1_mantissa = mul_result_mulToAdd_rData_rs1_mantissa;
  assign mul_result_mulToAdd_m2sPipe_payload_rs1_exponent = mul_result_mulToAdd_rData_rs1_exponent;
  assign mul_result_mulToAdd_m2sPipe_payload_rs1_sign = mul_result_mulToAdd_rData_rs1_sign;
  assign mul_result_mulToAdd_m2sPipe_payload_rs1_special = mul_result_mulToAdd_rData_rs1_special;
  assign mul_result_mulToAdd_m2sPipe_payload_rs2_mantissa = mul_result_mulToAdd_rData_rs2_mantissa;
  assign mul_result_mulToAdd_m2sPipe_payload_rs2_exponent = mul_result_mulToAdd_rData_rs2_exponent;
  assign mul_result_mulToAdd_m2sPipe_payload_rs2_sign = mul_result_mulToAdd_rData_rs2_sign;
  assign mul_result_mulToAdd_m2sPipe_payload_rs2_special = mul_result_mulToAdd_rData_rs2_special;
  assign mul_result_mulToAdd_m2sPipe_payload_rd = mul_result_mulToAdd_rData_rd;
  assign mul_result_mulToAdd_m2sPipe_payload_roundMode = mul_result_mulToAdd_rData_roundMode;
  assign mul_result_mulToAdd_m2sPipe_payload_format = mul_result_mulToAdd_rData_format;
  assign mul_result_mulToAdd_m2sPipe_payload_needCommit = mul_result_mulToAdd_rData_needCommit;
  assign decode_mulToAdd_valid = mul_result_mulToAdd_m2sPipe_valid;
  assign mul_result_mulToAdd_m2sPipe_ready = decode_mulToAdd_ready;
  assign decode_mulToAdd_payload_source = mul_result_mulToAdd_m2sPipe_payload_source;
  assign decode_mulToAdd_payload_rs1_mantissa = mul_result_mulToAdd_m2sPipe_payload_rs1_mantissa;
  assign decode_mulToAdd_payload_rs1_exponent = mul_result_mulToAdd_m2sPipe_payload_rs1_exponent;
  assign decode_mulToAdd_payload_rs1_sign = mul_result_mulToAdd_m2sPipe_payload_rs1_sign;
  assign decode_mulToAdd_payload_rs1_special = mul_result_mulToAdd_m2sPipe_payload_rs1_special;
  assign decode_mulToAdd_payload_rs2_mantissa = mul_result_mulToAdd_m2sPipe_payload_rs2_mantissa;
  assign decode_mulToAdd_payload_rs2_exponent = mul_result_mulToAdd_m2sPipe_payload_rs2_exponent;
  assign decode_mulToAdd_payload_rs2_sign = mul_result_mulToAdd_m2sPipe_payload_rs2_sign;
  assign decode_mulToAdd_payload_rs2_special = mul_result_mulToAdd_m2sPipe_payload_rs2_special;
  assign decode_mulToAdd_payload_rd = mul_result_mulToAdd_m2sPipe_payload_rd;
  assign decode_mulToAdd_payload_roundMode = mul_result_mulToAdd_m2sPipe_payload_roundMode;
  assign decode_mulToAdd_payload_format = mul_result_mulToAdd_m2sPipe_payload_format;
  assign decode_mulToAdd_payload_needCommit = mul_result_mulToAdd_m2sPipe_payload_needCommit;
  assign mul_result_mulToAdd_valid = (mul_norm_input_valid && mul_norm_input_payload_add);
  assign mul_result_mulToAdd_payload_source = mul_norm_input_payload_source;
  always @(*) begin
    mul_result_mulToAdd_payload_rs1_mantissa = {mul_norm_output_mantissa,mul_norm_scrap};
    if(mul_norm_NV) begin
      mul_result_mulToAdd_payload_rs1_mantissa[53] = 1'b0;
    end
  end

  assign mul_result_mulToAdd_payload_rs1_exponent = mul_norm_output_exponent;
  assign mul_result_mulToAdd_payload_rs1_sign = mul_norm_output_sign;
  assign mul_result_mulToAdd_payload_rs1_special = mul_norm_output_special;
  assign mul_result_mulToAdd_payload_rs2_exponent = mul_norm_input_payload_rs3_exponent;
  assign mul_result_mulToAdd_payload_rs2_sign = mul_norm_input_payload_rs3_sign;
  assign mul_result_mulToAdd_payload_rs2_special = mul_norm_input_payload_rs3_special;
  assign mul_result_mulToAdd_payload_rs2_mantissa = ({2'd0,mul_norm_input_payload_rs3_mantissa} <<< 2'd2);
  assign mul_result_mulToAdd_payload_rd = mul_norm_input_payload_rd;
  assign mul_result_mulToAdd_payload_roundMode = mul_norm_input_payload_roundMode;
  assign mul_result_mulToAdd_payload_needCommit = 1'b0;
  assign mul_result_mulToAdd_payload_format = mul_norm_input_payload_format;
  assign mul_norm_input_ready = ((mul_norm_input_payload_add ? mul_result_mulToAdd_ready : mul_result_output_ready) || mul_norm_input_payload_divSqrt);
  assign div_input_fire = (div_input_valid && div_input_ready);
  assign decode_div_ready = (! decode_div_rValid);
  assign div_input_valid = decode_div_rValid;
  assign div_input_payload_source = decode_div_rData_source;
  assign div_input_payload_rs1_mantissa = decode_div_rData_rs1_mantissa;
  assign div_input_payload_rs1_exponent = decode_div_rData_rs1_exponent;
  assign div_input_payload_rs1_sign = decode_div_rData_rs1_sign;
  assign div_input_payload_rs1_special = decode_div_rData_rs1_special;
  assign div_input_payload_rs2_mantissa = decode_div_rData_rs2_mantissa;
  assign div_input_payload_rs2_exponent = decode_div_rData_rs2_exponent;
  assign div_input_payload_rs2_sign = decode_div_rData_rs2_sign;
  assign div_input_payload_rs2_special = decode_div_rData_rs2_special;
  assign div_input_payload_rd = decode_div_rData_rd;
  assign div_input_payload_roundMode = decode_div_rData_roundMode;
  assign div_input_payload_format = decode_div_rData_format;
  always @(*) begin
    div_haltIt = 1'b1;
    if(div_divider_io_output_valid) begin
      div_haltIt = 1'b0;
    end
  end

  assign when_FpuCore_l221_4 = (div_input_fire && (div_input_payload_source == 1'b0));
  assign when_FpuCore_l221_5 = (div_input_fire && (div_input_payload_source == 1'b1));
  assign _zz_div_input_ready = (! (div_haltIt || (! div_isCommited)));
  assign div_input_ready = (div_output_ready && _zz_div_input_ready);
  assign div_output_valid = (div_input_valid && _zz_div_input_ready);
  assign div_dividerResult = div_divider_io_output_payload_result;
  assign div_dividerScrap = ((div_divider_io_output_payload_remain != 53'h0) || 1'b0);
  assign div_divider_io_input_fire = (div_divider_io_input_valid && div_divider_io_input_ready);
  assign when_FpuCore_l1056 = (! div_haltIt);
  assign div_divider_io_input_valid = (div_input_valid && (! div_cmdSent));
  assign div_output_payload_source = div_input_payload_source;
  assign div_output_payload_rd = div_input_payload_rd;
  assign div_output_payload_roundMode = div_input_payload_roundMode;
  assign div_output_payload_format = div_input_payload_format;
  assign div_needShift = (! div_dividerResult[54]);
  assign div_mantissa = (div_needShift ? div_dividerResult[52 : 0] : div_dividerResult[53 : 1]);
  assign div_scrap = (div_dividerScrap || ((! div_needShift) && div_dividerResult[0]));
  assign div_exponent = (_zz_div_exponent - _zz_div_exponent_4);
  always @(*) begin
    div_output_payload_value_special = 1'b0;
    if(div_forceNan) begin
      div_output_payload_value_special = 1'b1;
    end else begin
      if(div_forceOverflow) begin
        div_output_payload_value_special = 1'b1;
      end else begin
        if(div_forceZero) begin
          div_output_payload_value_special = 1'b1;
        end
      end
    end
  end

  assign div_output_payload_value_sign = (div_input_payload_rs1_sign ^ div_input_payload_rs2_sign);
  always @(*) begin
    div_output_payload_value_exponent = div_exponent[11:0];
    if(when_FpuCore_l1072) begin
      div_output_payload_value_exponent[11 : 9] = 3'b111;
    end
    if(when_FpuCore_l1089) begin
      div_output_payload_value_exponent[11 : 10] = 2'b11;
    end
    if(div_forceNan) begin
      div_output_payload_value_exponent[1 : 0] = 2'b10;
      div_output_payload_value_exponent[2] = 1'b1;
    end else begin
      if(div_forceOverflow) begin
        div_output_payload_value_exponent[1 : 0] = 2'b01;
      end else begin
        if(div_forceZero) begin
          div_output_payload_value_exponent[1 : 0] = 2'b00;
        end else begin
          if(div_forceUnderflow) begin
            div_output_payload_value_exponent = div_underflowExp[11:0];
          end
        end
      end
    end
  end

  always @(*) begin
    div_output_payload_value_mantissa = div_mantissa;
    if(div_forceNan) begin
      div_output_payload_value_mantissa[52] = 1'b1;
    end
  end

  assign div_output_payload_scrap = div_scrap;
  assign when_FpuCore_l1072 = (div_exponent[13 : 12] == 2'b11);
  assign div_underflowThreshold = ((div_input_payload_format == FpuFormat_DOUBLE) ? 14'h23cb : 14'h2768);
  assign div_underflowExp = ((div_input_payload_format == FpuFormat_DOUBLE) ? 14'h23ca : 14'h2767);
  assign div_forceUnderflow = (div_exponent < div_underflowThreshold);
  assign div_forceOverflow = ((div_input_payload_rs1_special && (div_input_payload_rs1_exponent[1 : 0] == 2'b01)) || (div_input_payload_rs2_special && (div_input_payload_rs2_exponent[1 : 0] == 2'b00)));
  assign div_infinitynan = (((div_input_payload_rs1_special && (div_input_payload_rs1_exponent[1 : 0] == 2'b00)) && (div_input_payload_rs2_special && (div_input_payload_rs2_exponent[1 : 0] == 2'b00))) || ((div_input_payload_rs1_special && (div_input_payload_rs1_exponent[1 : 0] == 2'b01)) && (div_input_payload_rs2_special && (div_input_payload_rs2_exponent[1 : 0] == 2'b01))));
  assign div_forceNan = (((div_input_payload_rs1_special && (div_input_payload_rs1_exponent[1 : 0] == 2'b10)) || (div_input_payload_rs2_special && (div_input_payload_rs2_exponent[1 : 0] == 2'b10))) || div_infinitynan);
  assign div_forceZero = ((div_input_payload_rs1_special && (div_input_payload_rs1_exponent[1 : 0] == 2'b00)) || (div_input_payload_rs2_special && (div_input_payload_rs2_exponent[1 : 0] == 2'b01)));
  always @(*) begin
    div_output_payload_NV = 1'b0;
    if(div_forceNan) begin
      if(when_FpuCore_l1093) begin
        div_output_payload_NV = 1'b1;
      end
    end
  end

  assign div_output_payload_DZ = (((! div_forceNan) && (! (div_input_payload_rs1_special && (div_input_payload_rs1_exponent[1 : 0] == 2'b01)))) && (div_input_payload_rs2_special && (div_input_payload_rs2_exponent[1 : 0] == 2'b00)));
  assign when_FpuCore_l1089 = (div_exponent[13 : 11] == 3'b111);
  assign when_FpuCore_l1093 = ((div_infinitynan || ((div_input_payload_rs1_special && (div_input_payload_rs1_exponent[1 : 0] == 2'b10)) && (! div_input_payload_rs1_mantissa[51]))) || ((div_input_payload_rs2_special && (div_input_payload_rs2_exponent[1 : 0] == 2'b10)) && (! div_input_payload_rs2_mantissa[51])));
  assign sqrt_input_fire = (sqrt_input_valid && sqrt_input_ready);
  assign decode_sqrt_ready = (! decode_sqrt_rValid);
  assign sqrt_input_valid = decode_sqrt_rValid;
  assign sqrt_input_payload_source = decode_sqrt_rData_source;
  assign sqrt_input_payload_rs1_mantissa = decode_sqrt_rData_rs1_mantissa;
  assign sqrt_input_payload_rs1_exponent = decode_sqrt_rData_rs1_exponent;
  assign sqrt_input_payload_rs1_sign = decode_sqrt_rData_rs1_sign;
  assign sqrt_input_payload_rs1_special = decode_sqrt_rData_rs1_special;
  assign sqrt_input_payload_rd = decode_sqrt_rData_rd;
  assign sqrt_input_payload_roundMode = decode_sqrt_rData_roundMode;
  assign sqrt_input_payload_format = decode_sqrt_rData_format;
  always @(*) begin
    sqrt_haltIt = 1'b1;
    if(sqrt_sqrt_io_output_valid) begin
      sqrt_haltIt = 1'b0;
    end
  end

  assign when_FpuCore_l221_6 = (sqrt_input_fire && (sqrt_input_payload_source == 1'b0));
  assign when_FpuCore_l221_7 = (sqrt_input_fire && (sqrt_input_payload_source == 1'b1));
  assign _zz_sqrt_input_ready = (! (sqrt_haltIt || (! sqrt_isCommited)));
  assign sqrt_input_ready = (sqrt_output_ready && _zz_sqrt_input_ready);
  assign sqrt_output_valid = (sqrt_input_valid && _zz_sqrt_input_ready);
  assign sqrt_needShift = (! sqrt_input_payload_rs1_exponent[0]);
  assign sqrt_sqrt_io_input_payload_a = (sqrt_needShift ? {{1'b1,sqrt_input_payload_rs1_mantissa},1'b0} : {2'b01,sqrt_input_payload_rs1_mantissa});
  assign sqrt_sqrt_io_input_fire = (sqrt_sqrt_io_input_valid && sqrt_sqrt_io_input_ready);
  assign when_FpuCore_l1118 = (! sqrt_haltIt);
  assign sqrt_sqrt_io_input_valid = (sqrt_input_valid && (! sqrt_cmdSent));
  assign sqrt_output_payload_source = sqrt_input_payload_source;
  assign sqrt_output_payload_rd = sqrt_input_payload_rd;
  assign sqrt_output_payload_roundMode = sqrt_input_payload_roundMode;
  assign sqrt_output_payload_format = sqrt_input_payload_format;
  assign sqrt_scrap = (sqrt_sqrt_io_output_payload_remain != 57'h0);
  always @(*) begin
    sqrt_output_payload_value_special = 1'b0;
    if(when_FpuCore_l1137) begin
      sqrt_output_payload_value_special = 1'b1;
    end
    if(sqrt_negative) begin
      sqrt_output_payload_value_special = 1'b1;
    end
    if(when_FpuCore_l1144) begin
      sqrt_output_payload_value_special = 1'b1;
    end
    if(when_FpuCore_l1148) begin
      sqrt_output_payload_value_special = 1'b1;
    end
  end

  assign sqrt_output_payload_value_sign = sqrt_input_payload_rs1_sign;
  always @(*) begin
    sqrt_output_payload_value_exponent = sqrt_exponent;
    if(when_FpuCore_l1137) begin
      sqrt_output_payload_value_exponent[1 : 0] = 2'b01;
    end
    if(sqrt_negative) begin
      sqrt_output_payload_value_exponent[1 : 0] = 2'b10;
      sqrt_output_payload_value_exponent[2] = 1'b1;
    end
    if(when_FpuCore_l1144) begin
      sqrt_output_payload_value_exponent[1 : 0] = 2'b10;
      sqrt_output_payload_value_exponent[2] = 1'b1;
    end
    if(when_FpuCore_l1148) begin
      sqrt_output_payload_value_exponent[1 : 0] = 2'b00;
    end
  end

  always @(*) begin
    sqrt_output_payload_value_mantissa = sqrt_sqrt_io_output_payload_result;
    if(sqrt_negative) begin
      sqrt_output_payload_value_mantissa[52] = 1'b1;
    end
    if(when_FpuCore_l1144) begin
      sqrt_output_payload_value_mantissa[52] = 1'b1;
    end
  end

  assign sqrt_output_payload_scrap = sqrt_scrap;
  always @(*) begin
    sqrt_output_payload_NV = 1'b0;
    if(sqrt_negative) begin
      sqrt_output_payload_NV = 1'b1;
    end
    if(when_FpuCore_l1144) begin
      sqrt_output_payload_NV = (! sqrt_input_payload_rs1_mantissa[51]);
    end
  end

  assign sqrt_output_payload_DZ = 1'b0;
  assign sqrt_negative = (((! (sqrt_input_payload_rs1_special && (sqrt_input_payload_rs1_exponent[1 : 0] == 2'b10))) && (! (sqrt_input_payload_rs1_special && (sqrt_input_payload_rs1_exponent[1 : 0] == 2'b00)))) && sqrt_input_payload_rs1_sign);
  assign when_FpuCore_l1137 = (sqrt_input_payload_rs1_special && (sqrt_input_payload_rs1_exponent[1 : 0] == 2'b01));
  assign when_FpuCore_l1144 = (sqrt_input_payload_rs1_special && (sqrt_input_payload_rs1_exponent[1 : 0] == 2'b10));
  assign when_FpuCore_l1148 = (sqrt_input_payload_rs1_special && (sqrt_input_payload_rs1_exponent[1 : 0] == 2'b00));
  assign add_preShifter_input_valid = decode_add_valid;
  assign decode_add_ready = add_preShifter_input_ready;
  assign add_preShifter_input_payload_source = decode_add_payload_source;
  assign add_preShifter_input_payload_rs1_mantissa = decode_add_payload_rs1_mantissa;
  assign add_preShifter_input_payload_rs1_exponent = decode_add_payload_rs1_exponent;
  assign add_preShifter_input_payload_rs1_sign = decode_add_payload_rs1_sign;
  assign add_preShifter_input_payload_rs1_special = decode_add_payload_rs1_special;
  assign add_preShifter_input_payload_rs2_mantissa = decode_add_payload_rs2_mantissa;
  assign add_preShifter_input_payload_rs2_exponent = decode_add_payload_rs2_exponent;
  assign add_preShifter_input_payload_rs2_sign = decode_add_payload_rs2_sign;
  assign add_preShifter_input_payload_rs2_special = decode_add_payload_rs2_special;
  assign add_preShifter_input_payload_rd = decode_add_payload_rd;
  assign add_preShifter_input_payload_roundMode = decode_add_payload_roundMode;
  assign add_preShifter_input_payload_format = decode_add_payload_format;
  assign add_preShifter_input_payload_needCommit = decode_add_payload_needCommit;
  assign add_preShifter_output_valid = add_preShifter_input_valid;
  assign add_preShifter_input_ready = add_preShifter_output_ready;
  assign add_preShifter_exp21 = ({1'b0,add_preShifter_input_payload_rs2_exponent} - {1'b0,add_preShifter_input_payload_rs1_exponent});
  assign add_preShifter_rs1ExponentBigger = ((add_preShifter_exp21[12] || (add_preShifter_input_payload_rs2_special && (add_preShifter_input_payload_rs2_exponent[1 : 0] == 2'b00))) && (! (add_preShifter_input_payload_rs1_special && (add_preShifter_input_payload_rs1_exponent[1 : 0] == 2'b00))));
  assign add_preShifter_rs1ExponentEqual = (add_preShifter_input_payload_rs1_exponent == add_preShifter_input_payload_rs2_exponent);
  assign add_preShifter_rs1MantissaBigger = (add_preShifter_input_payload_rs2_mantissa < add_preShifter_input_payload_rs1_mantissa);
  assign add_preShifter_absRs1Bigger = ((((add_preShifter_rs1ExponentBigger || (add_preShifter_rs1ExponentEqual && add_preShifter_rs1MantissaBigger)) && (! (add_preShifter_input_payload_rs1_special && (add_preShifter_input_payload_rs1_exponent[1 : 0] == 2'b00)))) || (add_preShifter_input_payload_rs1_special && (add_preShifter_input_payload_rs1_exponent[1 : 0] == 2'b01))) && (! (add_preShifter_input_payload_rs2_special && (add_preShifter_input_payload_rs2_exponent[1 : 0] == 2'b01))));
  assign add_preShifter_output_payload_source = add_preShifter_input_payload_source;
  assign add_preShifter_output_payload_rs1_mantissa = add_preShifter_input_payload_rs1_mantissa;
  assign add_preShifter_output_payload_rs1_exponent = add_preShifter_input_payload_rs1_exponent;
  assign add_preShifter_output_payload_rs1_sign = add_preShifter_input_payload_rs1_sign;
  assign add_preShifter_output_payload_rs1_special = add_preShifter_input_payload_rs1_special;
  assign add_preShifter_output_payload_rs2_mantissa = add_preShifter_input_payload_rs2_mantissa;
  assign add_preShifter_output_payload_rs2_exponent = add_preShifter_input_payload_rs2_exponent;
  assign add_preShifter_output_payload_rs2_sign = add_preShifter_input_payload_rs2_sign;
  assign add_preShifter_output_payload_rs2_special = add_preShifter_input_payload_rs2_special;
  assign add_preShifter_output_payload_rd = add_preShifter_input_payload_rd;
  assign add_preShifter_output_payload_roundMode = add_preShifter_input_payload_roundMode;
  assign add_preShifter_output_payload_format = add_preShifter_input_payload_format;
  assign add_preShifter_output_payload_needCommit = add_preShifter_input_payload_needCommit;
  assign add_preShifter_output_payload_absRs1Bigger = add_preShifter_absRs1Bigger;
  assign add_preShifter_output_payload_rs1ExponentBigger = add_preShifter_rs1ExponentBigger;
  always @(*) begin
    add_preShifter_output_ready = add_shifter_input_ready;
    if(when_Stream_l375_15) begin
      add_preShifter_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_15 = (! add_shifter_input_valid);
  assign add_shifter_input_valid = add_preShifter_output_rValid;
  assign add_shifter_input_payload_source = add_preShifter_output_rData_source;
  assign add_shifter_input_payload_rs1_mantissa = add_preShifter_output_rData_rs1_mantissa;
  assign add_shifter_input_payload_rs1_exponent = add_preShifter_output_rData_rs1_exponent;
  assign add_shifter_input_payload_rs1_sign = add_preShifter_output_rData_rs1_sign;
  assign add_shifter_input_payload_rs1_special = add_preShifter_output_rData_rs1_special;
  assign add_shifter_input_payload_rs2_mantissa = add_preShifter_output_rData_rs2_mantissa;
  assign add_shifter_input_payload_rs2_exponent = add_preShifter_output_rData_rs2_exponent;
  assign add_shifter_input_payload_rs2_sign = add_preShifter_output_rData_rs2_sign;
  assign add_shifter_input_payload_rs2_special = add_preShifter_output_rData_rs2_special;
  assign add_shifter_input_payload_rd = add_preShifter_output_rData_rd;
  assign add_shifter_input_payload_roundMode = add_preShifter_output_rData_roundMode;
  assign add_shifter_input_payload_format = add_preShifter_output_rData_format;
  assign add_shifter_input_payload_needCommit = add_preShifter_output_rData_needCommit;
  assign add_shifter_input_payload_absRs1Bigger = add_preShifter_output_rData_absRs1Bigger;
  assign add_shifter_input_payload_rs1ExponentBigger = add_preShifter_output_rData_rs1ExponentBigger;
  assign add_shifter_output_valid = add_shifter_input_valid;
  assign add_shifter_input_ready = add_shifter_output_ready;
  assign add_shifter_output_payload_source = add_shifter_input_payload_source;
  assign add_shifter_output_payload_rs1_mantissa = add_shifter_input_payload_rs1_mantissa;
  assign add_shifter_output_payload_rs1_exponent = add_shifter_input_payload_rs1_exponent;
  assign add_shifter_output_payload_rs1_sign = add_shifter_input_payload_rs1_sign;
  assign add_shifter_output_payload_rs1_special = add_shifter_input_payload_rs1_special;
  assign add_shifter_output_payload_rs2_mantissa = add_shifter_input_payload_rs2_mantissa;
  assign add_shifter_output_payload_rs2_exponent = add_shifter_input_payload_rs2_exponent;
  assign add_shifter_output_payload_rs2_sign = add_shifter_input_payload_rs2_sign;
  assign add_shifter_output_payload_rs2_special = add_shifter_input_payload_rs2_special;
  assign add_shifter_output_payload_rd = add_shifter_input_payload_rd;
  assign add_shifter_output_payload_roundMode = add_shifter_input_payload_roundMode;
  assign add_shifter_output_payload_format = add_shifter_input_payload_format;
  assign add_shifter_output_payload_needCommit = add_shifter_input_payload_needCommit;
  assign add_shifter_exp21 = ({1'b0,add_shifter_input_payload_rs2_exponent} - {1'b0,add_shifter_input_payload_rs1_exponent});
  assign _zz_add_shifter_shiftBy = add_shifter_exp21;
  assign add_shifter_shiftBy = (_zz_add_shifter_shiftBy_1 + _zz_add_shifter_shiftBy_3);
  assign add_shifter_shiftOverflow = (13'h0037 <= add_shifter_shiftBy);
  assign add_shifter_passThrough = ((add_shifter_shiftOverflow || (add_shifter_input_payload_rs1_special && (add_shifter_input_payload_rs1_exponent[1 : 0] == 2'b00))) || (add_shifter_input_payload_rs2_special && (add_shifter_input_payload_rs2_exponent[1 : 0] == 2'b00)));
  assign add_shifter_xySign = (add_shifter_input_payload_absRs1Bigger ? add_shifter_input_payload_rs1_sign : add_shifter_input_payload_rs2_sign);
  assign add_shifter_output_payload_xSign = (add_shifter_xySign ^ (add_shifter_input_payload_rs1ExponentBigger ? add_shifter_input_payload_rs1_sign : add_shifter_input_payload_rs2_sign));
  assign add_shifter_output_payload_ySign = (add_shifter_xySign ^ (add_shifter_input_payload_rs1ExponentBigger ? add_shifter_input_payload_rs2_sign : add_shifter_input_payload_rs1_sign));
  assign add_shifter_xMantissa = {1'b1,(add_shifter_input_payload_rs1ExponentBigger ? add_shifter_input_payload_rs1_mantissa : add_shifter_input_payload_rs2_mantissa)};
  assign add_shifter_yMantissaUnshifted = {1'b1,(add_shifter_input_payload_rs1ExponentBigger ? add_shifter_input_payload_rs2_mantissa : add_shifter_input_payload_rs1_mantissa)};
  assign add_shifter_yMantissa = add_shifter_yMantissaUnshifted;
  always @(*) begin
    add_shifter_roundingScrap = 1'b0;
    if(when_FpuCore_l1419) begin
      add_shifter_roundingScrap = 1'b1;
    end
    if(when_FpuCore_l1419_1) begin
      add_shifter_roundingScrap = 1'b1;
    end
    if(when_FpuCore_l1419_2) begin
      add_shifter_roundingScrap = 1'b1;
    end
    if(when_FpuCore_l1419_3) begin
      add_shifter_roundingScrap = 1'b1;
    end
    if(when_FpuCore_l1419_4) begin
      add_shifter_roundingScrap = 1'b1;
    end
    if(when_FpuCore_l1419_5) begin
      add_shifter_roundingScrap = 1'b1;
    end
    if(add_shifter_shiftOverflow) begin
      add_shifter_roundingScrap = 1'b1;
    end
    if(when_FpuCore_l1424) begin
      add_shifter_roundingScrap = 1'b0;
    end
  end

  assign when_FpuCore_l1419 = (add_shifter_shiftBy[5] && (add_shifter_yMantissa[31 : 0] != 32'h0));
  assign when_FpuCore_l1419_1 = (add_shifter_shiftBy[4] && (add_shifter_yMantissa_1[15 : 0] != 16'h0));
  assign when_FpuCore_l1419_2 = (add_shifter_shiftBy[3] && (add_shifter_yMantissa_2[7 : 0] != 8'h0));
  assign when_FpuCore_l1419_3 = (add_shifter_shiftBy[2] && (add_shifter_yMantissa_3[3 : 0] != 4'b0000));
  assign when_FpuCore_l1419_4 = (add_shifter_shiftBy[1] && (add_shifter_yMantissa_4[1 : 0] != 2'b00));
  assign when_FpuCore_l1419_5 = (add_shifter_shiftBy[0] && (add_shifter_yMantissa_5[0 : 0] != 1'b0));
  assign when_FpuCore_l1424 = (add_shifter_input_payload_rs1_special || add_shifter_input_payload_rs2_special);
  assign add_shifter_output_payload_xyExponent = (add_shifter_input_payload_rs1ExponentBigger ? add_shifter_input_payload_rs1_exponent : add_shifter_input_payload_rs2_exponent);
  assign add_shifter_output_payload_xMantissa = add_shifter_xMantissa;
  assign add_shifter_output_payload_yMantissa = add_shifter_yMantissa_6;
  assign add_shifter_output_payload_xySign = add_shifter_xySign;
  assign add_shifter_output_payload_roundingScrap = add_shifter_roundingScrap;
  always @(*) begin
    add_shifter_output_ready = add_math_input_ready;
    if(when_Stream_l375_16) begin
      add_shifter_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_16 = (! add_math_input_valid);
  assign add_math_input_valid = add_shifter_output_rValid;
  assign add_math_input_payload_source = add_shifter_output_rData_source;
  assign add_math_input_payload_rs1_mantissa = add_shifter_output_rData_rs1_mantissa;
  assign add_math_input_payload_rs1_exponent = add_shifter_output_rData_rs1_exponent;
  assign add_math_input_payload_rs1_sign = add_shifter_output_rData_rs1_sign;
  assign add_math_input_payload_rs1_special = add_shifter_output_rData_rs1_special;
  assign add_math_input_payload_rs2_mantissa = add_shifter_output_rData_rs2_mantissa;
  assign add_math_input_payload_rs2_exponent = add_shifter_output_rData_rs2_exponent;
  assign add_math_input_payload_rs2_sign = add_shifter_output_rData_rs2_sign;
  assign add_math_input_payload_rs2_special = add_shifter_output_rData_rs2_special;
  assign add_math_input_payload_rd = add_shifter_output_rData_rd;
  assign add_math_input_payload_roundMode = add_shifter_output_rData_roundMode;
  assign add_math_input_payload_format = add_shifter_output_rData_format;
  assign add_math_input_payload_needCommit = add_shifter_output_rData_needCommit;
  assign add_math_input_payload_xSign = add_shifter_output_rData_xSign;
  assign add_math_input_payload_ySign = add_shifter_output_rData_ySign;
  assign add_math_input_payload_xMantissa = add_shifter_output_rData_xMantissa;
  assign add_math_input_payload_yMantissa = add_shifter_output_rData_yMantissa;
  assign add_math_input_payload_xyExponent = add_shifter_output_rData_xyExponent;
  assign add_math_input_payload_xySign = add_shifter_output_rData_xySign;
  assign add_math_input_payload_roundingScrap = add_shifter_output_rData_roundingScrap;
  assign add_math_output_valid = add_math_input_valid;
  assign add_math_input_ready = add_math_output_ready;
  assign add_math_output_payload_source = add_math_input_payload_source;
  assign add_math_output_payload_rs1_mantissa = add_math_input_payload_rs1_mantissa;
  assign add_math_output_payload_rs1_exponent = add_math_input_payload_rs1_exponent;
  assign add_math_output_payload_rs1_sign = add_math_input_payload_rs1_sign;
  assign add_math_output_payload_rs1_special = add_math_input_payload_rs1_special;
  assign add_math_output_payload_rs2_mantissa = add_math_input_payload_rs2_mantissa;
  assign add_math_output_payload_rs2_exponent = add_math_input_payload_rs2_exponent;
  assign add_math_output_payload_rs2_sign = add_math_input_payload_rs2_sign;
  assign add_math_output_payload_rs2_special = add_math_input_payload_rs2_special;
  assign add_math_output_payload_rd = add_math_input_payload_rd;
  assign add_math_output_payload_roundMode = add_math_input_payload_roundMode;
  assign add_math_output_payload_format = add_math_input_payload_format;
  assign add_math_output_payload_needCommit = add_math_input_payload_needCommit;
  assign add_math_output_payload_xSign = add_math_input_payload_xSign;
  assign add_math_output_payload_ySign = add_math_input_payload_ySign;
  assign add_math_output_payload_xMantissa = add_math_input_payload_xMantissa;
  assign add_math_output_payload_yMantissa = add_math_input_payload_yMantissa;
  assign add_math_output_payload_xyExponent = add_math_input_payload_xyExponent;
  assign add_math_output_payload_xySign = add_math_input_payload_xySign;
  assign add_math_output_payload_roundingScrap = add_math_input_payload_roundingScrap;
  assign add_math_xSigned = _zz_add_math_xSigned;
  assign add_math_ySigned = _zz_add_math_ySigned;
  assign add_math_output_payload_xyMantissa = _zz_add_math_output_payload_xyMantissa[55 : 0];
  always @(*) begin
    add_math_output_ready = add_oh_input_ready;
    if(when_Stream_l375_17) begin
      add_math_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_17 = (! add_oh_input_valid);
  assign add_oh_input_valid = add_math_output_rValid;
  assign add_oh_input_payload_source = add_math_output_rData_source;
  assign add_oh_input_payload_rs1_mantissa = add_math_output_rData_rs1_mantissa;
  assign add_oh_input_payload_rs1_exponent = add_math_output_rData_rs1_exponent;
  assign add_oh_input_payload_rs1_sign = add_math_output_rData_rs1_sign;
  assign add_oh_input_payload_rs1_special = add_math_output_rData_rs1_special;
  assign add_oh_input_payload_rs2_mantissa = add_math_output_rData_rs2_mantissa;
  assign add_oh_input_payload_rs2_exponent = add_math_output_rData_rs2_exponent;
  assign add_oh_input_payload_rs2_sign = add_math_output_rData_rs2_sign;
  assign add_oh_input_payload_rs2_special = add_math_output_rData_rs2_special;
  assign add_oh_input_payload_rd = add_math_output_rData_rd;
  assign add_oh_input_payload_roundMode = add_math_output_rData_roundMode;
  assign add_oh_input_payload_format = add_math_output_rData_format;
  assign add_oh_input_payload_needCommit = add_math_output_rData_needCommit;
  assign add_oh_input_payload_xSign = add_math_output_rData_xSign;
  assign add_oh_input_payload_ySign = add_math_output_rData_ySign;
  assign add_oh_input_payload_xMantissa = add_math_output_rData_xMantissa;
  assign add_oh_input_payload_yMantissa = add_math_output_rData_yMantissa;
  assign add_oh_input_payload_xyExponent = add_math_output_rData_xyExponent;
  assign add_oh_input_payload_xySign = add_math_output_rData_xySign;
  assign add_oh_input_payload_roundingScrap = add_math_output_rData_roundingScrap;
  assign add_oh_input_payload_xyMantissa = add_math_output_rData_xyMantissa;
  assign add_oh_input_fire = (add_oh_input_valid && add_oh_input_ready);
  assign _zz_when_FpuCore_l221_1 = (add_oh_input_fire && add_oh_input_payload_needCommit);
  assign when_FpuCore_l221_8 = (_zz_when_FpuCore_l221_1 && (add_oh_input_payload_source == 1'b0));
  assign when_FpuCore_l221_9 = (_zz_when_FpuCore_l221_1 && (add_oh_input_payload_source == 1'b1));
  assign add_oh_isCommited = _zz_add_oh_isCommited;
  assign _zz_add_oh_input_ready = (! (add_oh_input_payload_needCommit && (! add_oh_isCommited)));
  assign add_oh_input_ready = (add_oh_output_ready && _zz_add_oh_input_ready);
  assign add_oh_output_valid = (add_oh_input_valid && _zz_add_oh_input_ready);
  assign add_oh_output_payload_source = add_oh_input_payload_source;
  assign add_oh_output_payload_rs1_mantissa = add_oh_input_payload_rs1_mantissa;
  assign add_oh_output_payload_rs1_exponent = add_oh_input_payload_rs1_exponent;
  assign add_oh_output_payload_rs1_sign = add_oh_input_payload_rs1_sign;
  assign add_oh_output_payload_rs1_special = add_oh_input_payload_rs1_special;
  assign add_oh_output_payload_rs2_mantissa = add_oh_input_payload_rs2_mantissa;
  assign add_oh_output_payload_rs2_exponent = add_oh_input_payload_rs2_exponent;
  assign add_oh_output_payload_rs2_sign = add_oh_input_payload_rs2_sign;
  assign add_oh_output_payload_rs2_special = add_oh_input_payload_rs2_special;
  assign add_oh_output_payload_rd = add_oh_input_payload_rd;
  assign add_oh_output_payload_roundMode = add_oh_input_payload_roundMode;
  assign add_oh_output_payload_format = add_oh_input_payload_format;
  assign add_oh_output_payload_needCommit = add_oh_input_payload_needCommit;
  assign add_oh_output_payload_xSign = add_oh_input_payload_xSign;
  assign add_oh_output_payload_ySign = add_oh_input_payload_ySign;
  assign add_oh_output_payload_xMantissa = add_oh_input_payload_xMantissa;
  assign add_oh_output_payload_yMantissa = add_oh_input_payload_yMantissa;
  assign add_oh_output_payload_xyExponent = add_oh_input_payload_xyExponent;
  assign add_oh_output_payload_xySign = add_oh_input_payload_xySign;
  assign add_oh_output_payload_roundingScrap = add_oh_input_payload_roundingScrap;
  assign add_oh_output_payload_xyMantissa = add_oh_input_payload_xyMantissa;
  assign _zz_add_oh_shift = {add_oh_output_payload_xyMantissa[0],{add_oh_output_payload_xyMantissa[1],{add_oh_output_payload_xyMantissa[2],{add_oh_output_payload_xyMantissa[3],{add_oh_output_payload_xyMantissa[4],{add_oh_output_payload_xyMantissa[5],{add_oh_output_payload_xyMantissa[6],{_zz__zz_add_oh_shift,{_zz__zz_add_oh_shift_1,_zz__zz_add_oh_shift_2}}}}}}}}};
  assign _zz_add_oh_shift_1 = (_zz_add_oh_shift & (~ _zz__zz_add_oh_shift_1_1));
  assign _zz_add_oh_shift_2 = _zz_add_oh_shift_1[3];
  assign _zz_add_oh_shift_3 = _zz_add_oh_shift_1[5];
  assign _zz_add_oh_shift_4 = _zz_add_oh_shift_1[6];
  assign _zz_add_oh_shift_5 = _zz_add_oh_shift_1[7];
  assign _zz_add_oh_shift_6 = _zz_add_oh_shift_1[9];
  assign _zz_add_oh_shift_7 = _zz_add_oh_shift_1[10];
  assign _zz_add_oh_shift_8 = _zz_add_oh_shift_1[11];
  assign _zz_add_oh_shift_9 = _zz_add_oh_shift_1[12];
  assign _zz_add_oh_shift_10 = _zz_add_oh_shift_1[13];
  assign _zz_add_oh_shift_11 = _zz_add_oh_shift_1[14];
  assign _zz_add_oh_shift_12 = _zz_add_oh_shift_1[15];
  assign _zz_add_oh_shift_13 = _zz_add_oh_shift_1[17];
  assign _zz_add_oh_shift_14 = _zz_add_oh_shift_1[18];
  assign _zz_add_oh_shift_15 = _zz_add_oh_shift_1[19];
  assign _zz_add_oh_shift_16 = _zz_add_oh_shift_1[20];
  assign _zz_add_oh_shift_17 = _zz_add_oh_shift_1[21];
  assign _zz_add_oh_shift_18 = _zz_add_oh_shift_1[22];
  assign _zz_add_oh_shift_19 = _zz_add_oh_shift_1[23];
  assign _zz_add_oh_shift_20 = _zz_add_oh_shift_1[24];
  assign _zz_add_oh_shift_21 = _zz_add_oh_shift_1[25];
  assign _zz_add_oh_shift_22 = _zz_add_oh_shift_1[26];
  assign _zz_add_oh_shift_23 = _zz_add_oh_shift_1[27];
  assign _zz_add_oh_shift_24 = _zz_add_oh_shift_1[28];
  assign _zz_add_oh_shift_25 = _zz_add_oh_shift_1[29];
  assign _zz_add_oh_shift_26 = _zz_add_oh_shift_1[30];
  assign _zz_add_oh_shift_27 = _zz_add_oh_shift_1[31];
  assign _zz_add_oh_shift_28 = _zz_add_oh_shift_1[33];
  assign _zz_add_oh_shift_29 = _zz_add_oh_shift_1[34];
  assign _zz_add_oh_shift_30 = _zz_add_oh_shift_1[35];
  assign _zz_add_oh_shift_31 = _zz_add_oh_shift_1[36];
  assign _zz_add_oh_shift_32 = _zz_add_oh_shift_1[37];
  assign _zz_add_oh_shift_33 = _zz_add_oh_shift_1[38];
  assign _zz_add_oh_shift_34 = _zz_add_oh_shift_1[39];
  assign _zz_add_oh_shift_35 = _zz_add_oh_shift_1[40];
  assign _zz_add_oh_shift_36 = _zz_add_oh_shift_1[41];
  assign _zz_add_oh_shift_37 = _zz_add_oh_shift_1[42];
  assign _zz_add_oh_shift_38 = _zz_add_oh_shift_1[43];
  assign _zz_add_oh_shift_39 = _zz_add_oh_shift_1[44];
  assign _zz_add_oh_shift_40 = _zz_add_oh_shift_1[45];
  assign _zz_add_oh_shift_41 = _zz_add_oh_shift_1[46];
  assign _zz_add_oh_shift_42 = _zz_add_oh_shift_1[47];
  assign _zz_add_oh_shift_43 = _zz_add_oh_shift_1[48];
  assign _zz_add_oh_shift_44 = _zz_add_oh_shift_1[49];
  assign _zz_add_oh_shift_45 = _zz_add_oh_shift_1[50];
  assign _zz_add_oh_shift_46 = _zz_add_oh_shift_1[51];
  assign _zz_add_oh_shift_47 = _zz_add_oh_shift_1[52];
  assign _zz_add_oh_shift_48 = _zz_add_oh_shift_1[53];
  assign _zz_add_oh_shift_49 = _zz_add_oh_shift_1[54];
  assign _zz_add_oh_shift_50 = _zz_add_oh_shift_1[55];
  assign _zz_add_oh_shift_51 = ((((((((((((((((_zz__zz_add_oh_shift_51 || _zz_add_oh_shift_21) || _zz_add_oh_shift_23) || _zz_add_oh_shift_25) || _zz_add_oh_shift_27) || _zz_add_oh_shift_28) || _zz_add_oh_shift_30) || _zz_add_oh_shift_32) || _zz_add_oh_shift_34) || _zz_add_oh_shift_36) || _zz_add_oh_shift_38) || _zz_add_oh_shift_40) || _zz_add_oh_shift_42) || _zz_add_oh_shift_44) || _zz_add_oh_shift_46) || _zz_add_oh_shift_48) || _zz_add_oh_shift_50);
  assign _zz_add_oh_shift_52 = ((((((((((((((((_zz__zz_add_oh_shift_52 || _zz_add_oh_shift_22) || _zz_add_oh_shift_23) || _zz_add_oh_shift_26) || _zz_add_oh_shift_27) || _zz_add_oh_shift_29) || _zz_add_oh_shift_30) || _zz_add_oh_shift_33) || _zz_add_oh_shift_34) || _zz_add_oh_shift_37) || _zz_add_oh_shift_38) || _zz_add_oh_shift_41) || _zz_add_oh_shift_42) || _zz_add_oh_shift_45) || _zz_add_oh_shift_46) || _zz_add_oh_shift_49) || _zz_add_oh_shift_50);
  assign _zz_add_oh_shift_53 = ((((((((((((((((_zz__zz_add_oh_shift_53 || _zz_add_oh_shift_24) || _zz_add_oh_shift_25) || _zz_add_oh_shift_26) || _zz_add_oh_shift_27) || _zz_add_oh_shift_31) || _zz_add_oh_shift_32) || _zz_add_oh_shift_33) || _zz_add_oh_shift_34) || _zz_add_oh_shift_39) || _zz_add_oh_shift_40) || _zz_add_oh_shift_41) || _zz_add_oh_shift_42) || _zz_add_oh_shift_47) || _zz_add_oh_shift_48) || _zz_add_oh_shift_49) || _zz_add_oh_shift_50);
  assign _zz_add_oh_shift_54 = (((((((((((((((((_zz__zz_add_oh_shift_54 || _zz_add_oh_shift_12) || _zz_add_oh_shift_20) || _zz_add_oh_shift_21) || _zz_add_oh_shift_22) || _zz_add_oh_shift_23) || _zz_add_oh_shift_24) || _zz_add_oh_shift_25) || _zz_add_oh_shift_26) || _zz_add_oh_shift_27) || _zz_add_oh_shift_35) || _zz_add_oh_shift_36) || _zz_add_oh_shift_37) || _zz_add_oh_shift_38) || _zz_add_oh_shift_39) || _zz_add_oh_shift_40) || _zz_add_oh_shift_41) || _zz_add_oh_shift_42);
  assign _zz_add_oh_shift_55 = (((((((((((((((((_zz__zz_add_oh_shift_55 || _zz_add_oh_shift_19) || _zz_add_oh_shift_20) || _zz_add_oh_shift_21) || _zz_add_oh_shift_22) || _zz_add_oh_shift_23) || _zz_add_oh_shift_24) || _zz_add_oh_shift_25) || _zz_add_oh_shift_26) || _zz_add_oh_shift_27) || _zz_add_oh_shift_43) || _zz_add_oh_shift_44) || _zz_add_oh_shift_45) || _zz_add_oh_shift_46) || _zz_add_oh_shift_47) || _zz_add_oh_shift_48) || _zz_add_oh_shift_49) || _zz_add_oh_shift_50);
  assign _zz_add_oh_shift_56 = ((((((((((((((((_zz__zz_add_oh_shift_56 || _zz_add_oh_shift_35) || _zz_add_oh_shift_36) || _zz_add_oh_shift_37) || _zz_add_oh_shift_38) || _zz_add_oh_shift_39) || _zz_add_oh_shift_40) || _zz_add_oh_shift_41) || _zz_add_oh_shift_42) || _zz_add_oh_shift_43) || _zz_add_oh_shift_44) || _zz_add_oh_shift_45) || _zz_add_oh_shift_46) || _zz_add_oh_shift_47) || _zz_add_oh_shift_48) || _zz_add_oh_shift_49) || _zz_add_oh_shift_50);
  assign add_oh_shift = {_zz_add_oh_shift_56,{_zz_add_oh_shift_55,{_zz_add_oh_shift_54,{_zz_add_oh_shift_53,{_zz_add_oh_shift_52,_zz_add_oh_shift_51}}}}};
  assign add_oh_output_payload_shift = add_oh_shift;
  always @(*) begin
    add_oh_output_ready = add_norm_input_ready;
    if(when_Stream_l375_18) begin
      add_oh_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_18 = (! add_norm_input_valid);
  assign add_norm_input_valid = add_oh_output_rValid;
  assign add_norm_input_payload_source = add_oh_output_rData_source;
  assign add_norm_input_payload_rs1_mantissa = add_oh_output_rData_rs1_mantissa;
  assign add_norm_input_payload_rs1_exponent = add_oh_output_rData_rs1_exponent;
  assign add_norm_input_payload_rs1_sign = add_oh_output_rData_rs1_sign;
  assign add_norm_input_payload_rs1_special = add_oh_output_rData_rs1_special;
  assign add_norm_input_payload_rs2_mantissa = add_oh_output_rData_rs2_mantissa;
  assign add_norm_input_payload_rs2_exponent = add_oh_output_rData_rs2_exponent;
  assign add_norm_input_payload_rs2_sign = add_oh_output_rData_rs2_sign;
  assign add_norm_input_payload_rs2_special = add_oh_output_rData_rs2_special;
  assign add_norm_input_payload_rd = add_oh_output_rData_rd;
  assign add_norm_input_payload_roundMode = add_oh_output_rData_roundMode;
  assign add_norm_input_payload_format = add_oh_output_rData_format;
  assign add_norm_input_payload_needCommit = add_oh_output_rData_needCommit;
  assign add_norm_input_payload_xSign = add_oh_output_rData_xSign;
  assign add_norm_input_payload_ySign = add_oh_output_rData_ySign;
  assign add_norm_input_payload_xMantissa = add_oh_output_rData_xMantissa;
  assign add_norm_input_payload_yMantissa = add_oh_output_rData_yMantissa;
  assign add_norm_input_payload_xyExponent = add_oh_output_rData_xyExponent;
  assign add_norm_input_payload_xySign = add_oh_output_rData_xySign;
  assign add_norm_input_payload_roundingScrap = add_oh_output_rData_roundingScrap;
  assign add_norm_input_payload_xyMantissa = add_oh_output_rData_xyMantissa;
  assign add_norm_input_payload_shift = add_oh_output_rData_shift;
  assign add_norm_output_valid = add_norm_input_valid;
  assign add_norm_input_ready = add_norm_output_ready;
  assign add_norm_output_payload_source = add_norm_input_payload_source;
  assign add_norm_output_payload_rs1_mantissa = add_norm_input_payload_rs1_mantissa;
  assign add_norm_output_payload_rs1_exponent = add_norm_input_payload_rs1_exponent;
  assign add_norm_output_payload_rs1_sign = add_norm_input_payload_rs1_sign;
  assign add_norm_output_payload_rs1_special = add_norm_input_payload_rs1_special;
  assign add_norm_output_payload_rs2_mantissa = add_norm_input_payload_rs2_mantissa;
  assign add_norm_output_payload_rs2_exponent = add_norm_input_payload_rs2_exponent;
  assign add_norm_output_payload_rs2_sign = add_norm_input_payload_rs2_sign;
  assign add_norm_output_payload_rs2_special = add_norm_input_payload_rs2_special;
  assign add_norm_output_payload_rd = add_norm_input_payload_rd;
  assign add_norm_output_payload_roundMode = add_norm_input_payload_roundMode;
  assign add_norm_output_payload_format = add_norm_input_payload_format;
  assign add_norm_output_payload_needCommit = add_norm_input_payload_needCommit;
  assign add_norm_output_payload_xySign = add_norm_input_payload_xySign;
  assign add_norm_output_payload_roundingScrap = add_norm_input_payload_roundingScrap;
  assign add_norm_output_payload_mantissa = (add_norm_input_payload_xyMantissa <<< add_norm_input_payload_shift);
  assign add_norm_output_payload_exponent = (_zz_add_norm_output_payload_exponent + 13'h0001);
  assign add_norm_output_payload_forceInfinity = ((add_norm_input_payload_rs1_special && (add_norm_input_payload_rs1_exponent[1 : 0] == 2'b01)) || (add_norm_input_payload_rs2_special && (add_norm_input_payload_rs2_exponent[1 : 0] == 2'b01)));
  assign add_norm_output_payload_forceZero = ((add_norm_input_payload_xyMantissa == 56'h0) || ((add_norm_input_payload_rs1_special && (add_norm_input_payload_rs1_exponent[1 : 0] == 2'b00)) && (add_norm_input_payload_rs2_special && (add_norm_input_payload_rs2_exponent[1 : 0] == 2'b00))));
  assign add_norm_output_payload_infinityNan = (((add_norm_input_payload_rs1_special && (add_norm_input_payload_rs1_exponent[1 : 0] == 2'b01)) && (add_norm_input_payload_rs2_special && (add_norm_input_payload_rs2_exponent[1 : 0] == 2'b01))) && (add_norm_input_payload_rs1_sign ^ add_norm_input_payload_rs2_sign));
  assign add_norm_output_payload_forceNan = (((add_norm_input_payload_rs1_special && (add_norm_input_payload_rs1_exponent[1 : 0] == 2'b10)) || (add_norm_input_payload_rs2_special && (add_norm_input_payload_rs2_exponent[1 : 0] == 2'b10))) || add_norm_output_payload_infinityNan);
  assign add_norm_output_payload_xyMantissaZero = (add_norm_input_payload_xyMantissa == 56'h0);
  assign add_result_input_valid = add_norm_output_valid;
  assign add_norm_output_ready = add_result_input_ready;
  assign add_result_input_payload_source = add_norm_output_payload_source;
  assign add_result_input_payload_rs1_mantissa = add_norm_output_payload_rs1_mantissa;
  assign add_result_input_payload_rs1_exponent = add_norm_output_payload_rs1_exponent;
  assign add_result_input_payload_rs1_sign = add_norm_output_payload_rs1_sign;
  assign add_result_input_payload_rs1_special = add_norm_output_payload_rs1_special;
  assign add_result_input_payload_rs2_mantissa = add_norm_output_payload_rs2_mantissa;
  assign add_result_input_payload_rs2_exponent = add_norm_output_payload_rs2_exponent;
  assign add_result_input_payload_rs2_sign = add_norm_output_payload_rs2_sign;
  assign add_result_input_payload_rs2_special = add_norm_output_payload_rs2_special;
  assign add_result_input_payload_rd = add_norm_output_payload_rd;
  assign add_result_input_payload_roundMode = add_norm_output_payload_roundMode;
  assign add_result_input_payload_format = add_norm_output_payload_format;
  assign add_result_input_payload_needCommit = add_norm_output_payload_needCommit;
  assign add_result_input_payload_mantissa = add_norm_output_payload_mantissa;
  assign add_result_input_payload_exponent = add_norm_output_payload_exponent;
  assign add_result_input_payload_infinityNan = add_norm_output_payload_infinityNan;
  assign add_result_input_payload_forceNan = add_norm_output_payload_forceNan;
  assign add_result_input_payload_forceZero = add_norm_output_payload_forceZero;
  assign add_result_input_payload_forceInfinity = add_norm_output_payload_forceInfinity;
  assign add_result_input_payload_xySign = add_norm_output_payload_xySign;
  assign add_result_input_payload_roundingScrap = add_norm_output_payload_roundingScrap;
  assign add_result_input_payload_xyMantissaZero = add_norm_output_payload_xyMantissaZero;
  assign add_result_output_valid = add_result_input_valid;
  assign add_result_input_ready = add_result_output_ready;
  assign add_result_output_payload_source = add_result_input_payload_source;
  assign add_result_output_payload_rd = add_result_input_payload_rd;
  always @(*) begin
    add_result_output_payload_value_sign = add_result_input_payload_xySign;
    if(!add_result_input_payload_forceNan) begin
      if(!add_result_input_payload_forceInfinity) begin
        if(add_result_input_payload_forceZero) begin
          if(when_FpuCore_l1513) begin
            add_result_output_payload_value_sign = (add_result_input_payload_rs1_sign && add_result_input_payload_rs2_sign);
          end
          if(when_FpuCore_l1516) begin
            add_result_output_payload_value_sign = 1'b1;
          end
        end
      end
    end
  end

  always @(*) begin
    add_result_output_payload_value_mantissa = _zz_add_result_output_payload_value_mantissa[52:0];
    if(add_result_input_payload_forceNan) begin
      add_result_output_payload_value_mantissa[52] = 1'b1;
    end
  end

  always @(*) begin
    add_result_output_payload_value_exponent = add_result_input_payload_exponent[11:0];
    if(add_result_input_payload_forceNan) begin
      add_result_output_payload_value_exponent[1 : 0] = 2'b10;
      add_result_output_payload_value_exponent[2] = 1'b1;
    end else begin
      if(add_result_input_payload_forceInfinity) begin
        add_result_output_payload_value_exponent[1 : 0] = 2'b01;
      end else begin
        if(add_result_input_payload_forceZero) begin
          add_result_output_payload_value_exponent[1 : 0] = 2'b00;
        end
      end
    end
  end

  always @(*) begin
    add_result_output_payload_value_special = 1'b0;
    if(add_result_input_payload_forceNan) begin
      add_result_output_payload_value_special = 1'b1;
    end else begin
      if(add_result_input_payload_forceInfinity) begin
        add_result_output_payload_value_special = 1'b1;
      end else begin
        if(add_result_input_payload_forceZero) begin
          add_result_output_payload_value_special = 1'b1;
        end
      end
    end
  end

  assign add_result_output_payload_roundMode = add_result_input_payload_roundMode;
  assign add_result_output_payload_format = add_result_input_payload_format;
  assign add_result_output_payload_scrap = ((add_result_input_payload_mantissa[1] || add_result_input_payload_mantissa[0]) || add_result_input_payload_roundingScrap);
  assign add_result_output_payload_NV = ((add_result_input_payload_infinityNan || ((add_result_input_payload_rs1_special && (add_result_input_payload_rs1_exponent[1 : 0] == 2'b10)) && (! add_result_input_payload_rs1_mantissa[53]))) || ((add_result_input_payload_rs2_special && (add_result_input_payload_rs2_exponent[1 : 0] == 2'b10)) && (! add_result_input_payload_rs2_mantissa[53])));
  assign add_result_output_payload_DZ = 1'b0;
  assign when_FpuCore_l1513 = (add_result_input_payload_xyMantissaZero || ((add_result_input_payload_rs1_special && (add_result_input_payload_rs1_exponent[1 : 0] == 2'b00)) && (add_result_input_payload_rs2_special && (add_result_input_payload_rs2_exponent[1 : 0] == 2'b00))));
  assign when_FpuCore_l1516 = ((add_result_input_payload_rs1_sign || add_result_input_payload_rs2_sign) && (add_result_input_payload_roundMode == FpuRoundMode_RDN));
  always @(*) begin
    load_s1_output_ready = load_s1_output_m2sPipe_ready;
    if(when_Stream_l375_19) begin
      load_s1_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_19 = (! load_s1_output_m2sPipe_valid);
  assign load_s1_output_m2sPipe_valid = load_s1_output_rValid;
  assign load_s1_output_m2sPipe_payload_source = load_s1_output_rData_source;
  assign load_s1_output_m2sPipe_payload_rd = load_s1_output_rData_rd;
  assign load_s1_output_m2sPipe_payload_value_mantissa = load_s1_output_rData_value_mantissa;
  assign load_s1_output_m2sPipe_payload_value_exponent = load_s1_output_rData_value_exponent;
  assign load_s1_output_m2sPipe_payload_value_sign = load_s1_output_rData_value_sign;
  assign load_s1_output_m2sPipe_payload_value_special = load_s1_output_rData_value_special;
  assign load_s1_output_m2sPipe_payload_scrap = load_s1_output_rData_scrap;
  assign load_s1_output_m2sPipe_payload_roundMode = load_s1_output_rData_roundMode;
  assign load_s1_output_m2sPipe_payload_format = load_s1_output_rData_format;
  assign load_s1_output_m2sPipe_payload_NV = load_s1_output_rData_NV;
  assign load_s1_output_m2sPipe_payload_DZ = load_s1_output_rData_DZ;
  always @(*) begin
    shortPip_output_ready = shortPip_output_m2sPipe_ready;
    if(when_Stream_l375_20) begin
      shortPip_output_ready = 1'b1;
    end
  end

  assign when_Stream_l375_20 = (! shortPip_output_m2sPipe_valid);
  assign shortPip_output_m2sPipe_valid = shortPip_output_rValid;
  assign shortPip_output_m2sPipe_payload_source = shortPip_output_rData_source;
  assign shortPip_output_m2sPipe_payload_rd = shortPip_output_rData_rd;
  assign shortPip_output_m2sPipe_payload_value_mantissa = shortPip_output_rData_value_mantissa;
  assign shortPip_output_m2sPipe_payload_value_exponent = shortPip_output_rData_value_exponent;
  assign shortPip_output_m2sPipe_payload_value_sign = shortPip_output_rData_value_sign;
  assign shortPip_output_m2sPipe_payload_value_special = shortPip_output_rData_value_special;
  assign shortPip_output_m2sPipe_payload_scrap = shortPip_output_rData_scrap;
  assign shortPip_output_m2sPipe_payload_roundMode = shortPip_output_rData_roundMode;
  assign shortPip_output_m2sPipe_payload_format = shortPip_output_rData_format;
  assign shortPip_output_m2sPipe_payload_NV = shortPip_output_rData_NV;
  assign shortPip_output_m2sPipe_payload_DZ = shortPip_output_rData_DZ;
  assign load_s1_output_m2sPipe_ready = streamArbiter_10_io_inputs_0_ready;
  assign sqrt_output_ready = streamArbiter_10_io_inputs_1_ready;
  assign div_output_ready = streamArbiter_10_io_inputs_2_ready;
  assign add_result_output_ready = streamArbiter_10_io_inputs_3_ready;
  assign mul_result_output_ready = streamArbiter_10_io_inputs_4_ready;
  assign shortPip_output_m2sPipe_ready = streamArbiter_10_io_inputs_5_ready;
  assign streamArbiter_10_io_output_combStage_valid = streamArbiter_10_io_output_valid;
  assign streamArbiter_10_io_output_combStage_payload_source = streamArbiter_10_io_output_payload_source;
  assign streamArbiter_10_io_output_combStage_payload_rd = streamArbiter_10_io_output_payload_rd;
  assign streamArbiter_10_io_output_combStage_payload_value_mantissa = streamArbiter_10_io_output_payload_value_mantissa;
  assign streamArbiter_10_io_output_combStage_payload_value_exponent = streamArbiter_10_io_output_payload_value_exponent;
  assign streamArbiter_10_io_output_combStage_payload_value_sign = streamArbiter_10_io_output_payload_value_sign;
  assign streamArbiter_10_io_output_combStage_payload_value_special = streamArbiter_10_io_output_payload_value_special;
  assign streamArbiter_10_io_output_combStage_payload_scrap = streamArbiter_10_io_output_payload_scrap;
  assign streamArbiter_10_io_output_combStage_payload_roundMode = streamArbiter_10_io_output_payload_roundMode;
  assign streamArbiter_10_io_output_combStage_payload_format = streamArbiter_10_io_output_payload_format;
  assign streamArbiter_10_io_output_combStage_payload_NV = streamArbiter_10_io_output_payload_NV;
  assign streamArbiter_10_io_output_combStage_payload_DZ = streamArbiter_10_io_output_payload_DZ;
  assign streamArbiter_10_io_output_combStage_ready = 1'b1;
  assign merge_arbitrated_valid = streamArbiter_10_io_output_combStage_valid;
  assign merge_arbitrated_payload_source = streamArbiter_10_io_output_combStage_payload_source;
  assign merge_arbitrated_payload_rd = streamArbiter_10_io_output_combStage_payload_rd;
  assign merge_arbitrated_payload_value_mantissa = streamArbiter_10_io_output_combStage_payload_value_mantissa;
  assign merge_arbitrated_payload_value_exponent = streamArbiter_10_io_output_combStage_payload_value_exponent;
  assign merge_arbitrated_payload_value_sign = streamArbiter_10_io_output_combStage_payload_value_sign;
  assign merge_arbitrated_payload_value_special = streamArbiter_10_io_output_combStage_payload_value_special;
  assign merge_arbitrated_payload_scrap = streamArbiter_10_io_output_combStage_payload_scrap;
  assign merge_arbitrated_payload_roundMode = streamArbiter_10_io_output_combStage_payload_roundMode;
  assign merge_arbitrated_payload_format = streamArbiter_10_io_output_combStage_payload_format;
  assign merge_arbitrated_payload_NV = streamArbiter_10_io_output_combStage_payload_NV;
  assign merge_arbitrated_payload_DZ = streamArbiter_10_io_output_combStage_payload_DZ;
  assign roundFront_output_valid = roundFront_input_valid;
  assign roundFront_output_payload_source = roundFront_input_payload_source;
  assign roundFront_output_payload_rd = roundFront_input_payload_rd;
  assign roundFront_output_payload_value_mantissa = roundFront_input_payload_value_mantissa;
  assign roundFront_output_payload_value_exponent = roundFront_input_payload_value_exponent;
  assign roundFront_output_payload_value_sign = roundFront_input_payload_value_sign;
  assign roundFront_output_payload_value_special = roundFront_input_payload_value_special;
  assign roundFront_output_payload_scrap = roundFront_input_payload_scrap;
  assign roundFront_output_payload_roundMode = roundFront_input_payload_roundMode;
  assign roundFront_output_payload_format = roundFront_input_payload_format;
  assign roundFront_output_payload_NV = roundFront_input_payload_NV;
  assign roundFront_output_payload_DZ = roundFront_input_payload_DZ;
  assign roundFront_manAggregate = {roundFront_input_payload_value_mantissa,roundFront_input_payload_scrap};
  assign roundFront_expBase = ((roundFront_input_payload_format == FpuFormat_DOUBLE) ? 11'h401 : 11'h781);
  assign roundFront_expDif = (_zz_roundFront_expDif - {1'b0,roundFront_input_payload_value_exponent});
  assign roundFront_expSubnormal = ((! roundFront_input_payload_value_special) && (! roundFront_expDif[12]));
  assign roundFront_discardCount = (roundFront_expSubnormal ? roundFront_expDif : 13'h0);
  assign when_FpuCore_l1551 = (roundFront_input_payload_format == FpuFormat_FLOAT);
  assign roundFront_discardCountTrunk = roundFront_discardCount_1[5:0];
  always @(*) begin
    roundFront_exactMask = {(6'h34 < roundFront_discardCountTrunk),{(6'h33 < roundFront_discardCountTrunk),{(6'h32 < roundFront_discardCountTrunk),{(6'h31 < roundFront_discardCountTrunk),{(_zz_roundFront_exactMask < roundFront_discardCountTrunk),{_zz_roundFront_exactMask_1,{_zz_roundFront_exactMask_2,_zz_roundFront_exactMask_3}}}}}}};
    if(when_FpuCore_l1559) begin
      roundFront_exactMask = 54'h3fffffffffffff;
    end
  end

  always @(*) begin
    roundFront_roundAdjusted = {_zz_roundFront_roundAdjusted[roundFront_discardCountTrunk],((roundFront_manAggregate & roundFront_exactMask) != 54'h0)};
    if(when_FpuCore_l1559) begin
      roundFront_roundAdjusted[1] = 1'b0;
    end
  end

  always @(*) begin
    roundFront_rneBit = _zz_roundFront_rneBit[roundFront_discardCountTrunk];
    if(when_FpuCore_l1559) begin
      roundFront_rneBit = 1'b0;
    end
  end

  assign when_FpuCore_l1559 = (13'h0036 <= roundFront_discardCount_1);
  always @(*) begin
    case(roundFront_input_payload_roundMode)
      FpuRoundMode_RNE : begin
        _zz_roundFront_mantissaIncrement = (roundFront_roundAdjusted[1] && (roundFront_roundAdjusted[0] || roundFront_rneBit));
      end
      FpuRoundMode_RTZ : begin
        _zz_roundFront_mantissaIncrement = 1'b0;
      end
      FpuRoundMode_RDN : begin
        _zz_roundFront_mantissaIncrement = ((roundFront_roundAdjusted != 2'b00) && roundFront_input_payload_value_sign);
      end
      FpuRoundMode_RUP : begin
        _zz_roundFront_mantissaIncrement = ((roundFront_roundAdjusted != 2'b00) && (! roundFront_input_payload_value_sign));
      end
      default : begin
        _zz_roundFront_mantissaIncrement = roundFront_roundAdjusted[1];
      end
    endcase
  end

  assign roundFront_mantissaIncrement = ((! roundFront_input_payload_value_special) && _zz_roundFront_mantissaIncrement);
  assign roundFront_output_payload_mantissaIncrement = roundFront_mantissaIncrement;
  assign roundFront_output_payload_roundAdjusted = roundFront_roundAdjusted;
  assign roundFront_output_payload_exactMask = roundFront_exactMask;
  assign roundBack_output_valid = roundBack_input_valid;
  assign roundBack_adderMantissa = (roundBack_input_payload_value_mantissa[52 : 1] & (roundBack_input_payload_mantissaIncrement ? (~ _zz_roundBack_adderMantissa) : 52'hfffffffffffff));
  assign roundBack_adderRightOp = _zz_roundBack_adderRightOp[51:0];
  assign _zz_roundBack_adder = {roundBack_input_payload_value_exponent,roundBack_adderMantissa};
  assign _zz_roundBack_adder_1 = roundBack_input_payload_mantissaIncrement;
  assign roundBack_adder = (_zz_roundBack_adder_2 + _zz_roundBack_adder_4);
  assign roundBack_masked = (roundBack_adder & (~ _zz_roundBack_masked));
  assign roundBack_math_special = roundBack_input_payload_value_special;
  assign roundBack_math_sign = roundBack_input_payload_value_sign;
  assign roundBack_math_exponent = roundBack_masked[63 : 52];
  assign roundBack_math_mantissa = roundBack_masked[51 : 0];
  always @(*) begin
    roundBack_patched_mantissa = roundBack_math_mantissa;
    if(when_FpuCore_l1619) begin
      if(when_FpuCore_l1629) begin
        roundBack_patched_mantissa = 52'hfffffffffffff;
      end
    end
    if(when_FpuCore_l1638) begin
      if(when_FpuCore_l1648) begin
        roundBack_patched_mantissa = 52'h0;
      end
    end
  end

  always @(*) begin
    roundBack_patched_exponent = roundBack_math_exponent;
    if(when_FpuCore_l1619) begin
      if(when_FpuCore_l1629) begin
        roundBack_patched_exponent = roundBack_ofThreshold;
      end else begin
        roundBack_patched_exponent[1 : 0] = 2'b01;
      end
    end
    if(when_FpuCore_l1638) begin
      if(when_FpuCore_l1648) begin
        roundBack_patched_exponent = {1'd0, roundBack_ufThreshold};
      end else begin
        roundBack_patched_exponent[1 : 0] = 2'b00;
      end
    end
  end

  assign roundBack_patched_sign = roundBack_math_sign;
  always @(*) begin
    roundBack_patched_special = roundBack_math_special;
    if(when_FpuCore_l1619) begin
      if(!when_FpuCore_l1629) begin
        roundBack_patched_special = 1'b1;
      end
    end
    if(when_FpuCore_l1638) begin
      if(!when_FpuCore_l1648) begin
        roundBack_patched_special = 1'b1;
      end
    end
  end

  always @(*) begin
    roundBack_nx = 1'b0;
    if(when_FpuCore_l1619) begin
      roundBack_nx = 1'b1;
    end
    if(when_FpuCore_l1638) begin
      roundBack_nx = 1'b1;
    end
    if(when_FpuCore_l1657) begin
      roundBack_nx = 1'b1;
    end
  end

  always @(*) begin
    roundBack_of = 1'b0;
    if(when_FpuCore_l1619) begin
      roundBack_of = 1'b1;
    end
  end

  always @(*) begin
    roundBack_uf = 1'b0;
    if(when_FpuCore_l1616) begin
      roundBack_uf = 1'b1;
    end
    if(when_FpuCore_l1638) begin
      roundBack_uf = 1'b1;
    end
  end

  assign roundBack_ufSubnormalThreshold = ((roundBack_input_payload_format == FpuFormat_DOUBLE) ? 11'h400 : 11'h780);
  assign roundBack_ufThreshold = ((roundBack_input_payload_format == FpuFormat_DOUBLE) ? 11'h3cd : 11'h76a);
  assign roundBack_ofThreshold = ((roundBack_input_payload_format == FpuFormat_DOUBLE) ? 12'hbfe : 12'h87e);
  always @(*) begin
    case(roundBack_input_payload_roundMode)
      FpuRoundMode_RNE : begin
        roundBack_threshold = 3'b110;
      end
      FpuRoundMode_RTZ : begin
        roundBack_threshold = 3'b110;
      end
      FpuRoundMode_RDN : begin
        roundBack_threshold = (roundBack_input_payload_value_sign ? 3'b101 : 3'b111);
      end
      FpuRoundMode_RUP : begin
        roundBack_threshold = (roundBack_input_payload_value_sign ? 3'b111 : 3'b101);
      end
      default : begin
        roundBack_threshold = 3'b110;
      end
    endcase
  end

  always @(*) begin
    roundBack_borringRound = {roundBack_input_payload_value_mantissa[1 : 0],roundBack_input_payload_scrap};
    if(when_FpuCore_l1613) begin
      roundBack_borringRound = {roundBack_input_payload_value_mantissa[30 : 29],(|roundBack_input_payload_value_mantissa[28 : 0])};
    end
  end

  assign when_FpuCore_l1613 = (roundBack_input_payload_format == FpuFormat_FLOAT);
  assign roundBack_borringCase = ((roundBack_input_payload_value_exponent == _zz_roundBack_borringCase) && (roundBack_borringRound < roundBack_threshold));
  assign when_FpuCore_l1616 = (((! roundBack_math_special) && ((roundBack_math_exponent <= _zz_when_FpuCore_l1616) || roundBack_borringCase)) && (roundBack_input_payload_roundAdjusted != 2'b00));
  assign when_FpuCore_l1619 = ((! roundBack_math_special) && (roundBack_ofThreshold < roundBack_math_exponent));
  always @(*) begin
    case(roundBack_input_payload_roundMode)
      FpuRoundMode_RNE : begin
        when_FpuCore_l1629 = 1'b0;
      end
      FpuRoundMode_RTZ : begin
        when_FpuCore_l1629 = 1'b1;
      end
      FpuRoundMode_RDN : begin
        when_FpuCore_l1629 = (! roundBack_math_sign);
      end
      FpuRoundMode_RUP : begin
        when_FpuCore_l1629 = roundBack_math_sign;
      end
      default : begin
        when_FpuCore_l1629 = 1'b0;
      end
    endcase
  end

  assign when_FpuCore_l1638 = ((! roundBack_math_special) && (roundBack_math_exponent < _zz_when_FpuCore_l1638));
  always @(*) begin
    case(roundBack_input_payload_roundMode)
      FpuRoundMode_RNE : begin
        when_FpuCore_l1648 = 1'b0;
      end
      FpuRoundMode_RTZ : begin
        when_FpuCore_l1648 = 1'b0;
      end
      FpuRoundMode_RDN : begin
        when_FpuCore_l1648 = roundBack_math_sign;
      end
      FpuRoundMode_RUP : begin
        when_FpuCore_l1648 = (! roundBack_math_sign);
      end
      default : begin
        when_FpuCore_l1648 = 1'b0;
      end
    endcase
  end

  assign when_FpuCore_l1657 = ((! roundBack_input_payload_value_special) && (roundBack_input_payload_roundAdjusted != 2'b00));
  assign roundBack_writes_0 = rf_scoreboards_0_writes_spinal_port1[0];
  assign roundBack_writes_1 = rf_scoreboards_1_writes_spinal_port1[0];
  assign roundBack_write = _zz_roundBack_write;
  assign roundBack_output_payload_NX = (roundBack_nx && roundBack_write);
  assign roundBack_output_payload_OF = (roundBack_of && roundBack_write);
  assign roundBack_output_payload_UF = (roundBack_uf && roundBack_write);
  assign roundBack_output_payload_NV = (roundBack_input_payload_NV && roundBack_write);
  assign roundBack_output_payload_DZ = (roundBack_input_payload_DZ && roundBack_write);
  assign roundBack_output_payload_source = roundBack_input_payload_source;
  assign roundBack_output_payload_rd = roundBack_input_payload_rd;
  assign roundBack_output_payload_write = roundBack_write;
  assign roundBack_output_payload_format = roundBack_input_payload_format;
  assign roundBack_output_payload_value_mantissa = roundBack_patched_mantissa;
  assign roundBack_output_payload_value_exponent = roundBack_patched_exponent;
  assign roundBack_output_payload_value_sign = roundBack_patched_sign;
  assign roundBack_output_payload_value_special = roundBack_patched_special;
  assign io_port_0_completion_valid = (writeback_input_valid && (writeback_input_payload_source == 1'b0));
  assign io_port_0_completion_payload_flags_NX = writeback_input_payload_NX;
  assign io_port_0_completion_payload_flags_OF = writeback_input_payload_OF;
  assign io_port_0_completion_payload_flags_UF = writeback_input_payload_UF;
  assign io_port_0_completion_payload_flags_NV = writeback_input_payload_NV;
  assign io_port_0_completion_payload_flags_DZ = writeback_input_payload_DZ;
  assign io_port_0_completion_payload_written = writeback_input_payload_write;
  assign io_port_1_completion_valid = (writeback_input_valid && (writeback_input_payload_source == 1'b1));
  assign io_port_1_completion_payload_flags_NX = writeback_input_payload_NX;
  assign io_port_1_completion_payload_flags_OF = writeback_input_payload_OF;
  assign io_port_1_completion_payload_flags_UF = writeback_input_payload_UF;
  assign io_port_1_completion_payload_flags_NV = writeback_input_payload_NV;
  assign io_port_1_completion_payload_flags_DZ = writeback_input_payload_DZ;
  assign io_port_1_completion_payload_written = writeback_input_payload_write;
  assign when_FpuCore_l1689 = (writeback_input_payload_source == 1'b0);
  assign when_FpuCore_l1689_1 = (writeback_input_payload_source == 1'b1);
  assign writeback_port_valid = (writeback_input_valid && writeback_input_payload_write);
  assign writeback_port_payload_address = {writeback_input_payload_source,writeback_input_payload_rd};
  always @(*) begin
    writeback_port_payload_data_value_mantissa = writeback_input_payload_value_mantissa;
    if(writeback_port_payload_data_boxed) begin
      writeback_port_payload_data_value_mantissa[28 : 0] = 29'h0;
    end
  end

  assign writeback_port_payload_data_value_exponent = writeback_input_payload_value_exponent;
  assign writeback_port_payload_data_value_sign = writeback_input_payload_value_sign;
  assign writeback_port_payload_data_value_special = writeback_input_payload_value_special;
  assign writeback_port_payload_data_boxed = (writeback_input_payload_format == FpuFormat_FLOAT);
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      rf_init_counter <= 6'h0;
      streamFork_3_io_outputs_1_rValidN <= 1'b1;
      streamFork_4_io_outputs_1_rValidN <= 1'b1;
      commitLogic_0_pending_counter <= 4'b0000;
      commitLogic_0_add_counter <= 4'b0000;
      commitLogic_0_mul_counter <= 4'b0000;
      commitLogic_0_div_counter <= 4'b0000;
      commitLogic_0_sqrt_counter <= 4'b0000;
      commitLogic_0_short_counter <= 4'b0000;
      commitLogic_1_pending_counter <= 4'b0000;
      commitLogic_1_add_counter <= 4'b0000;
      commitLogic_1_mul_counter <= 4'b0000;
      commitLogic_1_div_counter <= 4'b0000;
      commitLogic_1_sqrt_counter <= 4'b0000;
      commitLogic_1_short_counter <= 4'b0000;
      io_port_0_cmd_rValidN <= 1'b1;
      io_port_1_cmd_rValidN <= 1'b1;
      scheduler_0_output_rValid <= 1'b0;
      scheduler_1_output_rValid <= 1'b0;
      read_s0_rValid <= 1'b0;
      decode_load_rValidN <= 1'b1;
      decode_load_s2mPipe_rValid <= 1'b0;
      decode_load_s2mPipe_m2sPipe_rValid <= 1'b0;
      load_s0_output_rValid <= 1'b0;
      decode_shortPip_rValid <= 1'b0;
      shortPip_rspStreams_0_rValid <= 1'b0;
      shortPip_rspStreams_1_rValid <= 1'b0;
      decode_mul_rValid <= 1'b0;
      mul_preMul_output_rValid <= 1'b0;
      mul_mul_output_rValid <= 1'b0;
      mul_sum1_output_rValid <= 1'b0;
      mul_sum2_output_rValid <= 1'b0;
      mul_result_mulToAdd_rValid <= 1'b0;
      decode_div_rValid <= 1'b0;
      div_cmdSent <= 1'b0;
      decode_sqrt_rValid <= 1'b0;
      sqrt_cmdSent <= 1'b0;
      add_preShifter_output_rValid <= 1'b0;
      add_shifter_output_rValid <= 1'b0;
      add_math_output_rValid <= 1'b0;
      add_oh_output_rValid <= 1'b0;
      load_s1_output_rValid <= 1'b0;
      shortPip_output_rValid <= 1'b0;
      roundFront_input_valid <= 1'b0;
      roundBack_input_valid <= 1'b0;
      writeback_input_valid <= 1'b0;
    end else begin
      if(when_FpuCore_l163) begin
        rf_init_counter <= (rf_init_counter + 6'h01);
      end
      if(streamFork_3_io_outputs_1_valid) begin
        streamFork_3_io_outputs_1_rValidN <= 1'b0;
      end
      if(streamFork_3_io_outputs_1_s2mPipe_ready) begin
        streamFork_3_io_outputs_1_rValidN <= 1'b1;
      end
      if(streamFork_4_io_outputs_1_valid) begin
        streamFork_4_io_outputs_1_rValidN <= 1'b0;
      end
      if(streamFork_4_io_outputs_1_s2mPipe_ready) begin
        streamFork_4_io_outputs_1_rValidN <= 1'b1;
      end
      commitLogic_0_pending_counter <= (_zz_commitLogic_0_pending_counter - _zz_commitLogic_0_pending_counter_3);
      commitLogic_0_add_counter <= (_zz_commitLogic_0_add_counter - _zz_commitLogic_0_add_counter_3);
      commitLogic_0_mul_counter <= (_zz_commitLogic_0_mul_counter - _zz_commitLogic_0_mul_counter_3);
      commitLogic_0_div_counter <= (_zz_commitLogic_0_div_counter - _zz_commitLogic_0_div_counter_3);
      commitLogic_0_sqrt_counter <= (_zz_commitLogic_0_sqrt_counter - _zz_commitLogic_0_sqrt_counter_3);
      commitLogic_0_short_counter <= (_zz_commitLogic_0_short_counter - _zz_commitLogic_0_short_counter_3);
      commitLogic_1_pending_counter <= (_zz_commitLogic_1_pending_counter - _zz_commitLogic_1_pending_counter_3);
      commitLogic_1_add_counter <= (_zz_commitLogic_1_add_counter - _zz_commitLogic_1_add_counter_3);
      commitLogic_1_mul_counter <= (_zz_commitLogic_1_mul_counter - _zz_commitLogic_1_mul_counter_3);
      commitLogic_1_div_counter <= (_zz_commitLogic_1_div_counter - _zz_commitLogic_1_div_counter_3);
      commitLogic_1_sqrt_counter <= (_zz_commitLogic_1_sqrt_counter - _zz_commitLogic_1_sqrt_counter_3);
      commitLogic_1_short_counter <= (_zz_commitLogic_1_short_counter - _zz_commitLogic_1_short_counter_3);
      if(io_port_0_cmd_valid) begin
        io_port_0_cmd_rValidN <= 1'b0;
      end
      if(scheduler_0_input_ready) begin
        io_port_0_cmd_rValidN <= 1'b1;
      end
      if(io_port_1_cmd_valid) begin
        io_port_1_cmd_rValidN <= 1'b0;
      end
      if(scheduler_1_input_ready) begin
        io_port_1_cmd_rValidN <= 1'b1;
      end
      if(scheduler_0_output_ready) begin
        scheduler_0_output_rValid <= scheduler_0_output_valid;
      end
      if(scheduler_1_output_ready) begin
        scheduler_1_output_rValid <= scheduler_1_output_valid;
      end
      if(read_s0_ready) begin
        read_s0_rValid <= read_s0_valid;
      end
      if(decode_load_valid) begin
        decode_load_rValidN <= 1'b0;
      end
      if(decode_load_s2mPipe_ready) begin
        decode_load_rValidN <= 1'b1;
      end
      if(decode_load_s2mPipe_ready) begin
        decode_load_s2mPipe_rValid <= decode_load_s2mPipe_valid;
      end
      if(decode_load_s2mPipe_m2sPipe_ready) begin
        decode_load_s2mPipe_m2sPipe_rValid <= decode_load_s2mPipe_m2sPipe_valid;
      end
      if(load_s0_output_ready) begin
        load_s0_output_rValid <= load_s0_output_valid;
      end
      if(decode_shortPip_ready) begin
        decode_shortPip_rValid <= decode_shortPip_valid;
      end
      if(shortPip_rspStreams_0_ready) begin
        shortPip_rspStreams_0_rValid <= shortPip_rspStreams_0_valid;
      end
      if(shortPip_rspStreams_1_ready) begin
        shortPip_rspStreams_1_rValid <= shortPip_rspStreams_1_valid;
      end
      if(decode_mul_ready) begin
        decode_mul_rValid <= decode_mul_valid;
      end
      if(mul_preMul_output_ready) begin
        mul_preMul_output_rValid <= mul_preMul_output_valid;
      end
      if(mul_mul_output_ready) begin
        mul_mul_output_rValid <= mul_mul_output_valid;
      end
      if(mul_sum1_output_ready) begin
        mul_sum1_output_rValid <= mul_sum1_output_valid;
      end
      if(mul_sum2_output_ready) begin
        mul_sum2_output_rValid <= mul_sum2_output_valid;
      end
      if(mul_result_mulToAdd_ready) begin
        mul_result_mulToAdd_rValid <= mul_result_mulToAdd_valid;
      end
      if(decode_div_valid) begin
        decode_div_rValid <= 1'b1;
      end
      if(div_input_fire) begin
        decode_div_rValid <= 1'b0;
      end
      if(div_divider_io_input_fire) begin
        div_cmdSent <= 1'b1;
      end
      if(when_FpuCore_l1056) begin
        div_cmdSent <= 1'b0;
      end
      if(decode_sqrt_valid) begin
        decode_sqrt_rValid <= 1'b1;
      end
      if(sqrt_input_fire) begin
        decode_sqrt_rValid <= 1'b0;
      end
      if(sqrt_sqrt_io_input_fire) begin
        sqrt_cmdSent <= 1'b1;
      end
      if(when_FpuCore_l1118) begin
        sqrt_cmdSent <= 1'b0;
      end
      if(add_preShifter_output_ready) begin
        add_preShifter_output_rValid <= add_preShifter_output_valid;
      end
      if(add_shifter_output_ready) begin
        add_shifter_output_rValid <= add_shifter_output_valid;
      end
      if(add_math_output_ready) begin
        add_math_output_rValid <= add_math_output_valid;
      end
      if(add_oh_output_ready) begin
        add_oh_output_rValid <= add_oh_output_valid;
      end
      if(load_s1_output_ready) begin
        load_s1_output_rValid <= load_s1_output_valid;
      end
      if(shortPip_output_ready) begin
        shortPip_output_rValid <= shortPip_output_valid;
      end
      roundFront_input_valid <= merge_arbitrated_valid;
      roundBack_input_valid <= roundFront_output_valid;
      writeback_input_valid <= roundBack_output_valid;
      if(writeback_port_valid) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((! ((writeback_port_payload_data_value_exponent == 12'h0) && (! writeback_port_payload_data_value_special)))); // FpuCore.scala:L1718
          `else
            if(!(! ((writeback_port_payload_data_value_exponent == 12'h0) && (! writeback_port_payload_data_value_special)))) begin
              $display("FAILURE Special violation"); // FpuCore.scala:L1718
              $finish;
            end
          `endif
        `endif
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert((! ((writeback_port_payload_data_value_exponent == 12'hfff) && (! writeback_port_payload_data_value_special)))); // FpuCore.scala:L1719
          `else
            if(!(! ((writeback_port_payload_data_value_exponent == 12'hfff) && (! writeback_port_payload_data_value_special)))) begin
              $display("FAILURE Special violation"); // FpuCore.scala:L1719
              $finish;
            end
          `endif
        `endif
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(streamFork_3_io_outputs_1_rValidN) begin
      streamFork_3_io_outputs_1_rData_opcode <= streamFork_3_io_outputs_1_payload_opcode;
      streamFork_3_io_outputs_1_rData_rd <= streamFork_3_io_outputs_1_payload_rd;
      streamFork_3_io_outputs_1_rData_write <= streamFork_3_io_outputs_1_payload_write;
      streamFork_3_io_outputs_1_rData_value <= streamFork_3_io_outputs_1_payload_value;
    end
    if(streamFork_4_io_outputs_1_rValidN) begin
      streamFork_4_io_outputs_1_rData_opcode <= streamFork_4_io_outputs_1_payload_opcode;
      streamFork_4_io_outputs_1_rData_rd <= streamFork_4_io_outputs_1_payload_rd;
      streamFork_4_io_outputs_1_rData_write <= streamFork_4_io_outputs_1_payload_write;
      streamFork_4_io_outputs_1_rData_value <= streamFork_4_io_outputs_1_payload_value;
    end
    if(io_port_0_cmd_ready) begin
      io_port_0_cmd_rData_opcode <= io_port_0_cmd_payload_opcode;
      io_port_0_cmd_rData_arg <= io_port_0_cmd_payload_arg;
      io_port_0_cmd_rData_rs1 <= io_port_0_cmd_payload_rs1;
      io_port_0_cmd_rData_rs2 <= io_port_0_cmd_payload_rs2;
      io_port_0_cmd_rData_rs3 <= io_port_0_cmd_payload_rs3;
      io_port_0_cmd_rData_rd <= io_port_0_cmd_payload_rd;
      io_port_0_cmd_rData_format <= io_port_0_cmd_payload_format;
      io_port_0_cmd_rData_roundMode <= io_port_0_cmd_payload_roundMode;
    end
    if(io_port_1_cmd_ready) begin
      io_port_1_cmd_rData_opcode <= io_port_1_cmd_payload_opcode;
      io_port_1_cmd_rData_arg <= io_port_1_cmd_payload_arg;
      io_port_1_cmd_rData_rs1 <= io_port_1_cmd_payload_rs1;
      io_port_1_cmd_rData_rs2 <= io_port_1_cmd_payload_rs2;
      io_port_1_cmd_rData_rs3 <= io_port_1_cmd_payload_rs3;
      io_port_1_cmd_rData_rd <= io_port_1_cmd_payload_rd;
      io_port_1_cmd_rData_format <= io_port_1_cmd_payload_format;
      io_port_1_cmd_rData_roundMode <= io_port_1_cmd_payload_roundMode;
    end
    if(scheduler_0_output_ready) begin
      scheduler_0_output_rData_opcode <= scheduler_0_output_payload_opcode;
      scheduler_0_output_rData_arg <= scheduler_0_output_payload_arg;
      scheduler_0_output_rData_rs1 <= scheduler_0_output_payload_rs1;
      scheduler_0_output_rData_rs2 <= scheduler_0_output_payload_rs2;
      scheduler_0_output_rData_rs3 <= scheduler_0_output_payload_rs3;
      scheduler_0_output_rData_rd <= scheduler_0_output_payload_rd;
      scheduler_0_output_rData_format <= scheduler_0_output_payload_format;
      scheduler_0_output_rData_roundMode <= scheduler_0_output_payload_roundMode;
    end
    if(scheduler_1_output_ready) begin
      scheduler_1_output_rData_opcode <= scheduler_1_output_payload_opcode;
      scheduler_1_output_rData_arg <= scheduler_1_output_payload_arg;
      scheduler_1_output_rData_rs1 <= scheduler_1_output_payload_rs1;
      scheduler_1_output_rData_rs2 <= scheduler_1_output_payload_rs2;
      scheduler_1_output_rData_rs3 <= scheduler_1_output_payload_rs3;
      scheduler_1_output_rData_rd <= scheduler_1_output_payload_rd;
      scheduler_1_output_rData_format <= scheduler_1_output_payload_format;
      scheduler_1_output_rData_roundMode <= scheduler_1_output_payload_roundMode;
    end
    if(read_s0_ready) begin
      read_s0_rData_source <= read_s0_payload_source;
      read_s0_rData_opcode <= read_s0_payload_opcode;
      read_s0_rData_rs1 <= read_s0_payload_rs1;
      read_s0_rData_rs2 <= read_s0_payload_rs2;
      read_s0_rData_rs3 <= read_s0_payload_rs3;
      read_s0_rData_rd <= read_s0_payload_rd;
      read_s0_rData_arg <= read_s0_payload_arg;
      read_s0_rData_roundMode <= read_s0_payload_roundMode;
      read_s0_rData_format <= read_s0_payload_format;
    end
    if(decode_load_ready) begin
      decode_load_rData_source <= decode_load_payload_source;
      decode_load_rData_rd <= decode_load_payload_rd;
      decode_load_rData_i2f <= decode_load_payload_i2f;
      decode_load_rData_arg <= decode_load_payload_arg;
      decode_load_rData_roundMode <= decode_load_payload_roundMode;
      decode_load_rData_format <= decode_load_payload_format;
    end
    if(decode_load_s2mPipe_ready) begin
      decode_load_s2mPipe_rData_source <= decode_load_s2mPipe_payload_source;
      decode_load_s2mPipe_rData_rd <= decode_load_s2mPipe_payload_rd;
      decode_load_s2mPipe_rData_i2f <= decode_load_s2mPipe_payload_i2f;
      decode_load_s2mPipe_rData_arg <= decode_load_s2mPipe_payload_arg;
      decode_load_s2mPipe_rData_roundMode <= decode_load_s2mPipe_payload_roundMode;
      decode_load_s2mPipe_rData_format <= decode_load_s2mPipe_payload_format;
    end
    if(decode_load_s2mPipe_m2sPipe_ready) begin
      decode_load_s2mPipe_m2sPipe_rData_source <= decode_load_s2mPipe_m2sPipe_payload_source;
      decode_load_s2mPipe_m2sPipe_rData_rd <= decode_load_s2mPipe_m2sPipe_payload_rd;
      decode_load_s2mPipe_m2sPipe_rData_i2f <= decode_load_s2mPipe_m2sPipe_payload_i2f;
      decode_load_s2mPipe_m2sPipe_rData_arg <= decode_load_s2mPipe_m2sPipe_payload_arg;
      decode_load_s2mPipe_m2sPipe_rData_roundMode <= decode_load_s2mPipe_m2sPipe_payload_roundMode;
      decode_load_s2mPipe_m2sPipe_rData_format <= decode_load_s2mPipe_m2sPipe_payload_format;
    end
    if(load_s0_output_ready) begin
      load_s0_output_rData_source <= load_s0_output_payload_source;
      load_s0_output_rData_rd <= load_s0_output_payload_rd;
      load_s0_output_rData_value <= load_s0_output_payload_value;
      load_s0_output_rData_i2f <= load_s0_output_payload_i2f;
      load_s0_output_rData_arg <= load_s0_output_payload_arg;
      load_s0_output_rData_roundMode <= load_s0_output_payload_roundMode;
      load_s0_output_rData_format <= load_s0_output_payload_format;
    end
    if(when_FpuCore_l525) begin
      load_s1_fsm_shift_output <= load_s1_fsm_shift_input_6;
    end
    if(when_FpuCore_l529) begin
      if(load_s1_fsm_boot) begin
        if(when_FpuCore_l532) begin
          load_s0_output_rData_value[31 : 0] <= _zz_load_s0_output_rData_value_2;
          load_s1_fsm_patched <= 1'b1;
        end else begin
          load_s1_fsm_shift_by <= {_zz_load_s1_fsm_shift_by_52,{_zz_load_s1_fsm_shift_by_51,{_zz_load_s1_fsm_shift_by_50,{_zz_load_s1_fsm_shift_by_49,{_zz_load_s1_fsm_shift_by_48,_zz_load_s1_fsm_shift_by_47}}}}};
          load_s1_fsm_boot <= 1'b0;
          load_s1_fsm_i2fZero <= (load_s1_input_payload_value[31 : 0] == 32'h0);
        end
      end else begin
        load_s1_fsm_done <= 1'b1;
      end
    end
    if(when_FpuCore_l551) begin
      load_s1_fsm_done <= 1'b0;
      load_s1_fsm_boot <= 1'b1;
      load_s1_fsm_patched <= 1'b0;
    end
    if(decode_shortPip_ready) begin
      decode_shortPip_rData_source <= decode_shortPip_payload_source;
      decode_shortPip_rData_opcode <= decode_shortPip_payload_opcode;
      decode_shortPip_rData_rs1_mantissa <= decode_shortPip_payload_rs1_mantissa;
      decode_shortPip_rData_rs1_exponent <= decode_shortPip_payload_rs1_exponent;
      decode_shortPip_rData_rs1_sign <= decode_shortPip_payload_rs1_sign;
      decode_shortPip_rData_rs1_special <= decode_shortPip_payload_rs1_special;
      decode_shortPip_rData_rs2_mantissa <= decode_shortPip_payload_rs2_mantissa;
      decode_shortPip_rData_rs2_exponent <= decode_shortPip_payload_rs2_exponent;
      decode_shortPip_rData_rs2_sign <= decode_shortPip_payload_rs2_sign;
      decode_shortPip_rData_rs2_special <= decode_shortPip_payload_rs2_special;
      decode_shortPip_rData_rd <= decode_shortPip_payload_rd;
      decode_shortPip_rData_value <= decode_shortPip_payload_value;
      decode_shortPip_rData_arg <= decode_shortPip_payload_arg;
      decode_shortPip_rData_roundMode <= decode_shortPip_payload_roundMode;
      decode_shortPip_rData_format <= decode_shortPip_payload_format;
      decode_shortPip_rData_rs1Boxed <= decode_shortPip_payload_rs1Boxed;
      decode_shortPip_rData_rs2Boxed <= decode_shortPip_payload_rs2Boxed;
    end
    if(when_FpuCore_l646) begin
      shortPip_fsm_shift_scrap <= 1'b1;
    end
    if(when_FpuCore_l646_1) begin
      shortPip_fsm_shift_scrap <= 1'b1;
    end
    if(when_FpuCore_l646_2) begin
      shortPip_fsm_shift_scrap <= 1'b1;
    end
    if(when_FpuCore_l646_3) begin
      shortPip_fsm_shift_scrap <= 1'b1;
    end
    if(when_FpuCore_l646_4) begin
      shortPip_fsm_shift_scrap <= 1'b1;
    end
    if(when_FpuCore_l646_5) begin
      shortPip_fsm_shift_scrap <= 1'b1;
    end
    if(shortPip_fsm_boot) begin
      shortPip_fsm_shift_scrap <= 1'b0;
    end
    if(when_FpuCore_l652) begin
      shortPip_fsm_shift_output <= shortPip_fsm_shift_input_6;
    end
    if(when_FpuCore_l658) begin
      if(shortPip_fsm_boot) begin
        if(shortPip_fsm_isF2i) begin
          shortPip_fsm_shift_by <= _zz_shortPip_fsm_shift_by_2[5:0];
        end else begin
          shortPip_fsm_shift_by <= _zz_shortPip_fsm_shift_by_5[5:0];
        end
        shortPip_fsm_boot <= 1'b0;
      end else begin
        shortPip_fsm_done <= 1'b1;
      end
    end
    if(when_FpuCore_l672) begin
      shortPip_fsm_done <= 1'b0;
      shortPip_fsm_boot <= 1'b1;
    end
    if(shortPip_rspStreams_0_ready) begin
      shortPip_rspStreams_0_rData_value <= shortPip_rspStreams_0_payload_value;
      shortPip_rspStreams_0_rData_NV <= shortPip_rspStreams_0_payload_NV;
      shortPip_rspStreams_0_rData_NX <= shortPip_rspStreams_0_payload_NX;
    end
    if(shortPip_rspStreams_1_ready) begin
      shortPip_rspStreams_1_rData_value <= shortPip_rspStreams_1_payload_value;
      shortPip_rspStreams_1_rData_NV <= shortPip_rspStreams_1_payload_NV;
      shortPip_rspStreams_1_rData_NX <= shortPip_rspStreams_1_payload_NX;
    end
    if(decode_mul_ready) begin
      decode_mul_rData_source <= decode_mul_payload_source;
      decode_mul_rData_rs1_mantissa <= decode_mul_payload_rs1_mantissa;
      decode_mul_rData_rs1_exponent <= decode_mul_payload_rs1_exponent;
      decode_mul_rData_rs1_sign <= decode_mul_payload_rs1_sign;
      decode_mul_rData_rs1_special <= decode_mul_payload_rs1_special;
      decode_mul_rData_rs2_mantissa <= decode_mul_payload_rs2_mantissa;
      decode_mul_rData_rs2_exponent <= decode_mul_payload_rs2_exponent;
      decode_mul_rData_rs2_sign <= decode_mul_payload_rs2_sign;
      decode_mul_rData_rs2_special <= decode_mul_payload_rs2_special;
      decode_mul_rData_rs3_mantissa <= decode_mul_payload_rs3_mantissa;
      decode_mul_rData_rs3_exponent <= decode_mul_payload_rs3_exponent;
      decode_mul_rData_rs3_sign <= decode_mul_payload_rs3_sign;
      decode_mul_rData_rs3_special <= decode_mul_payload_rs3_special;
      decode_mul_rData_rd <= decode_mul_payload_rd;
      decode_mul_rData_add <= decode_mul_payload_add;
      decode_mul_rData_divSqrt <= decode_mul_payload_divSqrt;
      decode_mul_rData_msb1 <= decode_mul_payload_msb1;
      decode_mul_rData_msb2 <= decode_mul_payload_msb2;
      decode_mul_rData_roundMode <= decode_mul_payload_roundMode;
      decode_mul_rData_format <= decode_mul_payload_format;
    end
    if(mul_preMul_output_ready) begin
      mul_preMul_output_rData_source <= mul_preMul_output_payload_source;
      mul_preMul_output_rData_rs1_mantissa <= mul_preMul_output_payload_rs1_mantissa;
      mul_preMul_output_rData_rs1_exponent <= mul_preMul_output_payload_rs1_exponent;
      mul_preMul_output_rData_rs1_sign <= mul_preMul_output_payload_rs1_sign;
      mul_preMul_output_rData_rs1_special <= mul_preMul_output_payload_rs1_special;
      mul_preMul_output_rData_rs2_mantissa <= mul_preMul_output_payload_rs2_mantissa;
      mul_preMul_output_rData_rs2_exponent <= mul_preMul_output_payload_rs2_exponent;
      mul_preMul_output_rData_rs2_sign <= mul_preMul_output_payload_rs2_sign;
      mul_preMul_output_rData_rs2_special <= mul_preMul_output_payload_rs2_special;
      mul_preMul_output_rData_rs3_mantissa <= mul_preMul_output_payload_rs3_mantissa;
      mul_preMul_output_rData_rs3_exponent <= mul_preMul_output_payload_rs3_exponent;
      mul_preMul_output_rData_rs3_sign <= mul_preMul_output_payload_rs3_sign;
      mul_preMul_output_rData_rs3_special <= mul_preMul_output_payload_rs3_special;
      mul_preMul_output_rData_rd <= mul_preMul_output_payload_rd;
      mul_preMul_output_rData_add <= mul_preMul_output_payload_add;
      mul_preMul_output_rData_divSqrt <= mul_preMul_output_payload_divSqrt;
      mul_preMul_output_rData_msb1 <= mul_preMul_output_payload_msb1;
      mul_preMul_output_rData_msb2 <= mul_preMul_output_payload_msb2;
      mul_preMul_output_rData_roundMode <= mul_preMul_output_payload_roundMode;
      mul_preMul_output_rData_format <= mul_preMul_output_payload_format;
      mul_preMul_output_rData_exp <= mul_preMul_output_payload_exp;
    end
    if(mul_mul_output_ready) begin
      mul_mul_output_rData_source <= mul_mul_output_payload_source;
      mul_mul_output_rData_rs1_mantissa <= mul_mul_output_payload_rs1_mantissa;
      mul_mul_output_rData_rs1_exponent <= mul_mul_output_payload_rs1_exponent;
      mul_mul_output_rData_rs1_sign <= mul_mul_output_payload_rs1_sign;
      mul_mul_output_rData_rs1_special <= mul_mul_output_payload_rs1_special;
      mul_mul_output_rData_rs2_mantissa <= mul_mul_output_payload_rs2_mantissa;
      mul_mul_output_rData_rs2_exponent <= mul_mul_output_payload_rs2_exponent;
      mul_mul_output_rData_rs2_sign <= mul_mul_output_payload_rs2_sign;
      mul_mul_output_rData_rs2_special <= mul_mul_output_payload_rs2_special;
      mul_mul_output_rData_rs3_mantissa <= mul_mul_output_payload_rs3_mantissa;
      mul_mul_output_rData_rs3_exponent <= mul_mul_output_payload_rs3_exponent;
      mul_mul_output_rData_rs3_sign <= mul_mul_output_payload_rs3_sign;
      mul_mul_output_rData_rs3_special <= mul_mul_output_payload_rs3_special;
      mul_mul_output_rData_rd <= mul_mul_output_payload_rd;
      mul_mul_output_rData_add <= mul_mul_output_payload_add;
      mul_mul_output_rData_divSqrt <= mul_mul_output_payload_divSqrt;
      mul_mul_output_rData_msb1 <= mul_mul_output_payload_msb1;
      mul_mul_output_rData_msb2 <= mul_mul_output_payload_msb2;
      mul_mul_output_rData_roundMode <= mul_mul_output_payload_roundMode;
      mul_mul_output_rData_format <= mul_mul_output_payload_format;
      mul_mul_output_rData_exp <= mul_mul_output_payload_exp;
      mul_mul_output_rData_muls_0 <= mul_mul_output_payload_muls_0;
      mul_mul_output_rData_muls_1 <= mul_mul_output_payload_muls_1;
      mul_mul_output_rData_muls_2 <= mul_mul_output_payload_muls_2;
      mul_mul_output_rData_muls_3 <= mul_mul_output_payload_muls_3;
      mul_mul_output_rData_muls_4 <= mul_mul_output_payload_muls_4;
      mul_mul_output_rData_muls_5 <= mul_mul_output_payload_muls_5;
      mul_mul_output_rData_muls_6 <= mul_mul_output_payload_muls_6;
      mul_mul_output_rData_muls_7 <= mul_mul_output_payload_muls_7;
      mul_mul_output_rData_muls_8 <= mul_mul_output_payload_muls_8;
    end
    if(mul_sum1_output_ready) begin
      mul_sum1_output_rData_source <= mul_sum1_output_payload_source;
      mul_sum1_output_rData_rs1_mantissa <= mul_sum1_output_payload_rs1_mantissa;
      mul_sum1_output_rData_rs1_exponent <= mul_sum1_output_payload_rs1_exponent;
      mul_sum1_output_rData_rs1_sign <= mul_sum1_output_payload_rs1_sign;
      mul_sum1_output_rData_rs1_special <= mul_sum1_output_payload_rs1_special;
      mul_sum1_output_rData_rs2_mantissa <= mul_sum1_output_payload_rs2_mantissa;
      mul_sum1_output_rData_rs2_exponent <= mul_sum1_output_payload_rs2_exponent;
      mul_sum1_output_rData_rs2_sign <= mul_sum1_output_payload_rs2_sign;
      mul_sum1_output_rData_rs2_special <= mul_sum1_output_payload_rs2_special;
      mul_sum1_output_rData_rs3_mantissa <= mul_sum1_output_payload_rs3_mantissa;
      mul_sum1_output_rData_rs3_exponent <= mul_sum1_output_payload_rs3_exponent;
      mul_sum1_output_rData_rs3_sign <= mul_sum1_output_payload_rs3_sign;
      mul_sum1_output_rData_rs3_special <= mul_sum1_output_payload_rs3_special;
      mul_sum1_output_rData_rd <= mul_sum1_output_payload_rd;
      mul_sum1_output_rData_add <= mul_sum1_output_payload_add;
      mul_sum1_output_rData_divSqrt <= mul_sum1_output_payload_divSqrt;
      mul_sum1_output_rData_msb1 <= mul_sum1_output_payload_msb1;
      mul_sum1_output_rData_msb2 <= mul_sum1_output_payload_msb2;
      mul_sum1_output_rData_roundMode <= mul_sum1_output_payload_roundMode;
      mul_sum1_output_rData_format <= mul_sum1_output_payload_format;
      mul_sum1_output_rData_exp <= mul_sum1_output_payload_exp;
      mul_sum1_output_rData_muls2_0 <= mul_sum1_output_payload_muls2_0;
      mul_sum1_output_rData_muls2_1 <= mul_sum1_output_payload_muls2_1;
      mul_sum1_output_rData_muls2_2 <= mul_sum1_output_payload_muls2_2;
      mul_sum1_output_rData_muls2_3 <= mul_sum1_output_payload_muls2_3;
      mul_sum1_output_rData_muls2_4 <= mul_sum1_output_payload_muls2_4;
      mul_sum1_output_rData_mulC2 <= mul_sum1_output_payload_mulC2;
    end
    if(mul_sum2_output_ready) begin
      mul_sum2_output_rData_source <= mul_sum2_output_payload_source;
      mul_sum2_output_rData_rs1_mantissa <= mul_sum2_output_payload_rs1_mantissa;
      mul_sum2_output_rData_rs1_exponent <= mul_sum2_output_payload_rs1_exponent;
      mul_sum2_output_rData_rs1_sign <= mul_sum2_output_payload_rs1_sign;
      mul_sum2_output_rData_rs1_special <= mul_sum2_output_payload_rs1_special;
      mul_sum2_output_rData_rs2_mantissa <= mul_sum2_output_payload_rs2_mantissa;
      mul_sum2_output_rData_rs2_exponent <= mul_sum2_output_payload_rs2_exponent;
      mul_sum2_output_rData_rs2_sign <= mul_sum2_output_payload_rs2_sign;
      mul_sum2_output_rData_rs2_special <= mul_sum2_output_payload_rs2_special;
      mul_sum2_output_rData_rs3_mantissa <= mul_sum2_output_payload_rs3_mantissa;
      mul_sum2_output_rData_rs3_exponent <= mul_sum2_output_payload_rs3_exponent;
      mul_sum2_output_rData_rs3_sign <= mul_sum2_output_payload_rs3_sign;
      mul_sum2_output_rData_rs3_special <= mul_sum2_output_payload_rs3_special;
      mul_sum2_output_rData_rd <= mul_sum2_output_payload_rd;
      mul_sum2_output_rData_add <= mul_sum2_output_payload_add;
      mul_sum2_output_rData_divSqrt <= mul_sum2_output_payload_divSqrt;
      mul_sum2_output_rData_msb1 <= mul_sum2_output_payload_msb1;
      mul_sum2_output_rData_msb2 <= mul_sum2_output_payload_msb2;
      mul_sum2_output_rData_roundMode <= mul_sum2_output_payload_roundMode;
      mul_sum2_output_rData_format <= mul_sum2_output_payload_format;
      mul_sum2_output_rData_exp <= mul_sum2_output_payload_exp;
      mul_sum2_output_rData_mulC <= mul_sum2_output_payload_mulC;
    end
    if(mul_result_mulToAdd_ready) begin
      mul_result_mulToAdd_rData_source <= mul_result_mulToAdd_payload_source;
      mul_result_mulToAdd_rData_rs1_mantissa <= mul_result_mulToAdd_payload_rs1_mantissa;
      mul_result_mulToAdd_rData_rs1_exponent <= mul_result_mulToAdd_payload_rs1_exponent;
      mul_result_mulToAdd_rData_rs1_sign <= mul_result_mulToAdd_payload_rs1_sign;
      mul_result_mulToAdd_rData_rs1_special <= mul_result_mulToAdd_payload_rs1_special;
      mul_result_mulToAdd_rData_rs2_mantissa <= mul_result_mulToAdd_payload_rs2_mantissa;
      mul_result_mulToAdd_rData_rs2_exponent <= mul_result_mulToAdd_payload_rs2_exponent;
      mul_result_mulToAdd_rData_rs2_sign <= mul_result_mulToAdd_payload_rs2_sign;
      mul_result_mulToAdd_rData_rs2_special <= mul_result_mulToAdd_payload_rs2_special;
      mul_result_mulToAdd_rData_rd <= mul_result_mulToAdd_payload_rd;
      mul_result_mulToAdd_rData_roundMode <= mul_result_mulToAdd_payload_roundMode;
      mul_result_mulToAdd_rData_format <= mul_result_mulToAdd_payload_format;
      mul_result_mulToAdd_rData_needCommit <= mul_result_mulToAdd_payload_needCommit;
    end
    if(decode_div_ready) begin
      decode_div_rData_source <= decode_div_payload_source;
      decode_div_rData_rs1_mantissa <= decode_div_payload_rs1_mantissa;
      decode_div_rData_rs1_exponent <= decode_div_payload_rs1_exponent;
      decode_div_rData_rs1_sign <= decode_div_payload_rs1_sign;
      decode_div_rData_rs1_special <= decode_div_payload_rs1_special;
      decode_div_rData_rs2_mantissa <= decode_div_payload_rs2_mantissa;
      decode_div_rData_rs2_exponent <= decode_div_payload_rs2_exponent;
      decode_div_rData_rs2_sign <= decode_div_payload_rs2_sign;
      decode_div_rData_rs2_special <= decode_div_payload_rs2_special;
      decode_div_rData_rd <= decode_div_payload_rd;
      decode_div_rData_roundMode <= decode_div_payload_roundMode;
      decode_div_rData_format <= decode_div_payload_format;
    end
    div_isCommited <= _zz_div_isCommited;
    if(decode_sqrt_ready) begin
      decode_sqrt_rData_source <= decode_sqrt_payload_source;
      decode_sqrt_rData_rs1_mantissa <= decode_sqrt_payload_rs1_mantissa;
      decode_sqrt_rData_rs1_exponent <= decode_sqrt_payload_rs1_exponent;
      decode_sqrt_rData_rs1_sign <= decode_sqrt_payload_rs1_sign;
      decode_sqrt_rData_rs1_special <= decode_sqrt_payload_rs1_special;
      decode_sqrt_rData_rd <= decode_sqrt_payload_rd;
      decode_sqrt_rData_roundMode <= decode_sqrt_payload_roundMode;
      decode_sqrt_rData_format <= decode_sqrt_payload_format;
    end
    sqrt_isCommited <= _zz_sqrt_isCommited;
    sqrt_exponent <= (_zz_sqrt_exponent + _zz_sqrt_exponent_4);
    if(add_preShifter_output_ready) begin
      add_preShifter_output_rData_source <= add_preShifter_output_payload_source;
      add_preShifter_output_rData_rs1_mantissa <= add_preShifter_output_payload_rs1_mantissa;
      add_preShifter_output_rData_rs1_exponent <= add_preShifter_output_payload_rs1_exponent;
      add_preShifter_output_rData_rs1_sign <= add_preShifter_output_payload_rs1_sign;
      add_preShifter_output_rData_rs1_special <= add_preShifter_output_payload_rs1_special;
      add_preShifter_output_rData_rs2_mantissa <= add_preShifter_output_payload_rs2_mantissa;
      add_preShifter_output_rData_rs2_exponent <= add_preShifter_output_payload_rs2_exponent;
      add_preShifter_output_rData_rs2_sign <= add_preShifter_output_payload_rs2_sign;
      add_preShifter_output_rData_rs2_special <= add_preShifter_output_payload_rs2_special;
      add_preShifter_output_rData_rd <= add_preShifter_output_payload_rd;
      add_preShifter_output_rData_roundMode <= add_preShifter_output_payload_roundMode;
      add_preShifter_output_rData_format <= add_preShifter_output_payload_format;
      add_preShifter_output_rData_needCommit <= add_preShifter_output_payload_needCommit;
      add_preShifter_output_rData_absRs1Bigger <= add_preShifter_output_payload_absRs1Bigger;
      add_preShifter_output_rData_rs1ExponentBigger <= add_preShifter_output_payload_rs1ExponentBigger;
    end
    if(add_shifter_output_ready) begin
      add_shifter_output_rData_source <= add_shifter_output_payload_source;
      add_shifter_output_rData_rs1_mantissa <= add_shifter_output_payload_rs1_mantissa;
      add_shifter_output_rData_rs1_exponent <= add_shifter_output_payload_rs1_exponent;
      add_shifter_output_rData_rs1_sign <= add_shifter_output_payload_rs1_sign;
      add_shifter_output_rData_rs1_special <= add_shifter_output_payload_rs1_special;
      add_shifter_output_rData_rs2_mantissa <= add_shifter_output_payload_rs2_mantissa;
      add_shifter_output_rData_rs2_exponent <= add_shifter_output_payload_rs2_exponent;
      add_shifter_output_rData_rs2_sign <= add_shifter_output_payload_rs2_sign;
      add_shifter_output_rData_rs2_special <= add_shifter_output_payload_rs2_special;
      add_shifter_output_rData_rd <= add_shifter_output_payload_rd;
      add_shifter_output_rData_roundMode <= add_shifter_output_payload_roundMode;
      add_shifter_output_rData_format <= add_shifter_output_payload_format;
      add_shifter_output_rData_needCommit <= add_shifter_output_payload_needCommit;
      add_shifter_output_rData_xSign <= add_shifter_output_payload_xSign;
      add_shifter_output_rData_ySign <= add_shifter_output_payload_ySign;
      add_shifter_output_rData_xMantissa <= add_shifter_output_payload_xMantissa;
      add_shifter_output_rData_yMantissa <= add_shifter_output_payload_yMantissa;
      add_shifter_output_rData_xyExponent <= add_shifter_output_payload_xyExponent;
      add_shifter_output_rData_xySign <= add_shifter_output_payload_xySign;
      add_shifter_output_rData_roundingScrap <= add_shifter_output_payload_roundingScrap;
    end
    if(add_math_output_ready) begin
      add_math_output_rData_source <= add_math_output_payload_source;
      add_math_output_rData_rs1_mantissa <= add_math_output_payload_rs1_mantissa;
      add_math_output_rData_rs1_exponent <= add_math_output_payload_rs1_exponent;
      add_math_output_rData_rs1_sign <= add_math_output_payload_rs1_sign;
      add_math_output_rData_rs1_special <= add_math_output_payload_rs1_special;
      add_math_output_rData_rs2_mantissa <= add_math_output_payload_rs2_mantissa;
      add_math_output_rData_rs2_exponent <= add_math_output_payload_rs2_exponent;
      add_math_output_rData_rs2_sign <= add_math_output_payload_rs2_sign;
      add_math_output_rData_rs2_special <= add_math_output_payload_rs2_special;
      add_math_output_rData_rd <= add_math_output_payload_rd;
      add_math_output_rData_roundMode <= add_math_output_payload_roundMode;
      add_math_output_rData_format <= add_math_output_payload_format;
      add_math_output_rData_needCommit <= add_math_output_payload_needCommit;
      add_math_output_rData_xSign <= add_math_output_payload_xSign;
      add_math_output_rData_ySign <= add_math_output_payload_ySign;
      add_math_output_rData_xMantissa <= add_math_output_payload_xMantissa;
      add_math_output_rData_yMantissa <= add_math_output_payload_yMantissa;
      add_math_output_rData_xyExponent <= add_math_output_payload_xyExponent;
      add_math_output_rData_xySign <= add_math_output_payload_xySign;
      add_math_output_rData_roundingScrap <= add_math_output_payload_roundingScrap;
      add_math_output_rData_xyMantissa <= add_math_output_payload_xyMantissa;
    end
    if(add_oh_output_ready) begin
      add_oh_output_rData_source <= add_oh_output_payload_source;
      add_oh_output_rData_rs1_mantissa <= add_oh_output_payload_rs1_mantissa;
      add_oh_output_rData_rs1_exponent <= add_oh_output_payload_rs1_exponent;
      add_oh_output_rData_rs1_sign <= add_oh_output_payload_rs1_sign;
      add_oh_output_rData_rs1_special <= add_oh_output_payload_rs1_special;
      add_oh_output_rData_rs2_mantissa <= add_oh_output_payload_rs2_mantissa;
      add_oh_output_rData_rs2_exponent <= add_oh_output_payload_rs2_exponent;
      add_oh_output_rData_rs2_sign <= add_oh_output_payload_rs2_sign;
      add_oh_output_rData_rs2_special <= add_oh_output_payload_rs2_special;
      add_oh_output_rData_rd <= add_oh_output_payload_rd;
      add_oh_output_rData_roundMode <= add_oh_output_payload_roundMode;
      add_oh_output_rData_format <= add_oh_output_payload_format;
      add_oh_output_rData_needCommit <= add_oh_output_payload_needCommit;
      add_oh_output_rData_xSign <= add_oh_output_payload_xSign;
      add_oh_output_rData_ySign <= add_oh_output_payload_ySign;
      add_oh_output_rData_xMantissa <= add_oh_output_payload_xMantissa;
      add_oh_output_rData_yMantissa <= add_oh_output_payload_yMantissa;
      add_oh_output_rData_xyExponent <= add_oh_output_payload_xyExponent;
      add_oh_output_rData_xySign <= add_oh_output_payload_xySign;
      add_oh_output_rData_roundingScrap <= add_oh_output_payload_roundingScrap;
      add_oh_output_rData_xyMantissa <= add_oh_output_payload_xyMantissa;
      add_oh_output_rData_shift <= add_oh_output_payload_shift;
    end
    if(load_s1_output_ready) begin
      load_s1_output_rData_source <= load_s1_output_payload_source;
      load_s1_output_rData_rd <= load_s1_output_payload_rd;
      load_s1_output_rData_value_mantissa <= load_s1_output_payload_value_mantissa;
      load_s1_output_rData_value_exponent <= load_s1_output_payload_value_exponent;
      load_s1_output_rData_value_sign <= load_s1_output_payload_value_sign;
      load_s1_output_rData_value_special <= load_s1_output_payload_value_special;
      load_s1_output_rData_scrap <= load_s1_output_payload_scrap;
      load_s1_output_rData_roundMode <= load_s1_output_payload_roundMode;
      load_s1_output_rData_format <= load_s1_output_payload_format;
      load_s1_output_rData_NV <= load_s1_output_payload_NV;
      load_s1_output_rData_DZ <= load_s1_output_payload_DZ;
    end
    if(shortPip_output_ready) begin
      shortPip_output_rData_source <= shortPip_output_payload_source;
      shortPip_output_rData_rd <= shortPip_output_payload_rd;
      shortPip_output_rData_value_mantissa <= shortPip_output_payload_value_mantissa;
      shortPip_output_rData_value_exponent <= shortPip_output_payload_value_exponent;
      shortPip_output_rData_value_sign <= shortPip_output_payload_value_sign;
      shortPip_output_rData_value_special <= shortPip_output_payload_value_special;
      shortPip_output_rData_scrap <= shortPip_output_payload_scrap;
      shortPip_output_rData_roundMode <= shortPip_output_payload_roundMode;
      shortPip_output_rData_format <= shortPip_output_payload_format;
      shortPip_output_rData_NV <= shortPip_output_payload_NV;
      shortPip_output_rData_DZ <= shortPip_output_payload_DZ;
    end
    roundFront_input_payload_source <= merge_arbitrated_payload_source;
    roundFront_input_payload_rd <= merge_arbitrated_payload_rd;
    roundFront_input_payload_value_mantissa <= merge_arbitrated_payload_value_mantissa;
    roundFront_input_payload_value_exponent <= merge_arbitrated_payload_value_exponent;
    roundFront_input_payload_value_sign <= merge_arbitrated_payload_value_sign;
    roundFront_input_payload_value_special <= merge_arbitrated_payload_value_special;
    roundFront_input_payload_scrap <= merge_arbitrated_payload_scrap;
    roundFront_input_payload_roundMode <= merge_arbitrated_payload_roundMode;
    roundFront_input_payload_format <= merge_arbitrated_payload_format;
    roundFront_input_payload_NV <= merge_arbitrated_payload_NV;
    roundFront_input_payload_DZ <= merge_arbitrated_payload_DZ;
    roundBack_input_payload_source <= roundFront_output_payload_source;
    roundBack_input_payload_rd <= roundFront_output_payload_rd;
    roundBack_input_payload_value_mantissa <= roundFront_output_payload_value_mantissa;
    roundBack_input_payload_value_exponent <= roundFront_output_payload_value_exponent;
    roundBack_input_payload_value_sign <= roundFront_output_payload_value_sign;
    roundBack_input_payload_value_special <= roundFront_output_payload_value_special;
    roundBack_input_payload_scrap <= roundFront_output_payload_scrap;
    roundBack_input_payload_roundMode <= roundFront_output_payload_roundMode;
    roundBack_input_payload_format <= roundFront_output_payload_format;
    roundBack_input_payload_NV <= roundFront_output_payload_NV;
    roundBack_input_payload_DZ <= roundFront_output_payload_DZ;
    roundBack_input_payload_mantissaIncrement <= roundFront_output_payload_mantissaIncrement;
    roundBack_input_payload_roundAdjusted <= roundFront_output_payload_roundAdjusted;
    roundBack_input_payload_exactMask <= roundFront_output_payload_exactMask;
    writeback_input_payload_source <= roundBack_output_payload_source;
    writeback_input_payload_rd <= roundBack_output_payload_rd;
    writeback_input_payload_value_mantissa <= roundBack_output_payload_value_mantissa;
    writeback_input_payload_value_exponent <= roundBack_output_payload_value_exponent;
    writeback_input_payload_value_sign <= roundBack_output_payload_value_sign;
    writeback_input_payload_value_special <= roundBack_output_payload_value_special;
    writeback_input_payload_format <= roundBack_output_payload_format;
    writeback_input_payload_NV <= roundBack_output_payload_NV;
    writeback_input_payload_NX <= roundBack_output_payload_NX;
    writeback_input_payload_OF <= roundBack_output_payload_OF;
    writeback_input_payload_UF <= roundBack_output_payload_UF;
    writeback_input_payload_DZ <= roundBack_output_payload_DZ;
    writeback_input_payload_write <= roundBack_output_payload_write;
  end


endmodule

module VexRiscv_1 (
  output wire          dBus_cmd_valid,
  input  wire          dBus_cmd_ready,
  output wire          dBus_cmd_payload_wr,
  output wire          dBus_cmd_payload_uncached,
  output wire [31:0]   dBus_cmd_payload_address,
  output wire [63:0]   dBus_cmd_payload_data,
  output wire [7:0]    dBus_cmd_payload_mask,
  output wire [2:0]    dBus_cmd_payload_size,
  output wire          dBus_cmd_payload_exclusive,
  output wire          dBus_cmd_payload_last,
  input  wire          dBus_rsp_valid,
  input  wire [3:0]    dBus_rsp_payload_aggregated,
  input  wire          dBus_rsp_payload_last,
  input  wire [63:0]   dBus_rsp_payload_data,
  input  wire          dBus_rsp_payload_error,
  input  wire          dBus_rsp_payload_exclusive,
  input  wire          dBus_inv_valid,
  output wire          dBus_inv_ready,
  input  wire          dBus_inv_payload_last,
  input  wire          dBus_inv_payload_fragment_enable,
  input  wire [31:0]   dBus_inv_payload_fragment_address,
  output wire          dBus_ack_valid,
  input  wire          dBus_ack_ready,
  output wire          dBus_ack_payload_last,
  output wire          dBus_ack_payload_fragment_hit,
  input  wire          dBus_sync_valid,
  output wire          dBus_sync_ready,
  input  wire [3:0]    dBus_sync_payload_aggregated,
  input  wire          timerInterrupt,
  input  wire          externalInterrupt,
  input  wire          softwareInterrupt,
  output wire          debugBus_halted,
  output wire          debugBus_running,
  output wire          debugBus_unavailable,
  output reg           debugBus_exception,
  output wire          debugBus_commit,
  output reg           debugBus_ebreak,
  output wire          debugBus_redo,
  output wire          debugBus_regSuccess,
  input  wire          debugBus_ackReset,
  output wire          debugBus_haveReset,
  input  wire          debugBus_resume_cmd_valid,
  output reg           debugBus_resume_rsp_valid,
  input  wire          debugBus_haltReq,
  input  wire          debugBus_dmToHart_valid,
  input  wire [1:0]    debugBus_dmToHart_payload_op,
  input  wire [4:0]    debugBus_dmToHart_payload_address,
  input  wire [31:0]   debugBus_dmToHart_payload_data,
  input  wire [2:0]    debugBus_dmToHart_payload_size,
  output reg           debugBus_hartToDm_valid,
  output reg  [3:0]    debugBus_hartToDm_payload_address,
  output reg  [31:0]   debugBus_hartToDm_payload_data,
  output reg           FpuPlugin_port_cmd_valid /* verilator public */ ,
  input  wire          FpuPlugin_port_cmd_ready /* verilator public */ ,
  output reg  [3:0]    FpuPlugin_port_cmd_payload_opcode /* verilator public */ ,
  output wire [1:0]    FpuPlugin_port_cmd_payload_arg /* verilator public */ ,
  output wire [4:0]    FpuPlugin_port_cmd_payload_rs1 /* verilator public */ ,
  output reg  [4:0]    FpuPlugin_port_cmd_payload_rs2 /* verilator public */ ,
  output wire [4:0]    FpuPlugin_port_cmd_payload_rs3 /* verilator public */ ,
  output reg  [4:0]    FpuPlugin_port_cmd_payload_rd /* verilator public */ ,
  output reg  [0:0]    FpuPlugin_port_cmd_payload_format /* verilator public */ ,
  output wire [2:0]    FpuPlugin_port_cmd_payload_roundMode /* verilator public */ ,
  output reg           FpuPlugin_port_commit_valid /* verilator public */ ,
  input  wire          FpuPlugin_port_commit_ready /* verilator public */ ,
  output reg  [3:0]    FpuPlugin_port_commit_payload_opcode /* verilator public */ ,
  output reg  [4:0]    FpuPlugin_port_commit_payload_rd /* verilator public */ ,
  output reg           FpuPlugin_port_commit_payload_write /* verilator public */ ,
  output reg  [63:0]   FpuPlugin_port_commit_payload_value /* verilator public */ ,
  input  wire          FpuPlugin_port_rsp_valid /* verilator public */ ,
  output reg           FpuPlugin_port_rsp_ready /* verilator public */ ,
  input  wire [63:0]   FpuPlugin_port_rsp_payload_value /* verilator public */ ,
  input  wire          FpuPlugin_port_rsp_payload_NV /* verilator public */ ,
  input  wire          FpuPlugin_port_rsp_payload_NX /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_valid /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_NX /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_UF /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_OF /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_DZ /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_NV /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_written /* verilator public */ ,
  output wire          CfuPlugin_bus_cmd_valid,
  input  wire          CfuPlugin_bus_cmd_ready,
  output wire [9:0]    CfuPlugin_bus_cmd_payload_function_id,
  output wire [31:0]   CfuPlugin_bus_cmd_payload_inputs_0,
  output wire [31:0]   CfuPlugin_bus_cmd_payload_inputs_1,
  input  wire          CfuPlugin_bus_rsp_valid,
  output wire          CfuPlugin_bus_rsp_ready,
  input  wire [31:0]   CfuPlugin_bus_rsp_payload_outputs_0,
  output wire          iBus_cmd_valid,
  input  wire          iBus_cmd_ready,
  output reg  [31:0]   iBus_cmd_payload_address,
  output wire [2:0]    iBus_cmd_payload_size,
  input  wire          iBus_rsp_valid,
  input  wire [63:0]   iBus_rsp_payload_data,
  input  wire          iBus_rsp_payload_error,
  input  wire          systemCd_logic_outputReset,
  output reg           stoptime,
  input  wire          io_systemClk
);
  localparam FpuOpcode_LOAD = 4'd0;
  localparam FpuOpcode_STORE = 4'd1;
  localparam FpuOpcode_MUL = 4'd2;
  localparam FpuOpcode_ADD = 4'd3;
  localparam FpuOpcode_FMA = 4'd4;
  localparam FpuOpcode_I2F = 4'd5;
  localparam FpuOpcode_F2I = 4'd6;
  localparam FpuOpcode_CMP = 4'd7;
  localparam FpuOpcode_DIV = 4'd8;
  localparam FpuOpcode_SQRT = 4'd9;
  localparam FpuOpcode_MIN_MAX = 4'd10;
  localparam FpuOpcode_SGNJ = 4'd11;
  localparam FpuOpcode_FMV_X_W = 4'd12;
  localparam FpuOpcode_FMV_W_X = 4'd13;
  localparam FpuOpcode_FCLASS = 4'd14;
  localparam FpuOpcode_FCVT_X_X = 4'd15;
  localparam ShiftCtrlEnum_DISABLE_1 = 2'd0;
  localparam ShiftCtrlEnum_SLL_1 = 2'd1;
  localparam ShiftCtrlEnum_SRL_1 = 2'd2;
  localparam ShiftCtrlEnum_SRA_1 = 2'd3;
  localparam AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam Input2Kind_RS = 1'd0;
  localparam Input2Kind_IMM_I = 1'd1;
  localparam BranchCtrlEnum_INC = 2'd0;
  localparam BranchCtrlEnum_B = 2'd1;
  localparam BranchCtrlEnum_JAL = 2'd2;
  localparam BranchCtrlEnum_JALR = 2'd3;
  localparam EnvCtrlEnum_NONE = 2'd0;
  localparam EnvCtrlEnum_XRET = 2'd1;
  localparam EnvCtrlEnum_ECALL = 2'd2;
  localparam EnvCtrlEnum_EBREAK = 2'd3;
  localparam AluCtrlEnum_ADD_SUB = 2'd0;
  localparam AluCtrlEnum_SLT_SLTU = 2'd1;
  localparam AluCtrlEnum_BITWISE = 2'd2;
  localparam FpuFormat_FLOAT = 1'd0;
  localparam FpuFormat_DOUBLE = 1'd1;
  localparam Src2CtrlEnum_RS = 2'd0;
  localparam Src2CtrlEnum_IMI = 2'd1;
  localparam Src2CtrlEnum_IMS = 2'd2;
  localparam Src2CtrlEnum_PC = 2'd3;
  localparam Src1CtrlEnum_RS = 2'd0;
  localparam Src1CtrlEnum_IMU = 2'd1;
  localparam Src1CtrlEnum_PC_INCREMENT = 2'd2;
  localparam Src1CtrlEnum_URS1 = 2'd3;
  localparam DebugDmToHartOp_DATA = 2'd0;
  localparam DebugDmToHartOp_EXECUTE = 2'd1;
  localparam DebugDmToHartOp_REG_WRITE = 2'd2;
  localparam DebugDmToHartOp_REG_READ = 2'd3;
  localparam FpuRoundMode_RNE = 3'd0;
  localparam FpuRoundMode_RTZ = 3'd1;
  localparam FpuRoundMode_RDN = 3'd2;
  localparam FpuRoundMode_RUP = 3'd3;
  localparam FpuRoundMode_RMM = 3'd4;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_BOOT = 2'd0;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_IDLE = 2'd1;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_SINGLE = 2'd2;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 = 2'd3;
  localparam FpuPlugin_enumDef_BOOT = 3'd0;
  localparam FpuPlugin_enumDef_IDLE = 3'd1;
  localparam FpuPlugin_enumDef_CMD = 3'd2;
  localparam FpuPlugin_enumDef_RSP = 3'd3;
  localparam FpuPlugin_enumDef_RSP_0 = 3'd4;
  localparam FpuPlugin_enumDef_RSP_1 = 3'd5;
  localparam FpuPlugin_enumDef_COMMIT = 3'd6;
  localparam FpuPlugin_enumDef_DONE = 3'd7;

  wire                IBusCachedPlugin_cache_io_flush;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isRemoved;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isUser;
  reg                 IBusCachedPlugin_cache_io_cpu_fill_valid;
  wire                dataCache_2_io_cpu_execute_isValid;
  wire       [31:0]   dataCache_2_io_cpu_execute_address;
  reg                 dataCache_2_io_cpu_execute_args_isLrsc;
  wire                dataCache_2_io_cpu_execute_args_amoCtrl_swap;
  wire       [2:0]    dataCache_2_io_cpu_execute_args_amoCtrl_alu;
  wire                dataCache_2_io_cpu_memory_isValid;
  reg                 dataCache_2_io_cpu_memory_mmuRsp_isIoAccess;
  reg                 dataCache_2_io_cpu_writeBack_isValid;
  wire                dataCache_2_io_cpu_writeBack_isUser;
  reg        [63:0]   dataCache_2_io_cpu_writeBack_storeData;
  wire       [31:0]   dataCache_2_io_cpu_writeBack_address;
  reg                 dataCache_2_io_cpu_writeBack_fence_SW;
  reg                 dataCache_2_io_cpu_writeBack_fence_SR;
  reg                 dataCache_2_io_cpu_writeBack_fence_SO;
  reg                 dataCache_2_io_cpu_writeBack_fence_SI;
  reg                 dataCache_2_io_cpu_writeBack_fence_PW;
  reg                 dataCache_2_io_cpu_writeBack_fence_PR;
  reg                 dataCache_2_io_cpu_writeBack_fence_PO;
  reg                 dataCache_2_io_cpu_writeBack_fence_PI;
  wire       [3:0]    dataCache_2_io_cpu_writeBack_fence_FM;
  wire                dataCache_2_io_cpu_flush_valid;
  wire                dataCache_2_io_cpu_flush_payload_singleLine;
  wire       [5:0]    dataCache_2_io_cpu_flush_payload_lineId;
  reg        [31:0]   RegFilePlugin_regFile_spinal_port0;
  reg        [31:0]   RegFilePlugin_regFile_spinal_port1;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_haltIt;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_data;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress;
  wire                IBusCachedPlugin_cache_io_cpu_decode_error;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuException;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_data;
  wire                IBusCachedPlugin_cache_io_cpu_decode_cacheMiss;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_physicalAddress;
  wire                IBusCachedPlugin_cache_io_mem_cmd_valid;
  wire       [31:0]   IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  wire       [2:0]    IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  wire                dataCache_2_io_cpu_execute_haltIt;
  wire                dataCache_2_io_cpu_execute_refilling;
  wire                dataCache_2_io_cpu_memory_isWrite;
  wire                dataCache_2_io_cpu_writeBack_haltIt;
  wire       [63:0]   dataCache_2_io_cpu_writeBack_data;
  wire                dataCache_2_io_cpu_writeBack_mmuException;
  wire                dataCache_2_io_cpu_writeBack_unalignedAccess;
  wire                dataCache_2_io_cpu_writeBack_accessError;
  wire                dataCache_2_io_cpu_writeBack_isWrite;
  wire                dataCache_2_io_cpu_writeBack_keepMemRspData;
  wire                dataCache_2_io_cpu_writeBack_exclusiveOk;
  wire                dataCache_2_io_cpu_flush_ready;
  wire                dataCache_2_io_cpu_redo;
  wire                dataCache_2_io_cpu_writesPending;
  wire                dataCache_2_io_mem_cmd_valid;
  wire                dataCache_2_io_mem_cmd_payload_wr;
  wire                dataCache_2_io_mem_cmd_payload_uncached;
  wire       [31:0]   dataCache_2_io_mem_cmd_payload_address;
  wire       [63:0]   dataCache_2_io_mem_cmd_payload_data;
  wire       [7:0]    dataCache_2_io_mem_cmd_payload_mask;
  wire       [2:0]    dataCache_2_io_mem_cmd_payload_size;
  wire                dataCache_2_io_mem_cmd_payload_exclusive;
  wire                dataCache_2_io_mem_cmd_payload_last;
  wire                dataCache_2_io_mem_inv_ready;
  wire                dataCache_2_io_mem_ack_valid;
  wire                dataCache_2_io_mem_ack_payload_last;
  wire                dataCache_2_io_mem_ack_payload_fragment_hit;
  wire                dataCache_2_io_mem_sync_ready;
  wire                systemCd_logic_outputReset_buffercc_io_dataOut;
  wire       [31:0]   EfxCPUSp1_inst_result;
  wire       [31:0]   EfxCPUSp2_inst_result;
  wire       [51:0]   _zz_memory_MUL_LOW;
  wire       [51:0]   _zz_memory_MUL_LOW_1;
  wire       [51:0]   _zz_memory_MUL_LOW_2;
  wire       [32:0]   _zz_memory_MUL_LOW_3;
  wire       [51:0]   _zz_memory_MUL_LOW_4;
  wire       [49:0]   _zz_memory_MUL_LOW_5;
  wire       [51:0]   _zz_memory_MUL_LOW_6;
  wire       [49:0]   _zz_memory_MUL_LOW_7;
  wire       [31:0]   _zz_decode_FORMAL_PC_NEXT;
  wire       [2:0]    _zz_decode_FORMAL_PC_NEXT_1;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_1;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_2;
  wire                _zz_decode_LEGAL_INSTRUCTION_3;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_4;
  wire       [29:0]   _zz_decode_LEGAL_INSTRUCTION_5;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_6;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_7;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_8;
  wire                _zz_decode_LEGAL_INSTRUCTION_9;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_10;
  wire       [23:0]   _zz_decode_LEGAL_INSTRUCTION_11;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_12;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_13;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_14;
  wire                _zz_decode_LEGAL_INSTRUCTION_15;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_16;
  wire       [17:0]   _zz_decode_LEGAL_INSTRUCTION_17;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_18;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_19;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_20;
  wire                _zz_decode_LEGAL_INSTRUCTION_21;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_22;
  wire       [11:0]   _zz_decode_LEGAL_INSTRUCTION_23;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_24;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_25;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_26;
  wire                _zz_decode_LEGAL_INSTRUCTION_27;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_28;
  wire       [5:0]    _zz_decode_LEGAL_INSTRUCTION_29;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_30;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_31;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_32;
  wire                _zz_decode_LEGAL_INSTRUCTION_33;
  wire                _zz_decode_LEGAL_INSTRUCTION_34;
  wire       [2:0]    _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  reg        [31:0]   _zz_IBusCachedPlugin_jump_pcLoad_payload_4;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_5;
  wire       [31:0]   _zz_IBusCachedPlugin_fetchPc_pc;
  wire       [2:0]    _zz_IBusCachedPlugin_fetchPc_pc_1;
  wire       [31:0]   _zz_IBusCachedPlugin_decodePc_pcPlus;
  wire       [2:0]    _zz_IBusCachedPlugin_decodePc_pcPlus_1;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_28;
  wire       [0:0]    _zz_IBusCachedPlugin_decompressor_decompressed_29;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_30;
  wire       [31:0]   _zz_IBusCachedPlugin_decompressor_decompressed_31;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_32;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_33;
  wire       [6:0]    _zz_IBusCachedPlugin_decompressor_decompressed_34;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_35;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_36;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_37;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_38;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_39;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_40;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_41;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_42;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_43;
  wire       [25:0]   _zz_io_cpu_flush_payload_lineId;
  wire       [25:0]   _zz_io_cpu_flush_payload_lineId_1;
  wire       [2:0]    _zz_DBusCachedPlugin_exceptionBus_payload_code;
  wire       [2:0]    _zz_DBusCachedPlugin_exceptionBus_payload_code_1;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted;
  wire       [2:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_1;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_2;
  wire       [1:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_3;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_4;
  wire       [0:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_5;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_6;
  wire       [0:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_7;
  wire       [0:0]    _zz_writeBack_DBusCachedPlugin_rspRf;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_1;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_2;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_3;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_4;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_5;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_6;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_7;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_8;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_9;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_10;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_11;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_12;
  wire       [40:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_13;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_14;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_15;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_16;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_17;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_18;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_19;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_20;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_21;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_22;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_23;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_24;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_25;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_26;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_27;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_28;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_29;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_30;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_31;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_32;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_33;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_34;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_35;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_36;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_37;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_38;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_39;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_40;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_41;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_42;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_43;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_44;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_45;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_46;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_47;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_48;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_49;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_50;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_51;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_52;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_53;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_54;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_55;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_56;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_57;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_58;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_59;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_60;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_61;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_62;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_63;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_64;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_65;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_66;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_67;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_68;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_69;
  wire       [35:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_70;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_71;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_72;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_73;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_74;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_75;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_76;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_77;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_78;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_79;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_80;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_81;
  wire       [33:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_82;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_83;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_84;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_85;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_86;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_87;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_88;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_89;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_90;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_91;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_92;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_93;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_94;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_95;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_96;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_97;
  wire       [29:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_98;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_99;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_100;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_101;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_102;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_103;
  wire       [27:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_104;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_105;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_106;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_107;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_108;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_109;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_110;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_111;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_112;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_113;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_114;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_115;
  wire       [24:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_116;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_117;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_118;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_119;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_120;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_121;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_122;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_123;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_124;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_125;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_126;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_127;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_128;
  wire       [20:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_129;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_130;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_131;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_132;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_133;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_134;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_135;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_136;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_137;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_138;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_139;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_140;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_141;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_142;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_143;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_144;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_145;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_146;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_147;
  wire       [16:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_148;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_149;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_150;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_151;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_152;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_153;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_154;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_155;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_156;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_157;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_158;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_159;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_160;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_161;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_162;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_163;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_164;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_165;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_166;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_167;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_168;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_169;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_170;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_171;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_172;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_173;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_174;
  wire       [13:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_175;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_176;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_177;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_178;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_179;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_180;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_181;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_182;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_183;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_184;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_185;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_186;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_187;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_188;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_189;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_190;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_191;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_192;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_193;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_194;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_195;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_196;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_197;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_198;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_199;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_200;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_201;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_202;
  wire       [6:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_203;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_204;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_205;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_206;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_207;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_208;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_209;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_210;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_211;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_212;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_213;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_214;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_215;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_216;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_217;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_218;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_219;
  wire       [10:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_220;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_221;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_222;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_223;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_224;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_225;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_226;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_227;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_228;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_229;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_230;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_231;
  wire       [8:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_232;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_233;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_234;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_235;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_236;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_237;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_238;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_239;
  wire       [6:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_240;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_241;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_242;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_243;
  wire       [5:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_244;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_245;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_246;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_247;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_248;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_249;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_250;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_251;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_252;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_253;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_254;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_255;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_256;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_257;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_258;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_259;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_260;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_261;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_262;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_263;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_264;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_265;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_266;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_267;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_268;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_269;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_270;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_271;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_272;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_273;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_274;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_275;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_276;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_277;
  wire                _zz_RegFilePlugin_regFile_port;
  wire                _zz_decode_RegFilePlugin_rs1Data;
  wire                _zz_RegFilePlugin_regFile_port_1;
  wire                _zz_decode_RegFilePlugin_rs2Data;
  wire       [2:0]    _zz__zz_decode_SRC1;
  wire       [4:0]    _zz__zz_decode_SRC1_1;
  wire       [11:0]   _zz__zz_decode_SRC2_2;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_1;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_2;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_4;
  wire       [2:0]    _zz_CsrPlugin_timeout_counter_valueNext;
  wire       [0:0]    _zz_CsrPlugin_timeout_counter_valueNext_1;
  wire       [0:0]    _zz__zz_6;
  wire       [63:0]   _zz_CsrPlugin_counters_mcycle;
  wire       [0:0]    _zz_CsrPlugin_counters_mcycle_1;
  wire       [63:0]   _zz_CsrPlugin_counters_minstret;
  wire       [0:0]    _zz_CsrPlugin_counters_minstret_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1;
  wire                _zz_when;
  wire       [19:0]   _zz__zz_execute_BranchPlugin_branch_src2;
  wire       [11:0]   _zz__zz_execute_BranchPlugin_branch_src2_4;
  wire       [65:0]   _zz_writeBack_MulPlugin_result;
  wire       [65:0]   _zz_writeBack_MulPlugin_result_1;
  wire       [31:0]   _zz__zz_decode_RS2_2;
  wire       [31:0]   _zz__zz_decode_RS2_2_1;
  wire       [5:0]    _zz_memory_MulDivIterativePlugin_div_counter_valueNext;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_div_counter_valueNext_1;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder_1;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_outNumerator;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_1;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_2;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_3;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_4;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_div_result_5;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_rs1_2;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_rs1_3;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_rs2_1;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_rs2_2;
  wire       [5:0]    _zz_FpuPlugin_pendings;
  wire       [5:0]    _zz_FpuPlugin_pendings_1;
  wire       [5:0]    _zz_FpuPlugin_pendings_2;
  wire       [0:0]    _zz_FpuPlugin_pendings_3;
  wire       [5:0]    _zz_FpuPlugin_pendings_4;
  wire       [0:0]    _zz_FpuPlugin_pendings_5;
  wire       [5:0]    _zz_FpuPlugin_pendings_6;
  wire       [0:0]    _zz_FpuPlugin_pendings_7;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_17;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_18;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_19;
  wire       [7:0]    _zz_when_CsrPlugin_l1862;
  wire       [63:0]   writeBack_MEMORY_LOAD_DATA;
  wire       [51:0]   memory_MUL_LOW;
  wire       [31:0]   execute_SHIFT_RIGHT;
  wire       [31:0]   execute_REGFILE_WRITE_DATA;
  wire                memory_CfuPlugin_CFU_IN_FLIGHT;
  wire                execute_CfuPlugin_CFU_IN_FLIGHT;
  wire       [33:0]   memory_MUL_HH;
  wire       [33:0]   execute_MUL_HH;
  wire       [33:0]   execute_MUL_HL;
  wire       [33:0]   execute_MUL_LH;
  wire       [31:0]   execute_MUL_LL;
  wire       [31:0]   execute_BRANCH_CALC;
  wire                execute_BRANCH_DO;
  wire       [31:0]   execute_MEMORY_VIRTUAL_ADDRESS;
  wire       [31:0]   execute_MEMORY_STORE_DATA_RF;
  wire                memory_FPU_COMMIT_LOAD;
  wire                execute_FPU_COMMIT_LOAD;
  wire                decode_FPU_COMMIT_LOAD;
  wire                memory_FPU_FORKED;
  wire                execute_FPU_FORKED;
  wire                decode_FPU_FORKED;
  wire                decode_CSR_READ_OPCODE;
  wire                decode_CSR_WRITE_OPCODE;
  wire       [31:0]   decode_SRC2;
  wire       [31:0]   decode_SRC1;
  wire                decode_SRC2_FORCE_ZERO;
  wire       [31:0]   memory_RS1;
  wire       [1:0]    _zz_execute_to_memory_SHIFT_CTRL;
  wire       [1:0]    _zz_execute_to_memory_SHIFT_CTRL_1;
  wire       [1:0]    decode_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SHIFT_CTRL_1;
  wire       [1:0]    decode_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  wire       [0:0]    decode_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_decode_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1;
  wire                decode_CfuPlugin_CFU_ENABLE;
  wire       [3:0]    memory_FPU_OPCODE;
  wire       [3:0]    _zz_memory_FPU_OPCODE;
  wire       [3:0]    _zz_memory_to_writeBack_FPU_OPCODE;
  wire       [3:0]    _zz_memory_to_writeBack_FPU_OPCODE_1;
  wire       [3:0]    execute_FPU_OPCODE;
  wire       [3:0]    _zz_execute_FPU_OPCODE;
  wire       [3:0]    _zz_execute_to_memory_FPU_OPCODE;
  wire       [3:0]    _zz_execute_to_memory_FPU_OPCODE_1;
  wire       [3:0]    _zz_decode_to_execute_FPU_OPCODE;
  wire       [3:0]    _zz_decode_to_execute_FPU_OPCODE_1;
  wire                memory_FPU_RSP;
  wire                execute_FPU_RSP;
  wire                decode_FPU_RSP;
  wire                memory_FPU_COMMIT;
  wire                execute_FPU_COMMIT;
  wire                decode_FPU_COMMIT;
  wire                decode_IS_RS2_SIGNED;
  wire                decode_IS_RS1_SIGNED;
  wire                decode_IS_DIV;
  wire                memory_IS_MUL;
  wire                decode_IS_MUL;
  wire                decode_SRC_LESS_UNSIGNED;
  wire       [1:0]    decode_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_to_execute_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_to_execute_BRANCH_CTRL_1;
  wire       [1:0]    _zz_memory_to_writeBack_ENV_CTRL;
  wire       [1:0]    _zz_memory_to_writeBack_ENV_CTRL_1;
  wire       [1:0]    _zz_execute_to_memory_ENV_CTRL;
  wire       [1:0]    _zz_execute_to_memory_ENV_CTRL_1;
  wire       [1:0]    decode_ENV_CTRL;
  wire       [1:0]    _zz_decode_ENV_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ENV_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ENV_CTRL_1;
  wire                decode_IS_CSR;
  wire                memory_MEMORY_FENCE;
  wire                execute_MEMORY_FENCE;
  wire                decode_MEMORY_FENCE;
  wire                decode_MEMORY_MANAGMENT;
  wire                memory_MEMORY_AMO;
  wire                memory_MEMORY_LRSC;
  wire                execute_HAS_SIDE_EFFECT;
  wire                decode_HAS_SIDE_EFFECT;
  wire                decode_MEMORY_WR;
  wire                execute_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_EXECUTE_STAGE;
  wire       [1:0]    decode_ALU_CTRL;
  wire       [1:0]    _zz_decode_ALU_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_CTRL_1;
  wire                decode_MEMORY_FENCE_WR;
  wire                decode_MEMORY_FORCE_CONSTISTENCY;
  wire       [31:0]   writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   memory_FORMAL_PC_NEXT;
  wire       [31:0]   execute_FORMAL_PC_NEXT;
  wire       [31:0]   decode_FORMAL_PC_NEXT;
  wire       [31:0]   memory_SHIFT_RIGHT;
  wire       [1:0]    memory_SHIFT_CTRL;
  wire       [1:0]    _zz_memory_SHIFT_CTRL;
  wire       [1:0]    execute_SHIFT_CTRL;
  wire       [1:0]    _zz_execute_SHIFT_CTRL;
  wire       [31:0]   execute_SRC_ADD_SUB;
  wire       [1:0]    execute_ALU_CTRL;
  wire       [1:0]    _zz_execute_ALU_CTRL;
  wire       [1:0]    execute_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_execute_ALU_BITWISE_CTRL;
  reg                 _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
  reg                 _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
  wire                writeBack_CfuPlugin_CFU_IN_FLIGHT;
  wire       [0:0]    execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire                writeBack_HAS_SIDE_EFFECT;
  wire                memory_HAS_SIDE_EFFECT;
  wire                execute_LEGAL_INSTRUCTION;
  reg                 execute_CfuPlugin_CFU_ENABLE;
  reg                 _zz_memory_to_writeBack_FPU_FORKED;
  reg                 _zz_execute_to_memory_FPU_FORKED;
  reg                 _zz_decode_to_execute_FPU_FORKED;
  wire       [3:0]    writeBack_FPU_OPCODE;
  wire       [3:0]    _zz_writeBack_FPU_OPCODE;
  wire       [31:0]   writeBack_RS1;
  wire       [63:0]   _zz_writeBack_FpuPlugin_commit_payload_value;
  wire                writeBack_FPU_COMMIT_LOAD;
  reg                 DBusBypass0_cond;
  wire                writeBack_FPU_COMMIT;
  wire                writeBack_FPU_RSP;
  wire                writeBack_FPU_FORKED;
  wire       [0:0]    decode_FPU_FORMAT;
  wire       [0:0]    _zz_decode_FPU_FORMAT;
  wire       [1:0]    decode_FPU_ARG;
  wire       [3:0]    decode_FPU_OPCODE;
  wire       [3:0]    _zz_decode_FPU_OPCODE;
  reg                 decode_FPU_ENABLE;
  wire                execute_IS_RS1_SIGNED;
  wire                execute_IS_DIV;
  wire                execute_IS_RS2_SIGNED;
  wire                memory_IS_DIV;
  wire                writeBack_IS_MUL;
  wire       [33:0]   writeBack_MUL_HH;
  wire       [51:0]   writeBack_MUL_LOW;
  wire       [33:0]   memory_MUL_HL;
  wire       [33:0]   memory_MUL_LH;
  wire       [31:0]   memory_MUL_LL;
  wire                execute_IS_MUL;
  wire       [31:0]   memory_BRANCH_CALC;
  wire                memory_BRANCH_DO;
  wire       [31:0]   execute_PC;
  wire       [1:0]    execute_BRANCH_CTRL;
  wire       [1:0]    _zz_execute_BRANCH_CTRL;
  wire                execute_SRC_LESS;
  wire                execute_CSR_READ_OPCODE;
  wire                execute_CSR_WRITE_OPCODE;
  wire                execute_IS_CSR;
  wire       [1:0]    memory_ENV_CTRL;
  wire       [1:0]    _zz_memory_ENV_CTRL;
  wire       [1:0]    execute_ENV_CTRL;
  wire       [1:0]    _zz_execute_ENV_CTRL;
  wire       [1:0]    writeBack_ENV_CTRL;
  wire       [1:0]    _zz_writeBack_ENV_CTRL;
  reg                 CsrPlugin_running_aheadValue;
  wire                decode_RS2_USE;
  wire                decode_RS1_USE;
  reg        [31:0]   _zz_decode_RS2;
  wire                execute_REGFILE_WRITE_VALID;
  wire                execute_BYPASSABLE_EXECUTE_STAGE;
  reg        [31:0]   _zz_decode_RS2_1;
  wire                memory_REGFILE_WRITE_VALID;
  wire                memory_BYPASSABLE_MEMORY_STAGE;
  wire                writeBack_REGFILE_WRITE_VALID;
  reg        [31:0]   decode_RS2;
  reg        [31:0]   decode_RS1;
  wire                execute_SRC_LESS_UNSIGNED;
  wire                execute_SRC2_FORCE_ZERO;
  wire       [31:0]   execute_SRC2;
  wire                execute_SRC_USE_SUB_LESS;
  wire       [31:0]   execute_SRC1;
  wire       [31:0]   _zz_decode_to_execute_PC;
  wire       [31:0]   _zz_decode_to_execute_RS2;
  wire       [1:0]    decode_SRC2_CTRL;
  wire       [1:0]    _zz_decode_SRC2_CTRL;
  wire       [31:0]   _zz_decode_to_execute_RS1;
  wire       [1:0]    decode_SRC1_CTRL;
  wire       [1:0]    _zz_decode_SRC1_CTRL;
  wire                decode_SRC_USE_SUB_LESS;
  wire                decode_SRC_ADD_ZERO;
  wire       [31:0]   _zz_lastStageRegFileWrite_payload_address;
  wire                _zz_lastStageRegFileWrite_valid;
  reg                 _zz_1;
  wire       [31:0]   decode_INSTRUCTION_ANTICIPATED;
  reg                 decode_REGFILE_WRITE_VALID;
  reg                 decode_LEGAL_INSTRUCTION;
  wire       [1:0]    _zz_decode_SHIFT_CTRL_1;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL_1;
  wire       [0:0]    _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1;
  wire       [0:0]    _zz_decode_FPU_FORMAT_1;
  wire       [3:0]    _zz_decode_FPU_OPCODE_1;
  wire                _zz_decode_FPU_ENABLE;
  wire       [1:0]    _zz_decode_BRANCH_CTRL_1;
  wire       [1:0]    _zz_decode_ENV_CTRL_1;
  wire       [1:0]    _zz_decode_SRC2_CTRL_1;
  wire       [1:0]    _zz_decode_ALU_CTRL_1;
  wire       [1:0]    _zz_decode_SRC1_CTRL_1;
  reg        [31:0]   _zz_decode_RS2_2;
  wire                writeBack_MEMORY_WR;
  wire                writeBack_MEMORY_FENCE;
  wire                writeBack_MEMORY_AMO;
  wire                writeBack_MEMORY_LRSC;
  wire       [31:0]   writeBack_MEMORY_STORE_DATA_RF;
  wire       [31:0]   writeBack_REGFILE_WRITE_DATA;
  wire                writeBack_MEMORY_ENABLE;
  wire       [31:0]   memory_PC;
  wire       [31:0]   memory_MEMORY_STORE_DATA_RF;
  wire       [31:0]   memory_REGFILE_WRITE_DATA;
  wire       [31:0]   memory_INSTRUCTION;
  wire                memory_MEMORY_WR;
  wire                memory_MEMORY_ENABLE;
  wire                execute_MEMORY_FENCE_WR;
  wire       [31:0]   memory_MEMORY_VIRTUAL_ADDRESS;
  wire                execute_MEMORY_AMO;
  wire                execute_MEMORY_LRSC;
  wire                execute_MEMORY_FORCE_CONSTISTENCY;
  (* keep , syn_keep *) wire       [31:0]   execute_RS1 /* synthesis syn_keep = 1 */ ;
  wire                execute_MEMORY_MANAGMENT;
  (* keep , syn_keep *) wire       [31:0]   execute_RS2 /* synthesis syn_keep = 1 */ ;
  wire                execute_MEMORY_WR;
  wire       [31:0]   execute_SRC_ADD;
  wire                execute_MEMORY_ENABLE;
  wire       [31:0]   execute_INSTRUCTION;
  wire                decode_MEMORY_AMO;
  wire                decode_MEMORY_LRSC;
  reg                 _zz_decode_MEMORY_FORCE_CONSTISTENCY;
  wire                decode_MEMORY_ENABLE;
  wire                decode_FLUSH_ALL;
  reg                 IBusCachedPlugin_rsp_issueDetected_4;
  reg                 IBusCachedPlugin_rsp_issueDetected_3;
  reg                 IBusCachedPlugin_rsp_issueDetected_2;
  reg                 IBusCachedPlugin_rsp_issueDetected_1;
  reg        [31:0]   _zz_memory_to_writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   decode_PC;
  wire       [31:0]   decode_INSTRUCTION;
  wire                decode_IS_RVC;
  wire       [31:0]   writeBack_PC;
  wire       [31:0]   writeBack_INSTRUCTION;
  reg                 decode_arbitration_haltItself;
  reg                 decode_arbitration_haltByOther;
  reg                 decode_arbitration_removeIt;
  wire                decode_arbitration_flushIt;
  reg                 decode_arbitration_flushNext;
  reg                 decode_arbitration_isValid;
  wire                decode_arbitration_isStuck;
  wire                decode_arbitration_isStuckByOthers;
  wire                decode_arbitration_isFlushed;
  wire                decode_arbitration_isMoving;
  wire                decode_arbitration_isFiring;
  reg                 execute_arbitration_haltItself;
  reg                 execute_arbitration_haltByOther;
  reg                 execute_arbitration_removeIt;
  wire                execute_arbitration_flushIt;
  reg                 execute_arbitration_flushNext;
  reg                 execute_arbitration_isValid;
  wire                execute_arbitration_isStuck;
  wire                execute_arbitration_isStuckByOthers;
  wire                execute_arbitration_isFlushed;
  wire                execute_arbitration_isMoving;
  wire                execute_arbitration_isFiring;
  reg                 memory_arbitration_haltItself;
  reg                 memory_arbitration_haltByOther;
  reg                 memory_arbitration_removeIt;
  wire                memory_arbitration_flushIt;
  reg                 memory_arbitration_flushNext;
  reg                 memory_arbitration_isValid;
  wire                memory_arbitration_isStuck;
  wire                memory_arbitration_isStuckByOthers;
  wire                memory_arbitration_isFlushed;
  wire                memory_arbitration_isMoving;
  wire                memory_arbitration_isFiring;
  reg                 writeBack_arbitration_haltItself;
  reg                 writeBack_arbitration_haltByOther;
  reg                 writeBack_arbitration_removeIt;
  reg                 writeBack_arbitration_flushIt;
  reg                 writeBack_arbitration_flushNext;
  reg                 writeBack_arbitration_isValid;
  wire                writeBack_arbitration_isStuck;
  wire                writeBack_arbitration_isStuckByOthers;
  wire                writeBack_arbitration_isFlushed;
  wire                writeBack_arbitration_isMoving;
  wire                writeBack_arbitration_isFiring;
  wire       [31:0]   lastStageInstruction /* verilator public */ ;
  wire       [31:0]   lastStagePc /* verilator public */ ;
  wire                lastStageIsValid /* verilator public */ ;
  wire                lastStageIsFiring /* verilator public */ ;
  reg                 IBusCachedPlugin_fetcherHalt;
  wire                IBusCachedPlugin_forceNoDecodeCond;
  reg                 IBusCachedPlugin_incomingInstruction;
  wire                IBusCachedPlugin_pcValids_0;
  wire                IBusCachedPlugin_pcValids_1;
  wire                IBusCachedPlugin_pcValids_2;
  wire                IBusCachedPlugin_pcValids_3;
  reg                 IBusCachedPlugin_decodeExceptionPort_valid;
  reg        [3:0]    IBusCachedPlugin_decodeExceptionPort_payload_code;
  wire       [31:0]   IBusCachedPlugin_decodeExceptionPort_payload_badAddr;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   IBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                IBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                IBusCachedPlugin_mmuBus_rsp_isPaging;
  wire                IBusCachedPlugin_mmuBus_rsp_allowRead;
  wire                IBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire                IBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                IBusCachedPlugin_mmuBus_rsp_exception;
  wire                IBusCachedPlugin_mmuBus_rsp_refilling;
  wire                IBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                IBusCachedPlugin_mmuBus_end;
  wire                IBusCachedPlugin_mmuBus_busy;
  wire                DBusCachedPlugin_trigger_valid;
  wire                DBusCachedPlugin_trigger_load;
  wire                DBusCachedPlugin_trigger_store;
  wire       [31:0]   DBusCachedPlugin_trigger_virtual;
  wire       [31:0]   DBusCachedPlugin_trigger_writeData;
  wire       [31:0]   DBusCachedPlugin_trigger_readData;
  wire                DBusCachedPlugin_trigger_readDataValid;
  wire       [1:0]    DBusCachedPlugin_trigger_size;
  wire       [31:0]   DBusCachedPlugin_trigger_dpc;
  wire                DBusCachedPlugin_trigger_hit;
  wire                DBusCachedPlugin_trigger_hitBefore;
  wire                DBusCachedPlugin_writesPending;
  wire                DBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                DBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   DBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   DBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                DBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                DBusCachedPlugin_mmuBus_rsp_isPaging;
  wire                DBusCachedPlugin_mmuBus_rsp_allowRead;
  wire                DBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire                DBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                DBusCachedPlugin_mmuBus_rsp_exception;
  wire                DBusCachedPlugin_mmuBus_rsp_refilling;
  wire                DBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                DBusCachedPlugin_mmuBus_end;
  wire                DBusCachedPlugin_mmuBus_busy;
  reg                 DBusCachedPlugin_redoBranch_valid;
  wire       [31:0]   DBusCachedPlugin_redoBranch_payload;
  reg                 DBusCachedPlugin_exceptionBus_valid;
  reg        [3:0]    DBusCachedPlugin_exceptionBus_payload_code;
  wire       [31:0]   DBusCachedPlugin_exceptionBus_payload_badAddr;
  wire                decodeExceptionPort_valid;
  wire       [3:0]    decodeExceptionPort_payload_code;
  wire       [31:0]   decodeExceptionPort_payload_badAddr;
  wire       [31:0]   CsrPlugin_csrMapping_readDataSignal;
  wire       [31:0]   CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   CsrPlugin_csrMapping_writeDataSignal;
  reg                 CsrPlugin_csrMapping_allowCsrSignal;
  wire                CsrPlugin_csrMapping_hazardFree;
  reg                 CsrPlugin_csrMapping_doForceFailCsr;
  wire                CsrPlugin_inWfi /* verilator public */ ;
  reg                 CsrPlugin_thirdPartyWake;
  reg                 CsrPlugin_jumpInterface_valid;
  reg        [31:0]   CsrPlugin_jumpInterface_payload;
  wire                CsrPlugin_exceptionPendings_0;
  wire                CsrPlugin_exceptionPendings_1;
  wire                CsrPlugin_exceptionPendings_2;
  wire                CsrPlugin_exceptionPendings_3;
  wire                contextSwitching;
  reg        [1:0]    CsrPlugin_privilege;
  wire                CsrPlugin_forceMachineWire;
  reg                 CsrPlugin_selfException_valid;
  reg        [3:0]    CsrPlugin_selfException_payload_code;
  wire       [31:0]   CsrPlugin_selfException_payload_badAddr;
  reg                 CsrPlugin_allowInterrupts;
  wire                CsrPlugin_allowException;
  wire                CsrPlugin_allowEbreakException;
  reg                 CsrPlugin_xretAwayFromMachine;
  wire                fpuAccess_start;
  wire       [4:0]    fpuAccess_regId;
  wire       [2:0]    fpuAccess_size;
  wire                fpuAccess_write;
  wire       [63:0]   fpuAccess_writeData;
  reg        [31:0]   fpuAccess_readData;
  reg                 fpuAccess_readDataValid;
  reg        [0:0]    fpuAccess_readDataChunk;
  reg                 fpuAccess_done;
  wire                CsrPlugin_injectionPort_valid;
  reg                 CsrPlugin_injectionPort_ready;
  wire       [31:0]   CsrPlugin_injectionPort_payload;
  wire                debugMode;
  wire                BranchPlugin_jumpInterface_valid;
  wire       [31:0]   BranchPlugin_jumpInterface_payload;
  reg                 BranchPlugin_inDebugNoFetchFlag;
  wire                IBusCachedPlugin_externalFlush;
  wire                IBusCachedPlugin_jump_pcLoad_valid;
  wire       [31:0]   IBusCachedPlugin_jump_pcLoad_payload;
  wire       [2:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload;
  wire       [2:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  wire                _zz_IBusCachedPlugin_jump_pcLoad_payload_2;
  wire                _zz_IBusCachedPlugin_jump_pcLoad_payload_3;
  wire                IBusCachedPlugin_fetchPc_output_valid;
  wire                IBusCachedPlugin_fetchPc_output_ready;
  wire       [31:0]   IBusCachedPlugin_fetchPc_output_payload;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pcReg /* verilator public */ ;
  reg                 IBusCachedPlugin_fetchPc_correction;
  reg                 IBusCachedPlugin_fetchPc_correctionReg;
  wire                IBusCachedPlugin_fetchPc_output_fire;
  wire                IBusCachedPlugin_fetchPc_corrected;
  reg                 IBusCachedPlugin_fetchPc_pcRegPropagate;
  reg                 IBusCachedPlugin_fetchPc_booted;
  reg                 IBusCachedPlugin_fetchPc_inc;
  wire                when_Fetcher_l133;
  wire                when_Fetcher_l133_1;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pc;
  wire                IBusCachedPlugin_fetchPc_redo_valid;
  reg        [31:0]   IBusCachedPlugin_fetchPc_redo_payload;
  reg                 IBusCachedPlugin_fetchPc_flushed;
  wire                when_Fetcher_l160;
  reg                 IBusCachedPlugin_decodePc_flushed;
  reg        [31:0]   IBusCachedPlugin_decodePc_pcReg /* verilator public */ ;
  wire       [31:0]   IBusCachedPlugin_decodePc_pcPlus;
  reg                 IBusCachedPlugin_decodePc_injectedDecode;
  wire                when_Fetcher_l182;
  wire                when_Fetcher_l194;
  reg                 IBusCachedPlugin_iBusRsp_redoFetch;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_0_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_1_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_2_halt;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire                IBusCachedPlugin_iBusRsp_flush;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  reg        [31:0]   _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 IBusCachedPlugin_iBusRsp_readyForError;
  wire                IBusCachedPlugin_iBusRsp_output_valid;
  wire                IBusCachedPlugin_iBusRsp_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_pc;
  wire                IBusCachedPlugin_iBusRsp_output_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  wire                IBusCachedPlugin_iBusRsp_output_payload_isRvc;
  wire                when_Fetcher_l242;
  wire                IBusCachedPlugin_decompressor_input_valid;
  wire                IBusCachedPlugin_decompressor_input_ready;
  wire       [31:0]   IBusCachedPlugin_decompressor_input_payload_pc;
  wire                IBusCachedPlugin_decompressor_input_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_decompressor_input_payload_rsp_inst;
  wire                IBusCachedPlugin_decompressor_input_payload_isRvc;
  wire                IBusCachedPlugin_decompressor_output_valid;
  wire                IBusCachedPlugin_decompressor_output_ready;
  wire       [31:0]   IBusCachedPlugin_decompressor_output_payload_pc;
  wire                IBusCachedPlugin_decompressor_output_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_decompressor_output_payload_rsp_inst;
  wire                IBusCachedPlugin_decompressor_output_payload_isRvc;
  wire                IBusCachedPlugin_decompressor_flushNext;
  wire                IBusCachedPlugin_decompressor_consumeCurrent;
  reg                 IBusCachedPlugin_decompressor_bufferValid;
  reg        [15:0]   IBusCachedPlugin_decompressor_bufferData;
  wire                IBusCachedPlugin_decompressor_isInputLowRvc;
  wire                IBusCachedPlugin_decompressor_isInputHighRvc;
  reg                 IBusCachedPlugin_decompressor_throw2BytesReg;
  wire                IBusCachedPlugin_decompressor_throw2Bytes;
  wire                IBusCachedPlugin_decompressor_unaligned;
  reg                 IBusCachedPlugin_decompressor_bufferValidLatch;
  reg                 IBusCachedPlugin_decompressor_throw2BytesLatch;
  wire                IBusCachedPlugin_decompressor_bufferValidPatched;
  wire                IBusCachedPlugin_decompressor_throw2BytesPatched;
  wire       [31:0]   IBusCachedPlugin_decompressor_raw;
  wire                IBusCachedPlugin_decompressor_isRvc;
  wire       [15:0]   _zz_IBusCachedPlugin_decompressor_decompressed;
  reg        [31:0]   IBusCachedPlugin_decompressor_decompressed;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_1;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_2;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_3;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_4;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_5;
  reg        [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_6;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_7;
  reg        [9:0]    _zz_IBusCachedPlugin_decompressor_decompressed_8;
  wire       [20:0]   _zz_IBusCachedPlugin_decompressor_decompressed_9;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_10;
  reg        [14:0]   _zz_IBusCachedPlugin_decompressor_decompressed_11;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_12;
  reg        [2:0]    _zz_IBusCachedPlugin_decompressor_decompressed_13;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_14;
  reg        [9:0]    _zz_IBusCachedPlugin_decompressor_decompressed_15;
  wire       [20:0]   _zz_IBusCachedPlugin_decompressor_decompressed_16;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_17;
  reg        [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_18;
  wire       [12:0]   _zz_IBusCachedPlugin_decompressor_decompressed_19;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_20;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_21;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_22;
  wire       [4:0]    switch_Misc_l44;
  wire                when_Misc_l47;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_23;
  wire       [1:0]    switch_Misc_l241;
  wire       [1:0]    switch_Misc_l241_1;
  reg        [2:0]    _zz_IBusCachedPlugin_decompressor_decompressed_24;
  reg        [2:0]    _zz_IBusCachedPlugin_decompressor_decompressed_25;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_26;
  reg        [6:0]    _zz_IBusCachedPlugin_decompressor_decompressed_27;
  wire                IBusCachedPlugin_decompressor_output_fire;
  wire                IBusCachedPlugin_decompressor_bufferFill;
  wire                when_Fetcher_l285;
  wire                when_Fetcher_l288;
  wire                when_Fetcher_l293;
  wire                IBusCachedPlugin_injector_decodeInput_valid;
  wire                IBusCachedPlugin_injector_decodeInput_ready;
  wire       [31:0]   IBusCachedPlugin_injector_decodeInput_payload_pc;
  wire                IBusCachedPlugin_injector_decodeInput_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  wire                IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  reg                 _zz_IBusCachedPlugin_injector_decodeInput_valid;
  reg        [31:0]   _zz_IBusCachedPlugin_injector_decodeInput_payload_pc;
  reg                 _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_error;
  reg        [31:0]   _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  reg                 _zz_IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_0;
  wire                when_Fetcher_l331;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_1;
  wire                when_Fetcher_l331_1;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_2;
  wire                when_Fetcher_l331_2;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_3;
  wire                when_Fetcher_l331_3;
  reg        [31:0]   IBusCachedPlugin_injector_formal_rawInDecode;
  reg        [31:0]   IBusCachedPlugin_rspCounter;
  wire                IBusCachedPlugin_s0_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s1_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s2_tightlyCoupledHit;
  wire                IBusCachedPlugin_rsp_iBusRspOutputHalt;
  wire                IBusCachedPlugin_rsp_issueDetected;
  reg                 IBusCachedPlugin_rsp_redoFetch;
  wire                when_IBusCachedPlugin_l245;
  wire                when_IBusCachedPlugin_l250;
  wire                when_IBusCachedPlugin_l256;
  wire                when_IBusCachedPlugin_l262;
  wire                when_IBusCachedPlugin_l273;
  wire                dataCache_2_io_mem_cmd_s2mPipe_valid;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_ready;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_wr;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_uncached;
  wire       [31:0]   dataCache_2_io_mem_cmd_s2mPipe_payload_address;
  wire       [63:0]   dataCache_2_io_mem_cmd_s2mPipe_payload_data;
  wire       [7:0]    dataCache_2_io_mem_cmd_s2mPipe_payload_mask;
  wire       [2:0]    dataCache_2_io_mem_cmd_s2mPipe_payload_size;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_exclusive;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_last;
  reg                 dataCache_2_io_mem_cmd_rValidN;
  reg                 dataCache_2_io_mem_cmd_rData_wr;
  reg                 dataCache_2_io_mem_cmd_rData_uncached;
  reg        [31:0]   dataCache_2_io_mem_cmd_rData_address;
  reg        [63:0]   dataCache_2_io_mem_cmd_rData_data;
  reg        [7:0]    dataCache_2_io_mem_cmd_rData_mask;
  reg        [2:0]    dataCache_2_io_mem_cmd_rData_size;
  reg                 dataCache_2_io_mem_cmd_rData_exclusive;
  reg                 dataCache_2_io_mem_cmd_rData_last;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_ready;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_wr;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached;
  wire       [31:0]   dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_address;
  wire       [63:0]   dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_data;
  wire       [7:0]    dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_mask;
  wire       [2:0]    dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_size;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_exclusive;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_last;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rValid;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_wr;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_uncached;
  reg        [31:0]   dataCache_2_io_mem_cmd_s2mPipe_rData_address;
  reg        [63:0]   dataCache_2_io_mem_cmd_s2mPipe_rData_data;
  reg        [7:0]    dataCache_2_io_mem_cmd_s2mPipe_rData_mask;
  reg        [2:0]    dataCache_2_io_mem_cmd_s2mPipe_rData_size;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_exclusive;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_last;
  wire                when_Stream_l375;
  reg                 dBus_rsp_valid_regNext;
  reg                 dBus_rsp_payload_exclusive_regNext;
  reg                 dBus_rsp_payload_error_regNext;
  reg                 dBus_rsp_payload_last_regNext;
  reg        [3:0]    dBus_rsp_payload_aggregated_regNext;
  wire                when_DBusCachedPlugin_l334;
  reg        [63:0]   dBus_rsp_payload_data_regNextWhen;
  reg        [31:0]   DBusCachedPlugin_rspCounter;
  wire                when_DBusCachedPlugin_l356;
  wire                when_DBusCachedPlugin_l364;
  wire       [1:0]    execute_DBusCachedPlugin_size;
  reg        [31:0]   _zz_execute_MEMORY_STORE_DATA_RF;
  wire                dataCache_2_io_cpu_flush_isStall;
  wire                when_DBusCachedPlugin_l398;
  wire                when_DBusCachedPlugin_l414;
  wire                when_DBusCachedPlugin_l427;
  wire                when_DBusCachedPlugin_l476;
  wire       [11:0]   _zz_io_cpu_writeBack_fence_SW;
  reg                 writeBack_DBusCachedPlugin_fence_aquire;
  wire                when_DBusCachedPlugin_l518;
  wire                when_DBusCachedPlugin_l531;
  wire                when_DBusCachedPlugin_l535;
  wire                when_DBusCachedPlugin_l552;
  wire                when_DBusCachedPlugin_l572;
  wire       [63:0]   writeBack_DBusCachedPlugin_rspData;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_0;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_1;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_2;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_3;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_4;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_5;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_6;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_7;
  reg        [63:0]   writeBack_DBusCachedPlugin_rspShifted;
  reg        [31:0]   writeBack_DBusCachedPlugin_rspRf;
  wire                when_DBusCachedPlugin_l589;
  wire       [1:0]    switch_Misc_l241_2;
  wire                _zz_writeBack_DBusCachedPlugin_rspFormated;
  reg        [31:0]   _zz_writeBack_DBusCachedPlugin_rspFormated_1;
  wire                _zz_writeBack_DBusCachedPlugin_rspFormated_2;
  reg        [31:0]   _zz_writeBack_DBusCachedPlugin_rspFormated_3;
  reg        [31:0]   writeBack_DBusCachedPlugin_rspFormated;
  wire                when_DBusCachedPlugin_l599;
  wire       [47:0]   _zz_decode_CfuPlugin_CFU_ENABLE;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_1;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_2;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_3;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_4;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_5;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_6;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_7;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_8;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_9;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_10;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_11;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_12;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_13;
  wire       [1:0]    _zz_decode_SRC1_CTRL_2;
  wire       [1:0]    _zz_decode_ALU_CTRL_2;
  wire       [1:0]    _zz_decode_SRC2_CTRL_2;
  wire       [1:0]    _zz_decode_ENV_CTRL_2;
  wire       [1:0]    _zz_decode_BRANCH_CTRL_2;
  wire       [3:0]    _zz_decode_FPU_OPCODE_2;
  wire       [0:0]    _zz_decode_FPU_FORMAT_2;
  wire       [0:0]    _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL_2;
  wire       [1:0]    _zz_decode_SHIFT_CTRL_2;
  wire                when_RegFilePlugin_l63;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress1;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress2;
  wire       [31:0]   decode_RegFilePlugin_rs1Data;
  wire       [31:0]   decode_RegFilePlugin_rs2Data;
  reg                 lastStageRegFileWrite_valid /* verilator public */ ;
  reg        [4:0]    lastStageRegFileWrite_payload_address /* verilator public */ ;
  reg        [31:0]   lastStageRegFileWrite_payload_data /* verilator public */ ;
  reg                 _zz_5;
  reg        [31:0]   _zz_decode_SRC1;
  wire                _zz_decode_SRC2;
  reg        [19:0]   _zz_decode_SRC2_1;
  wire                _zz_decode_SRC2_2;
  reg        [19:0]   _zz_decode_SRC2_3;
  reg        [31:0]   _zz_decode_SRC2_4;
  reg        [31:0]   execute_SrcPlugin_addSub;
  wire                execute_SrcPlugin_less;
  reg                 HazardSimplePlugin_src0Hazard;
  reg                 HazardSimplePlugin_src1Hazard;
  wire                HazardSimplePlugin_writeBackWrites_valid;
  wire       [4:0]    HazardSimplePlugin_writeBackWrites_payload_address;
  wire       [31:0]   HazardSimplePlugin_writeBackWrites_payload_data;
  reg                 HazardSimplePlugin_writeBackBuffer_valid;
  reg        [4:0]    HazardSimplePlugin_writeBackBuffer_payload_address;
  reg        [31:0]   HazardSimplePlugin_writeBackBuffer_payload_data;
  wire                HazardSimplePlugin_addr0Match;
  wire                HazardSimplePlugin_addr1Match;
  wire                when_HazardSimplePlugin_l47;
  wire                when_HazardSimplePlugin_l48;
  wire                when_HazardSimplePlugin_l51;
  wire                when_HazardSimplePlugin_l45;
  wire                when_HazardSimplePlugin_l57;
  wire                when_HazardSimplePlugin_l58;
  wire                when_HazardSimplePlugin_l48_1;
  wire                when_HazardSimplePlugin_l51_1;
  wire                when_HazardSimplePlugin_l45_1;
  wire                when_HazardSimplePlugin_l57_1;
  wire                when_HazardSimplePlugin_l58_1;
  wire                when_HazardSimplePlugin_l48_2;
  wire                when_HazardSimplePlugin_l51_2;
  wire                when_HazardSimplePlugin_l45_2;
  wire                when_HazardSimplePlugin_l57_2;
  wire                when_HazardSimplePlugin_l58_2;
  wire                when_HazardSimplePlugin_l105;
  wire                when_HazardSimplePlugin_l108;
  wire                when_HazardSimplePlugin_l113;
  reg                 when_CsrPlugin_l836;
  reg        [1:0]    _zz_CsrPlugin_privilege;
  reg                 CsrPlugin_running;
  wire                when_CsrPlugin_l729;
  reg                 CsrPlugin_reseting;
  reg                 _zz_debugBus_haveReset;
  reg                 CsrPlugin_running_aheadValue_regNext;
  wire                CsrPlugin_enterHalt;
  reg                 CsrPlugin_doHalt;
  wire                when_CsrPlugin_l747;
  wire                CsrPlugin_forceResume;
  reg                 _zz_CsrPlugin_doResume;
  wire                CsrPlugin_doResume;
  reg                 CsrPlugin_timeout_state;
  reg                 CsrPlugin_timeout_stateRise;
  wire                CsrPlugin_timeout_counter_willIncrement;
  reg                 CsrPlugin_timeout_counter_willClear;
  reg        [2:0]    CsrPlugin_timeout_counter_valueNext;
  reg        [2:0]    CsrPlugin_timeout_counter_value;
  wire                CsrPlugin_timeout_counter_willOverflowIfInc;
  wire                CsrPlugin_timeout_counter_willOverflow;
  wire                when_CsrPlugin_l753;
  reg                 _zz_debugBus_hartToDm_valid;
  reg        [31:0]   CsrPlugin_dataCsrw_value_0;
  reg        [31:0]   CsrPlugin_dataCsrw_value_1;
  wire                when_CsrPlugin_l768;
  wire       [1:0]    _zz_6;
  wire                CsrPlugin_inject_cmd_valid;
  wire       [1:0]    CsrPlugin_inject_cmd_payload_op;
  wire       [4:0]    CsrPlugin_inject_cmd_payload_address;
  wire       [31:0]   CsrPlugin_inject_cmd_payload_data;
  wire       [2:0]    CsrPlugin_inject_cmd_payload_size;
  wire                CsrPlugin_inject_cmd_toStream_valid;
  reg                 CsrPlugin_inject_cmd_toStream_ready;
  wire       [1:0]    CsrPlugin_inject_cmd_toStream_payload_op;
  wire       [4:0]    CsrPlugin_inject_cmd_toStream_payload_address;
  wire       [31:0]   CsrPlugin_inject_cmd_toStream_payload_data;
  wire       [2:0]    CsrPlugin_inject_cmd_toStream_payload_size;
  wire                CsrPlugin_inject_buffer_valid;
  reg                 CsrPlugin_inject_buffer_ready;
  wire       [1:0]    CsrPlugin_inject_buffer_payload_op;
  wire       [4:0]    CsrPlugin_inject_buffer_payload_address;
  wire       [31:0]   CsrPlugin_inject_buffer_payload_data;
  wire       [2:0]    CsrPlugin_inject_buffer_payload_size;
  reg                 CsrPlugin_inject_cmd_toStream_rValid;
  reg        [1:0]    CsrPlugin_inject_cmd_toStream_rData_op;
  reg        [4:0]    CsrPlugin_inject_cmd_toStream_rData_address;
  reg        [31:0]   CsrPlugin_inject_cmd_toStream_rData_data;
  reg        [2:0]    CsrPlugin_inject_cmd_toStream_rData_size;
  wire                when_Stream_l375_1;
  wire                CsrPlugin_injectionPort_fire;
  reg                 CsrPlugin_inject_pending;
  wire                when_CsrPlugin_l804;
  wire                when_CsrPlugin_l804_1;
  reg        [31:0]   CsrPlugin_dpc;
  reg        [1:0]    CsrPlugin_dcsr_prv;
  reg                 CsrPlugin_dcsr_step;
  wire                CsrPlugin_dcsr_nmip;
  wire                CsrPlugin_dcsr_mprven;
  reg        [2:0]    CsrPlugin_dcsr_cause;
  reg                 CsrPlugin_dcsr_stoptime;
  reg                 CsrPlugin_dcsr_stopcount;
  reg                 CsrPlugin_dcsr_stepie;
  reg                 CsrPlugin_dcsr_ebreakm;
  wire       [3:0]    CsrPlugin_dcsr_xdebugver;
  wire                CsrPlugin_dcsr_stepLogic_wantExit;
  reg                 CsrPlugin_dcsr_stepLogic_wantStart;
  wire                CsrPlugin_dcsr_stepLogic_wantKill;
  reg        [1:0]    CsrPlugin_dcsr_stepLogic_stateReg;
  reg        [1:0]    CsrPlugin_dcsr_stepLogic_stateNext;
  wire                when_CsrPlugin_l830;
  wire                when_CsrPlugin_l848;
  wire                when_CsrPlugin_l880;
  wire       [1:0]    CsrPlugin_misa_base;
  wire       [25:0]   CsrPlugin_misa_extensions;
  reg        [1:0]    CsrPlugin_mtvec_mode;
  reg        [29:0]   CsrPlugin_mtvec_base;
  reg        [31:0]   CsrPlugin_mepc;
  reg                 CsrPlugin_mstatus_MIE;
  reg                 CsrPlugin_mstatus_MPIE;
  reg        [1:0]    CsrPlugin_mstatus_MPP;
  reg                 CsrPlugin_mip_MEIP;
  reg                 CsrPlugin_mip_MTIP;
  reg                 CsrPlugin_mip_MSIP;
  reg                 CsrPlugin_mie_MEIE;
  reg                 CsrPlugin_mie_MTIE;
  reg                 CsrPlugin_mie_MSIE;
  reg        [31:0]   CsrPlugin_mscratch;
  reg                 CsrPlugin_mcause_interrupt;
  reg        [3:0]    CsrPlugin_mcause_exceptionCode;
  reg        [31:0]   CsrPlugin_mtval;
  reg        [63:0]   CsrPlugin_counters_mcycle;
  reg        [63:0]   CsrPlugin_counters_minstret;
  wire                _zz_when_CsrPlugin_l1446;
  wire                _zz_when_CsrPlugin_l1446_1;
  wire                _zz_when_CsrPlugin_l1446_2;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  reg        [3:0]    CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  reg        [31:0]   CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
  wire       [1:0]    _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  wire                _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire                when_CsrPlugin_l1403;
  wire                when_CsrPlugin_l1403_1;
  wire                when_CsrPlugin_l1403_2;
  wire                when_CsrPlugin_l1403_3;
  wire                when_CsrPlugin_l1416;
  reg                 CsrPlugin_interrupt_valid;
  reg        [3:0]    CsrPlugin_interrupt_code /* verilator public */ ;
  reg        [1:0]    CsrPlugin_interrupt_targetPrivilege;
  wire                when_CsrPlugin_l1440;
  wire                when_CsrPlugin_l1446;
  wire                when_CsrPlugin_l1446_1;
  wire                when_CsrPlugin_l1446_2;
  wire                when_CsrPlugin_l1459;
  wire                CsrPlugin_exception;
  wire                CsrPlugin_lastStageWasWfi;
  reg                 CsrPlugin_pipelineLiberator_pcValids_0;
  reg                 CsrPlugin_pipelineLiberator_pcValids_1;
  reg                 CsrPlugin_pipelineLiberator_pcValids_2;
  wire                CsrPlugin_pipelineLiberator_active;
  wire                when_CsrPlugin_l1479;
  wire                when_CsrPlugin_l1479_1;
  wire                when_CsrPlugin_l1479_2;
  wire                when_CsrPlugin_l1484;
  reg                 CsrPlugin_pipelineLiberator_done;
  wire                when_CsrPlugin_l1490;
  wire                CsrPlugin_interruptJump /* verilator public */ ;
  reg                 CsrPlugin_hadException /* verilator public */ ;
  reg        [1:0]    CsrPlugin_targetPrivilege;
  reg        [3:0]    CsrPlugin_trapCause;
  reg                 CsrPlugin_trapCauseEbreakDebug;
  wire                when_CsrPlugin_l1517;
  wire                when_CsrPlugin_l1519;
  reg        [1:0]    CsrPlugin_xtvec_mode;
  reg        [29:0]   CsrPlugin_xtvec_base;
  reg                 CsrPlugin_trapEnterDebug;
  wire                when_CsrPlugin_l1533;
  wire                when_CsrPlugin_l1534;
  wire                when_CsrPlugin_l1542;
  wire                when_CsrPlugin_l1572;
  wire                when_CsrPlugin_l1600;
  wire       [1:0]    switch_CsrPlugin_l1604;
  wire                when_CsrPlugin_l1612;
  reg                 execute_CsrPlugin_wfiWake;
  wire                when_CsrPlugin_l1671;
  wire                execute_CsrPlugin_blockedBySideEffects;
  reg                 execute_CsrPlugin_illegalAccess;
  reg                 execute_CsrPlugin_illegalInstruction;
  wire                when_CsrPlugin_l1684;
  wire                when_CsrPlugin_l1691;
  wire                when_CsrPlugin_l1692;
  wire                when_CsrPlugin_l1699;
  wire                when_CsrPlugin_l1709;
  reg                 execute_CsrPlugin_writeInstruction;
  reg                 execute_CsrPlugin_readInstruction;
  wire                execute_CsrPlugin_writeEnable;
  wire                execute_CsrPlugin_readEnable;
  wire       [31:0]   execute_CsrPlugin_readToWriteData;
  wire                switch_Misc_l241_3;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_writeDataSignal;
  wire                when_CsrPlugin_l1731;
  wire                when_CsrPlugin_l1735;
  wire       [11:0]   execute_CsrPlugin_csrAddress;
  wire                execute_BranchPlugin_eq;
  wire       [2:0]    switch_Misc_l241_4;
  reg                 _zz_execute_BRANCH_DO;
  reg                 _zz_execute_BRANCH_DO_1;
  wire       [31:0]   execute_BranchPlugin_branch_src1;
  wire                _zz_execute_BranchPlugin_branch_src2;
  reg        [10:0]   _zz_execute_BranchPlugin_branch_src2_1;
  wire                _zz_execute_BranchPlugin_branch_src2_2;
  reg        [19:0]   _zz_execute_BranchPlugin_branch_src2_3;
  wire                _zz_execute_BranchPlugin_branch_src2_4;
  reg        [18:0]   _zz_execute_BranchPlugin_branch_src2_5;
  reg        [31:0]   _zz_execute_BranchPlugin_branch_src2_6;
  wire       [31:0]   execute_BranchPlugin_branch_src2;
  wire       [31:0]   execute_BranchPlugin_branchAdder;
  reg                 execute_MulPlugin_aSigned;
  reg                 execute_MulPlugin_bSigned;
  wire       [31:0]   execute_MulPlugin_a;
  wire       [31:0]   execute_MulPlugin_b;
  reg        [0:0]    execute_MulPlugin_delayLogic_counter;
  wire                when_MulPlugin_l65;
  wire                when_MulPlugin_l70;
  wire       [1:0]    switch_MulPlugin_l87;
  wire       [15:0]   execute_MulPlugin_aULow;
  wire       [15:0]   execute_MulPlugin_bULow;
  wire       [16:0]   execute_MulPlugin_aSLow;
  wire       [16:0]   execute_MulPlugin_bSLow;
  wire       [16:0]   execute_MulPlugin_aHigh;
  wire       [16:0]   execute_MulPlugin_bHigh;
  reg        [31:0]   execute_MulPlugin_withOuputBuffer_mul_ll;
  reg        [33:0]   execute_MulPlugin_withOuputBuffer_mul_lh;
  reg        [33:0]   execute_MulPlugin_withOuputBuffer_mul_hl;
  reg        [33:0]   execute_MulPlugin_withOuputBuffer_mul_hh;
  wire       [65:0]   writeBack_MulPlugin_result;
  wire                when_MulPlugin_l147;
  wire       [1:0]    switch_MulPlugin_l148;
  reg        [32:0]   memory_MulDivIterativePlugin_rs1;
  reg        [31:0]   memory_MulDivIterativePlugin_rs2;
  reg        [64:0]   memory_MulDivIterativePlugin_accumulator;
  wire                memory_MulDivIterativePlugin_frontendOk;
  reg                 memory_MulDivIterativePlugin_div_needRevert;
  reg                 memory_MulDivIterativePlugin_div_counter_willIncrement;
  reg                 memory_MulDivIterativePlugin_div_counter_willClear;
  reg        [5:0]    memory_MulDivIterativePlugin_div_counter_valueNext;
  reg        [5:0]    memory_MulDivIterativePlugin_div_counter_value;
  wire                memory_MulDivIterativePlugin_div_counter_willOverflowIfInc;
  wire                memory_MulDivIterativePlugin_div_counter_willOverflow;
  reg                 memory_MulDivIterativePlugin_div_done;
  wire                when_MulDivIterativePlugin_l126;
  wire                when_MulDivIterativePlugin_l126_1;
  reg        [31:0]   memory_MulDivIterativePlugin_div_result;
  wire                when_MulDivIterativePlugin_l128;
  wire                when_MulDivIterativePlugin_l129;
  wire                when_MulDivIterativePlugin_l132;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted;
  wire       [32:0]   memory_MulDivIterativePlugin_div_stage_0_remainderShifted;
  wire       [32:0]   memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator;
  wire       [31:0]   memory_MulDivIterativePlugin_div_stage_0_outRemainder;
  wire       [31:0]   memory_MulDivIterativePlugin_div_stage_0_outNumerator;
  wire                when_MulDivIterativePlugin_l151;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_result;
  wire                when_MulDivIterativePlugin_l162;
  wire                _zz_memory_MulDivIterativePlugin_rs2;
  wire                _zz_memory_MulDivIterativePlugin_rs1;
  reg        [32:0]   _zz_memory_MulDivIterativePlugin_rs1_1;
  reg        [5:0]    FpuPlugin_pendings;
  wire                FpuPlugin_port_cmd_fire;
  wire                FpuPlugin_port_rsp_fire;
  wire                FpuPlugin_hasPending;
  reg                 FpuPlugin_flags_NX;
  reg                 FpuPlugin_flags_UF;
  reg                 FpuPlugin_flags_OF;
  reg                 FpuPlugin_flags_DZ;
  reg                 FpuPlugin_flags_NV;
  wire                when_FpuPlugin_l215;
  wire                when_FpuPlugin_l216;
  wire                when_FpuPlugin_l217;
  wire                when_FpuPlugin_l218;
  wire                when_FpuPlugin_l219;
  reg        [2:0]    FpuPlugin_rm;
  wire                FpuPlugin_csrActive;
  wire                when_FpuPlugin_l229;
  reg        [1:0]    FpuPlugin_fs;
  wire                FpuPlugin_sd;
  wire                when_FpuPlugin_l234;
  reg                 _zz_when_FpuPlugin_l237;
  reg                 _zz_when_FpuPlugin_l237_1;
  reg                 _zz_when_FpuPlugin_l237_2;
  wire                when_FpuPlugin_l237;
  reg                 FpuPlugin_accessFpuCsr;
  wire                when_FpuPlugin_l253;
  reg                 _zz_decode_FPU_FORKED;
  wire                decode_FpuPlugin_trap;
  reg                 decode_FpuPlugin_forked;
  wire                when_FpuPlugin_l268;
  wire                when_FpuPlugin_l268_1;
  wire                decode_FpuPlugin_hazard;
  wire                when_FpuPlugin_l272;
  wire                when_FpuPlugin_l273;
  wire                FpuPlugin_port_cmd_isStall;
  wire       [2:0]    decode_FpuPlugin_iRoundMode;
  wire       [2:0]    decode_FpuPlugin_roundMode;
  wire       [2:0]    _zz_FpuPlugin_port_cmd_payload_roundMode;
  wire       [2:0]    _zz_FpuPlugin_port_cmd_payload_roundMode_1;
  wire                writeBack_FpuPlugin_isRsp;
  wire                writeBack_FpuPlugin_isCommit;
  reg        [63:0]   writeBack_FpuPlugin_storeFormated;
  wire                when_FpuPlugin_l306;
  wire       [63:0]   DBusBypass0_value;
  wire                when_FpuPlugin_l315;
  wire                when_FpuPlugin_l318;
  wire                when_FpuPlugin_l323;
  wire                when_FpuPlugin_l325;
  wire                writeBack_FpuPlugin_commit_valid /* verilator public */ ;
  wire                writeBack_FpuPlugin_commit_ready /* verilator public */ ;
  wire       [3:0]    writeBack_FpuPlugin_commit_payload_opcode /* verilator public */ ;
  wire       [4:0]    writeBack_FpuPlugin_commit_payload_rd /* verilator public */ ;
  wire                writeBack_FpuPlugin_commit_payload_write /* verilator public */ ;
  reg        [63:0]   writeBack_FpuPlugin_commit_payload_value /* verilator public */ ;
  wire                when_FpuPlugin_l339;
  wire                writeBack_FpuPlugin_commit_s2mPipe_valid;
  wire                writeBack_FpuPlugin_commit_s2mPipe_ready;
  wire       [3:0]    writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
  wire       [4:0]    writeBack_FpuPlugin_commit_s2mPipe_payload_rd;
  wire                writeBack_FpuPlugin_commit_s2mPipe_payload_write;
  wire       [63:0]   writeBack_FpuPlugin_commit_s2mPipe_payload_value;
  reg                 writeBack_FpuPlugin_commit_rValidN;
  reg        [3:0]    writeBack_FpuPlugin_commit_rData_opcode;
  reg        [4:0]    writeBack_FpuPlugin_commit_rData_rd;
  reg                 writeBack_FpuPlugin_commit_rData_write;
  reg        [63:0]   writeBack_FpuPlugin_commit_rData_value;
  wire       [3:0]    _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
  wire                FpuPlugin_wantExit;
  reg                 FpuPlugin_wantStart;
  wire                FpuPlugin_wantKill;
  wire                when_FpuPlugin_l350;
  wire                when_CfuPlugin_l192;
  wire                execute_CfuPlugin_hazard;
  wire                execute_CfuPlugin_scheduleWish;
  wire                execute_CfuPlugin_schedule;
  wire                when_CfuPlugin_l196;
  reg                 execute_CfuPlugin_hold;
  reg                 execute_CfuPlugin_fired;
  wire                CfuPlugin_bus_cmd_fire;
  wire                when_CfuPlugin_l199;
  wire                when_CfuPlugin_l203;
  wire       [9:0]    execute_CfuPlugin_functionsIds_0;
  wire                _zz_CfuPlugin_bus_cmd_payload_inputs_1;
  reg        [23:0]   _zz_CfuPlugin_bus_cmd_payload_inputs_1_1;
  reg        [31:0]   _zz_CfuPlugin_bus_cmd_payload_inputs_1_2;
  wire                writeBack_CfuPlugin_rsp_valid;
  reg                 writeBack_CfuPlugin_rsp_ready;
  wire       [31:0]   writeBack_CfuPlugin_rsp_payload_outputs_0;
  reg                 CfuPlugin_bus_rsp_rValidN;
  reg        [31:0]   CfuPlugin_bus_rsp_rData_outputs_0;
  wire                when_CfuPlugin_l239;
  reg        [31:0]   _zz_decode_RS2_3;
  wire                when_Pipeline_l124;
  reg        [31:0]   decode_to_execute_PC;
  wire                when_Pipeline_l124_1;
  reg        [31:0]   execute_to_memory_PC;
  wire                when_Pipeline_l124_2;
  reg        [31:0]   memory_to_writeBack_PC;
  wire                when_Pipeline_l124_3;
  reg        [31:0]   decode_to_execute_INSTRUCTION;
  wire                when_Pipeline_l124_4;
  reg        [31:0]   execute_to_memory_INSTRUCTION;
  wire                when_Pipeline_l124_5;
  reg        [31:0]   memory_to_writeBack_INSTRUCTION;
  wire                when_Pipeline_l124_6;
  reg        [31:0]   decode_to_execute_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_7;
  reg        [31:0]   execute_to_memory_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_8;
  reg        [31:0]   memory_to_writeBack_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_9;
  reg                 decode_to_execute_MEMORY_FORCE_CONSTISTENCY;
  wire                when_Pipeline_l124_10;
  reg                 decode_to_execute_LEGAL_INSTRUCTION;
  wire                when_Pipeline_l124_11;
  reg                 decode_to_execute_MEMORY_FENCE_WR;
  wire                when_Pipeline_l124_12;
  reg                 decode_to_execute_SRC_USE_SUB_LESS;
  wire                when_Pipeline_l124_13;
  reg                 decode_to_execute_MEMORY_ENABLE;
  wire                when_Pipeline_l124_14;
  reg                 execute_to_memory_MEMORY_ENABLE;
  wire                when_Pipeline_l124_15;
  reg                 memory_to_writeBack_MEMORY_ENABLE;
  wire                when_Pipeline_l124_16;
  reg        [1:0]    decode_to_execute_ALU_CTRL;
  wire                when_Pipeline_l124_17;
  reg                 decode_to_execute_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_18;
  reg                 execute_to_memory_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_19;
  reg                 memory_to_writeBack_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_20;
  reg                 decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  wire                when_Pipeline_l124_21;
  reg                 decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_22;
  reg                 execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_23;
  reg                 decode_to_execute_MEMORY_WR;
  wire                when_Pipeline_l124_24;
  reg                 execute_to_memory_MEMORY_WR;
  wire                when_Pipeline_l124_25;
  reg                 memory_to_writeBack_MEMORY_WR;
  wire                when_Pipeline_l124_26;
  reg                 decode_to_execute_HAS_SIDE_EFFECT;
  wire                when_Pipeline_l124_27;
  reg                 execute_to_memory_HAS_SIDE_EFFECT;
  wire                when_Pipeline_l124_28;
  reg                 memory_to_writeBack_HAS_SIDE_EFFECT;
  wire                when_Pipeline_l124_29;
  reg                 decode_to_execute_MEMORY_LRSC;
  wire                when_Pipeline_l124_30;
  reg                 execute_to_memory_MEMORY_LRSC;
  wire                when_Pipeline_l124_31;
  reg                 memory_to_writeBack_MEMORY_LRSC;
  wire                when_Pipeline_l124_32;
  reg                 decode_to_execute_MEMORY_AMO;
  wire                when_Pipeline_l124_33;
  reg                 execute_to_memory_MEMORY_AMO;
  wire                when_Pipeline_l124_34;
  reg                 memory_to_writeBack_MEMORY_AMO;
  wire                when_Pipeline_l124_35;
  reg                 decode_to_execute_MEMORY_MANAGMENT;
  wire                when_Pipeline_l124_36;
  reg                 decode_to_execute_MEMORY_FENCE;
  wire                when_Pipeline_l124_37;
  reg                 execute_to_memory_MEMORY_FENCE;
  wire                when_Pipeline_l124_38;
  reg                 memory_to_writeBack_MEMORY_FENCE;
  wire                when_Pipeline_l124_39;
  reg                 decode_to_execute_IS_CSR;
  wire                when_Pipeline_l124_40;
  reg        [1:0]    decode_to_execute_ENV_CTRL;
  wire                when_Pipeline_l124_41;
  reg        [1:0]    execute_to_memory_ENV_CTRL;
  wire                when_Pipeline_l124_42;
  reg        [1:0]    memory_to_writeBack_ENV_CTRL;
  wire                when_Pipeline_l124_43;
  reg        [1:0]    decode_to_execute_BRANCH_CTRL;
  wire                when_Pipeline_l124_44;
  reg                 decode_to_execute_SRC_LESS_UNSIGNED;
  wire                when_Pipeline_l124_45;
  reg                 decode_to_execute_IS_MUL;
  wire                when_Pipeline_l124_46;
  reg                 execute_to_memory_IS_MUL;
  wire                when_Pipeline_l124_47;
  reg                 memory_to_writeBack_IS_MUL;
  wire                when_Pipeline_l124_48;
  reg                 decode_to_execute_IS_DIV;
  wire                when_Pipeline_l124_49;
  reg                 execute_to_memory_IS_DIV;
  wire                when_Pipeline_l124_50;
  reg                 decode_to_execute_IS_RS1_SIGNED;
  wire                when_Pipeline_l124_51;
  reg                 decode_to_execute_IS_RS2_SIGNED;
  wire                when_Pipeline_l124_52;
  reg                 decode_to_execute_FPU_COMMIT;
  wire                when_Pipeline_l124_53;
  reg                 execute_to_memory_FPU_COMMIT;
  wire                when_Pipeline_l124_54;
  reg                 memory_to_writeBack_FPU_COMMIT;
  wire                when_Pipeline_l124_55;
  reg                 decode_to_execute_FPU_RSP;
  wire                when_Pipeline_l124_56;
  reg                 execute_to_memory_FPU_RSP;
  wire                when_Pipeline_l124_57;
  reg                 memory_to_writeBack_FPU_RSP;
  wire                when_Pipeline_l124_58;
  reg        [3:0]    decode_to_execute_FPU_OPCODE;
  wire                when_Pipeline_l124_59;
  reg        [3:0]    execute_to_memory_FPU_OPCODE;
  wire                when_Pipeline_l124_60;
  reg        [3:0]    memory_to_writeBack_FPU_OPCODE;
  wire                when_Pipeline_l124_61;
  reg                 decode_to_execute_CfuPlugin_CFU_ENABLE;
  wire                when_Pipeline_l124_62;
  reg        [0:0]    decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire                when_Pipeline_l124_63;
  reg        [1:0]    decode_to_execute_ALU_BITWISE_CTRL;
  wire                when_Pipeline_l124_64;
  reg        [1:0]    decode_to_execute_SHIFT_CTRL;
  wire                when_Pipeline_l124_65;
  reg        [1:0]    execute_to_memory_SHIFT_CTRL;
  wire                when_Pipeline_l124_66;
  reg        [31:0]   decode_to_execute_RS1;
  wire                when_Pipeline_l124_67;
  reg        [31:0]   execute_to_memory_RS1;
  wire                when_Pipeline_l124_68;
  reg        [31:0]   memory_to_writeBack_RS1;
  wire                when_Pipeline_l124_69;
  reg        [31:0]   decode_to_execute_RS2;
  wire                when_Pipeline_l124_70;
  reg                 decode_to_execute_SRC2_FORCE_ZERO;
  wire                when_Pipeline_l124_71;
  reg        [31:0]   decode_to_execute_SRC1;
  wire                when_Pipeline_l124_72;
  reg        [31:0]   decode_to_execute_SRC2;
  wire                when_Pipeline_l124_73;
  reg                 decode_to_execute_CSR_WRITE_OPCODE;
  wire                when_Pipeline_l124_74;
  reg                 decode_to_execute_CSR_READ_OPCODE;
  wire                when_Pipeline_l124_75;
  reg                 decode_to_execute_FPU_FORKED;
  wire                when_Pipeline_l124_76;
  reg                 execute_to_memory_FPU_FORKED;
  wire                when_Pipeline_l124_77;
  reg                 memory_to_writeBack_FPU_FORKED;
  wire                when_Pipeline_l124_78;
  reg                 decode_to_execute_FPU_COMMIT_LOAD;
  wire                when_Pipeline_l124_79;
  reg                 execute_to_memory_FPU_COMMIT_LOAD;
  wire                when_Pipeline_l124_80;
  reg                 memory_to_writeBack_FPU_COMMIT_LOAD;
  wire                when_Pipeline_l124_81;
  reg        [31:0]   execute_to_memory_MEMORY_STORE_DATA_RF;
  wire                when_Pipeline_l124_82;
  reg        [31:0]   memory_to_writeBack_MEMORY_STORE_DATA_RF;
  wire                when_Pipeline_l124_83;
  (* keep , syn_keep *) reg        [31:0]   execute_to_memory_MEMORY_VIRTUAL_ADDRESS /* synthesis syn_keep = 1 */ ;
  wire                when_Pipeline_l124_84;
  reg                 execute_to_memory_BRANCH_DO;
  wire                when_Pipeline_l124_85;
  reg        [31:0]   execute_to_memory_BRANCH_CALC;
  wire                when_Pipeline_l124_86;
  reg        [31:0]   execute_to_memory_MUL_LL;
  wire                when_Pipeline_l124_87;
  reg        [33:0]   execute_to_memory_MUL_LH;
  wire                when_Pipeline_l124_88;
  reg        [33:0]   execute_to_memory_MUL_HL;
  wire                when_Pipeline_l124_89;
  reg        [33:0]   execute_to_memory_MUL_HH;
  wire                when_Pipeline_l124_90;
  reg        [33:0]   memory_to_writeBack_MUL_HH;
  wire                when_Pipeline_l124_91;
  reg                 execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
  wire                when_Pipeline_l124_92;
  reg                 memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
  wire                when_Pipeline_l124_93;
  reg        [31:0]   execute_to_memory_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_94;
  reg        [31:0]   memory_to_writeBack_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_95;
  reg        [31:0]   execute_to_memory_SHIFT_RIGHT;
  wire                when_Pipeline_l124_96;
  reg        [51:0]   memory_to_writeBack_MUL_LOW;
  wire                when_Pipeline_l151;
  wire                when_Pipeline_l154;
  wire                when_Pipeline_l151_1;
  wire                when_Pipeline_l154_1;
  wire                when_Pipeline_l151_2;
  wire                when_Pipeline_l154_2;
  reg        [2:0]    IBusCachedPlugin_injector_port_state;
  wire                when_Fetcher_l373;
  wire                when_Fetcher_l391;
  wire                when_Fetcher_l411;
  wire                when_CsrPlugin_l1813;
  reg                 execute_CsrPlugin_csr_1972;
  wire                when_CsrPlugin_l1813_1;
  reg                 execute_CsrPlugin_csr_1969;
  wire                when_CsrPlugin_l1813_2;
  reg                 execute_CsrPlugin_csr_1968;
  wire                when_CsrPlugin_l1813_3;
  reg                 execute_CsrPlugin_csr_3857;
  wire                when_CsrPlugin_l1813_4;
  reg                 execute_CsrPlugin_csr_3858;
  wire                when_CsrPlugin_l1813_5;
  reg                 execute_CsrPlugin_csr_3859;
  wire                when_CsrPlugin_l1813_6;
  reg                 execute_CsrPlugin_csr_3860;
  wire                when_CsrPlugin_l1813_7;
  reg                 execute_CsrPlugin_csr_769;
  wire                when_CsrPlugin_l1813_8;
  reg                 execute_CsrPlugin_csr_768;
  wire                when_CsrPlugin_l1813_9;
  reg                 execute_CsrPlugin_csr_836;
  wire                when_CsrPlugin_l1813_10;
  reg                 execute_CsrPlugin_csr_772;
  wire                when_CsrPlugin_l1813_11;
  reg                 execute_CsrPlugin_csr_773;
  wire                when_CsrPlugin_l1813_12;
  reg                 execute_CsrPlugin_csr_833;
  wire                when_CsrPlugin_l1813_13;
  reg                 execute_CsrPlugin_csr_832;
  wire                when_CsrPlugin_l1813_14;
  reg                 execute_CsrPlugin_csr_834;
  wire                when_CsrPlugin_l1813_15;
  reg                 execute_CsrPlugin_csr_835;
  wire                when_CsrPlugin_l1813_16;
  reg                 execute_CsrPlugin_csr_3;
  wire                when_CsrPlugin_l1813_17;
  reg                 execute_CsrPlugin_csr_2;
  wire                when_CsrPlugin_l1813_18;
  reg                 execute_CsrPlugin_csr_1;
  wire                when_CsrPlugin_l1813_19;
  reg                 execute_CsrPlugin_csr_256;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_1;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_3;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_4;
  wire       [1:0]    switch_CsrPlugin_l1167;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_5;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_6;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_7;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_8;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_9;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_10;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_11;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_12;
  wire       [4:0]    _zz_FpuPlugin_flags_NX;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_13;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_14;
  wire       [4:0]    _zz_FpuPlugin_flags_NX_1;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_15;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_16;
  wire                when_CsrPlugin_l1846;
  wire       [11:0]   _zz_when_CsrPlugin_l1853;
  wire                when_CsrPlugin_l1853;
  reg                 when_CsrPlugin_l1863;
  wire                when_CsrPlugin_l1861;
  wire                when_CsrPlugin_l1862;
  wire                when_CsrPlugin_l1869;
  reg        [2:0]    FpuPlugin_stateReg;
  reg        [2:0]    FpuPlugin_stateNext;
  reg        [0:0]    _zz_FpuPlugin_port_cmd_payload_format;
  wire                when_FpuPlugin_l402;
  `ifndef SYNTHESIS
  reg [71:0] _zz_execute_to_memory_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_to_memory_SHIFT_CTRL_1_string;
  reg [71:0] decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_1_string;
  reg [39:0] decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string;
  reg [39:0] decode_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string;
  reg [63:0] memory_FPU_OPCODE_string;
  reg [63:0] _zz_memory_FPU_OPCODE_string;
  reg [63:0] _zz_memory_to_writeBack_FPU_OPCODE_string;
  reg [63:0] _zz_memory_to_writeBack_FPU_OPCODE_1_string;
  reg [63:0] execute_FPU_OPCODE_string;
  reg [63:0] _zz_execute_FPU_OPCODE_string;
  reg [63:0] _zz_execute_to_memory_FPU_OPCODE_string;
  reg [63:0] _zz_execute_to_memory_FPU_OPCODE_1_string;
  reg [63:0] _zz_decode_to_execute_FPU_OPCODE_string;
  reg [63:0] _zz_decode_to_execute_FPU_OPCODE_1_string;
  reg [31:0] decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_1_string;
  reg [47:0] _zz_memory_to_writeBack_ENV_CTRL_string;
  reg [47:0] _zz_memory_to_writeBack_ENV_CTRL_1_string;
  reg [47:0] _zz_execute_to_memory_ENV_CTRL_string;
  reg [47:0] _zz_execute_to_memory_ENV_CTRL_1_string;
  reg [47:0] decode_ENV_CTRL_string;
  reg [47:0] _zz_decode_ENV_CTRL_string;
  reg [47:0] _zz_decode_to_execute_ENV_CTRL_string;
  reg [47:0] _zz_decode_to_execute_ENV_CTRL_1_string;
  reg [63:0] decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_1_string;
  reg [71:0] memory_SHIFT_CTRL_string;
  reg [71:0] _zz_memory_SHIFT_CTRL_string;
  reg [71:0] execute_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_SHIFT_CTRL_string;
  reg [63:0] execute_ALU_CTRL_string;
  reg [63:0] _zz_execute_ALU_CTRL_string;
  reg [39:0] execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [63:0] writeBack_FPU_OPCODE_string;
  reg [63:0] _zz_writeBack_FPU_OPCODE_string;
  reg [47:0] decode_FPU_FORMAT_string;
  reg [47:0] _zz_decode_FPU_FORMAT_string;
  reg [63:0] decode_FPU_OPCODE_string;
  reg [63:0] _zz_decode_FPU_OPCODE_string;
  reg [31:0] execute_BRANCH_CTRL_string;
  reg [31:0] _zz_execute_BRANCH_CTRL_string;
  reg [47:0] memory_ENV_CTRL_string;
  reg [47:0] _zz_memory_ENV_CTRL_string;
  reg [47:0] execute_ENV_CTRL_string;
  reg [47:0] _zz_execute_ENV_CTRL_string;
  reg [47:0] writeBack_ENV_CTRL_string;
  reg [47:0] _zz_writeBack_ENV_CTRL_string;
  reg [23:0] decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_SRC2_CTRL_string;
  reg [95:0] decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_SRC1_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_1_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_1_string;
  reg [39:0] _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string;
  reg [47:0] _zz_decode_FPU_FORMAT_1_string;
  reg [63:0] _zz_decode_FPU_OPCODE_1_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_1_string;
  reg [47:0] _zz_decode_ENV_CTRL_1_string;
  reg [23:0] _zz_decode_SRC2_CTRL_1_string;
  reg [63:0] _zz_decode_ALU_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_1_string;
  reg [71:0] debugBus_dmToHart_payload_op_string;
  reg [63:0] FpuPlugin_port_cmd_payload_opcode_string;
  reg [47:0] FpuPlugin_port_cmd_payload_format_string;
  reg [23:0] FpuPlugin_port_cmd_payload_roundMode_string;
  reg [63:0] FpuPlugin_port_commit_payload_opcode_string;
  reg [95:0] _zz_decode_SRC1_CTRL_2_string;
  reg [63:0] _zz_decode_ALU_CTRL_2_string;
  reg [23:0] _zz_decode_SRC2_CTRL_2_string;
  reg [47:0] _zz_decode_ENV_CTRL_2_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_2_string;
  reg [63:0] _zz_decode_FPU_OPCODE_2_string;
  reg [47:0] _zz_decode_FPU_FORMAT_2_string;
  reg [39:0] _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_2_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_2_string;
  reg [71:0] CsrPlugin_inject_cmd_payload_op_string;
  reg [71:0] CsrPlugin_inject_cmd_toStream_payload_op_string;
  reg [71:0] CsrPlugin_inject_buffer_payload_op_string;
  reg [71:0] CsrPlugin_inject_cmd_toStream_rData_op_string;
  reg [47:0] CsrPlugin_dcsr_stepLogic_stateReg_string;
  reg [47:0] CsrPlugin_dcsr_stepLogic_stateNext_string;
  reg [23:0] _zz_FpuPlugin_port_cmd_payload_roundMode_string;
  reg [23:0] _zz_FpuPlugin_port_cmd_payload_roundMode_1_string;
  reg [63:0] writeBack_FpuPlugin_commit_payload_opcode_string;
  reg [63:0] writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string;
  reg [63:0] writeBack_FpuPlugin_commit_rData_opcode_string;
  reg [63:0] _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string;
  reg [63:0] decode_to_execute_ALU_CTRL_string;
  reg [47:0] decode_to_execute_ENV_CTRL_string;
  reg [47:0] execute_to_memory_ENV_CTRL_string;
  reg [47:0] memory_to_writeBack_ENV_CTRL_string;
  reg [31:0] decode_to_execute_BRANCH_CTRL_string;
  reg [63:0] decode_to_execute_FPU_OPCODE_string;
  reg [63:0] execute_to_memory_FPU_OPCODE_string;
  reg [63:0] memory_to_writeBack_FPU_OPCODE_string;
  reg [39:0] decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [71:0] decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] execute_to_memory_SHIFT_CTRL_string;
  reg [47:0] FpuPlugin_stateReg_string;
  reg [47:0] FpuPlugin_stateNext_string;
  reg [47:0] _zz_FpuPlugin_port_cmd_payload_format_string;
  `endif

  reg [31:0] RegFilePlugin_regFile [0:31] /* verilator public */ ;

  assign _zz_when = (|{decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid});
  assign _zz_memory_MUL_LOW = ($signed(_zz_memory_MUL_LOW_1) + $signed(_zz_memory_MUL_LOW_4));
  assign _zz_memory_MUL_LOW_1 = ($signed(52'h0) + $signed(_zz_memory_MUL_LOW_2));
  assign _zz_memory_MUL_LOW_3 = {1'b0,memory_MUL_LL};
  assign _zz_memory_MUL_LOW_2 = {{19{_zz_memory_MUL_LOW_3[32]}}, _zz_memory_MUL_LOW_3};
  assign _zz_memory_MUL_LOW_5 = ({16'd0,memory_MUL_LH} <<< 5'd16);
  assign _zz_memory_MUL_LOW_4 = {{2{_zz_memory_MUL_LOW_5[49]}}, _zz_memory_MUL_LOW_5};
  assign _zz_memory_MUL_LOW_7 = ({16'd0,memory_MUL_HL} <<< 5'd16);
  assign _zz_memory_MUL_LOW_6 = {{2{_zz_memory_MUL_LOW_7[49]}}, _zz_memory_MUL_LOW_7};
  assign _zz_decode_FORMAL_PC_NEXT_1 = (decode_IS_RVC ? 3'b010 : 3'b100);
  assign _zz_decode_FORMAL_PC_NEXT = {29'd0, _zz_decode_FORMAL_PC_NEXT_1};
  assign _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload - 3'b001);
  assign _zz_IBusCachedPlugin_fetchPc_pc_1 = {IBusCachedPlugin_fetchPc_inc,2'b00};
  assign _zz_IBusCachedPlugin_fetchPc_pc = {29'd0, _zz_IBusCachedPlugin_fetchPc_pc_1};
  assign _zz_IBusCachedPlugin_decodePc_pcPlus_1 = (decode_IS_RVC ? 3'b010 : 3'b100);
  assign _zz_IBusCachedPlugin_decodePc_pcPlus = {29'd0, _zz_IBusCachedPlugin_decodePc_pcPlus_1};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_31 = {{_zz_IBusCachedPlugin_decompressor_decompressed_11,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},12'h0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_38 = {{{3'b000,_zz_IBusCachedPlugin_decompressor_decompressed[9 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},3'b000};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_39 = {{{3'b000,_zz_IBusCachedPlugin_decompressor_decompressed[9 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},3'b000};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_40 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_41 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_42 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_43 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_io_cpu_flush_payload_lineId = _zz_io_cpu_flush_payload_lineId_1;
  assign _zz_io_cpu_flush_payload_lineId_1 = (execute_RS1 >>> 3'd6);
  assign _zz_DBusCachedPlugin_exceptionBus_payload_code = (writeBack_MEMORY_WR ? 3'b111 : 3'b101);
  assign _zz_DBusCachedPlugin_exceptionBus_payload_code_1 = (writeBack_MEMORY_WR ? 3'b110 : 3'b100);
  assign _zz_writeBack_DBusCachedPlugin_rspRf = (! dataCache_2_io_cpu_writeBack_exclusiveOk);
  assign _zz__zz_decode_SRC1 = (decode_IS_RVC ? 3'b010 : 3'b100);
  assign _zz__zz_decode_SRC1_1 = decode_INSTRUCTION[19 : 15];
  assign _zz__zz_decode_SRC2_2 = {decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]};
  assign _zz_execute_SrcPlugin_addSub = ($signed(_zz_execute_SrcPlugin_addSub_1) + $signed(_zz_execute_SrcPlugin_addSub_4));
  assign _zz_execute_SrcPlugin_addSub_1 = ($signed(_zz_execute_SrcPlugin_addSub_2) + $signed(_zz_execute_SrcPlugin_addSub_3));
  assign _zz_execute_SrcPlugin_addSub_2 = execute_SRC1;
  assign _zz_execute_SrcPlugin_addSub_3 = (execute_SRC_USE_SUB_LESS ? (~ execute_SRC2) : execute_SRC2);
  assign _zz_execute_SrcPlugin_addSub_4 = (execute_SRC_USE_SUB_LESS ? 32'h00000001 : 32'h0);
  assign _zz_CsrPlugin_timeout_counter_valueNext_1 = CsrPlugin_timeout_counter_willIncrement;
  assign _zz_CsrPlugin_timeout_counter_valueNext = {2'd0, _zz_CsrPlugin_timeout_counter_valueNext_1};
  assign _zz__zz_6 = debugBus_dmToHart_payload_address[0:0];
  assign _zz_CsrPlugin_counters_mcycle_1 = ((! debugMode) || (! CsrPlugin_dcsr_stopcount));
  assign _zz_CsrPlugin_counters_mcycle = {63'd0, _zz_CsrPlugin_counters_mcycle_1};
  assign _zz_CsrPlugin_counters_minstret_1 = ((! debugMode) || (! CsrPlugin_dcsr_stopcount));
  assign _zz_CsrPlugin_counters_minstret = {63'd0, _zz_CsrPlugin_counters_minstret_1};
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code & (~ _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1));
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code - 2'b01);
  assign _zz__zz_execute_BranchPlugin_branch_src2 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]};
  assign _zz__zz_execute_BranchPlugin_branch_src2_4 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]};
  assign _zz_writeBack_MulPlugin_result = {{14{writeBack_MUL_LOW[51]}}, writeBack_MUL_LOW};
  assign _zz_writeBack_MulPlugin_result_1 = ({32'd0,writeBack_MUL_HH} <<< 6'd32);
  assign _zz__zz_decode_RS2_2 = writeBack_MUL_LOW[31 : 0];
  assign _zz__zz_decode_RS2_2_1 = writeBack_MulPlugin_result[63 : 32];
  assign _zz_memory_MulDivIterativePlugin_div_counter_valueNext_1 = memory_MulDivIterativePlugin_div_counter_willIncrement;
  assign _zz_memory_MulDivIterativePlugin_div_counter_valueNext = {5'd0, _zz_memory_MulDivIterativePlugin_div_counter_valueNext_1};
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator = {1'd0, memory_MulDivIterativePlugin_rs2};
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder = memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator[31:0];
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder_1 = memory_MulDivIterativePlugin_div_stage_0_remainderShifted[31:0];
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_outNumerator = {_zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted,(! memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator[32])};
  assign _zz_memory_MulDivIterativePlugin_div_result_1 = _zz_memory_MulDivIterativePlugin_div_result_2;
  assign _zz_memory_MulDivIterativePlugin_div_result_2 = _zz_memory_MulDivIterativePlugin_div_result_3;
  assign _zz_memory_MulDivIterativePlugin_div_result_3 = ({memory_MulDivIterativePlugin_div_needRevert,(memory_MulDivIterativePlugin_div_needRevert ? (~ _zz_memory_MulDivIterativePlugin_div_result) : _zz_memory_MulDivIterativePlugin_div_result)} + _zz_memory_MulDivIterativePlugin_div_result_4);
  assign _zz_memory_MulDivIterativePlugin_div_result_5 = memory_MulDivIterativePlugin_div_needRevert;
  assign _zz_memory_MulDivIterativePlugin_div_result_4 = {32'd0, _zz_memory_MulDivIterativePlugin_div_result_5};
  assign _zz_memory_MulDivIterativePlugin_rs1_3 = _zz_memory_MulDivIterativePlugin_rs1;
  assign _zz_memory_MulDivIterativePlugin_rs1_2 = {32'd0, _zz_memory_MulDivIterativePlugin_rs1_3};
  assign _zz_memory_MulDivIterativePlugin_rs2_2 = _zz_memory_MulDivIterativePlugin_rs2;
  assign _zz_memory_MulDivIterativePlugin_rs2_1 = {31'd0, _zz_memory_MulDivIterativePlugin_rs2_2};
  assign _zz_FpuPlugin_pendings = (_zz_FpuPlugin_pendings_1 - _zz_FpuPlugin_pendings_4);
  assign _zz_FpuPlugin_pendings_1 = (FpuPlugin_pendings + _zz_FpuPlugin_pendings_2);
  assign _zz_FpuPlugin_pendings_3 = FpuPlugin_port_cmd_fire;
  assign _zz_FpuPlugin_pendings_2 = {5'd0, _zz_FpuPlugin_pendings_3};
  assign _zz_FpuPlugin_pendings_5 = FpuPlugin_port_completion_valid;
  assign _zz_FpuPlugin_pendings_4 = {5'd0, _zz_FpuPlugin_pendings_5};
  assign _zz_FpuPlugin_pendings_7 = FpuPlugin_port_rsp_fire;
  assign _zz_FpuPlugin_pendings_6 = {5'd0, _zz_FpuPlugin_pendings_7};
  assign _zz_when_CsrPlugin_l1862 = (execute_CsrPlugin_csrAddress >>> 3'd4);
  assign _zz_decode_RegFilePlugin_rs1Data = 1'b1;
  assign _zz_decode_RegFilePlugin_rs2Data = 1'b1;
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_5 = {_zz_IBusCachedPlugin_jump_pcLoad_payload_3,_zz_IBusCachedPlugin_jump_pcLoad_payload_2};
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_1 = dataCache_2_io_cpu_writeBack_address[2 : 0];
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_3 = dataCache_2_io_cpu_writeBack_address[2 : 1];
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_5 = dataCache_2_io_cpu_writeBack_address[2 : 2];
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_7 = dataCache_2_io_cpu_writeBack_address[2 : 2];
  assign _zz_decode_LEGAL_INSTRUCTION = 32'h0000007f;
  assign _zz_decode_LEGAL_INSTRUCTION_1 = (decode_INSTRUCTION & 32'h0000007f);
  assign _zz_decode_LEGAL_INSTRUCTION_2 = 32'h0000000b;
  assign _zz_decode_LEGAL_INSTRUCTION_3 = ((decode_INSTRUCTION & 32'h0000107f) == 32'h00001073);
  assign _zz_decode_LEGAL_INSTRUCTION_4 = ((decode_INSTRUCTION & 32'h0000207f) == 32'h00002073);
  assign _zz_decode_LEGAL_INSTRUCTION_5 = {((decode_INSTRUCTION & 32'h0000407f) == 32'h00004063),{((decode_INSTRUCTION & 32'h0000207f) == 32'h00002013),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_6) == 32'h00002007),{(_zz_decode_LEGAL_INSTRUCTION_7 == _zz_decode_LEGAL_INSTRUCTION_8),{_zz_decode_LEGAL_INSTRUCTION_9,{_zz_decode_LEGAL_INSTRUCTION_10,_zz_decode_LEGAL_INSTRUCTION_11}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_6 = 32'h0000605f;
  assign _zz_decode_LEGAL_INSTRUCTION_7 = (decode_INSTRUCTION & 32'h0000705b);
  assign _zz_decode_LEGAL_INSTRUCTION_8 = 32'h00002003;
  assign _zz_decode_LEGAL_INSTRUCTION_9 = ((decode_INSTRUCTION & 32'h0000107f) == 32'h00000013);
  assign _zz_decode_LEGAL_INSTRUCTION_10 = ((decode_INSTRUCTION & 32'h0000603f) == 32'h00000023);
  assign _zz_decode_LEGAL_INSTRUCTION_11 = {((decode_INSTRUCTION & 32'h0000207f) == 32'h00000003),{((decode_INSTRUCTION & 32'h0000707b) == 32'h00000063),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_12) == 32'h0000000f),{(_zz_decode_LEGAL_INSTRUCTION_13 == _zz_decode_LEGAL_INSTRUCTION_14),{_zz_decode_LEGAL_INSTRUCTION_15,{_zz_decode_LEGAL_INSTRUCTION_16,_zz_decode_LEGAL_INSTRUCTION_17}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_12 = 32'h0000607f;
  assign _zz_decode_LEGAL_INSTRUCTION_13 = (decode_INSTRUCTION & 32'he400007f);
  assign _zz_decode_LEGAL_INSTRUCTION_14 = 32'h00000053;
  assign _zz_decode_LEGAL_INSTRUCTION_15 = ((decode_INSTRUCTION & 32'h1800707f) == 32'h0000202f);
  assign _zz_decode_LEGAL_INSTRUCTION_16 = ((decode_INSTRUCTION & 32'hfc00007f) == 32'h00000033);
  assign _zz_decode_LEGAL_INSTRUCTION_17 = {((decode_INSTRUCTION & 32'he800707f) == 32'h0800202f),{((decode_INSTRUCTION & 32'h7c00607f) == 32'h20000053),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_18) == 32'h20000053),{(_zz_decode_LEGAL_INSTRUCTION_19 == _zz_decode_LEGAL_INSTRUCTION_20),{_zz_decode_LEGAL_INSTRUCTION_21,{_zz_decode_LEGAL_INSTRUCTION_22,_zz_decode_LEGAL_INSTRUCTION_23}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_18 = 32'h7c00507f;
  assign _zz_decode_LEGAL_INSTRUCTION_19 = (decode_INSTRUCTION & 32'hf400607f);
  assign _zz_decode_LEGAL_INSTRUCTION_20 = 32'h20000053;
  assign _zz_decode_LEGAL_INSTRUCTION_21 = ((decode_INSTRUCTION & 32'h01f0707f) == 32'h0000500f);
  assign _zz_decode_LEGAL_INSTRUCTION_22 = ((decode_INSTRUCTION & 32'hbe00705f) == 32'h00005013);
  assign _zz_decode_LEGAL_INSTRUCTION_23 = {((decode_INSTRUCTION & 32'hfe00305f) == 32'h00001013),{((decode_INSTRUCTION & 32'hede0007f) == 32'hc0000053),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_24) == 32'h00000033),{(_zz_decode_LEGAL_INSTRUCTION_25 == _zz_decode_LEGAL_INSTRUCTION_26),{_zz_decode_LEGAL_INSTRUCTION_27,{_zz_decode_LEGAL_INSTRUCTION_28,_zz_decode_LEGAL_INSTRUCTION_29}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_24 = 32'hbe00707f;
  assign _zz_decode_LEGAL_INSTRUCTION_25 = (decode_INSTRUCTION & 32'hfdf0007f);
  assign _zz_decode_LEGAL_INSTRUCTION_26 = 32'h58000053;
  assign _zz_decode_LEGAL_INSTRUCTION_27 = ((decode_INSTRUCTION & 32'h7ff0007f) == 32'h42000053);
  assign _zz_decode_LEGAL_INSTRUCTION_28 = ((decode_INSTRUCTION & 32'h7ff0007f) == 32'h40100053);
  assign _zz_decode_LEGAL_INSTRUCTION_29 = {((decode_INSTRUCTION & 32'hf9f0707f) == 32'h1000202f),{((decode_INSTRUCTION & 32'hfdf0707f) == 32'he0001053),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_30) == 32'he0000053),{(_zz_decode_LEGAL_INSTRUCTION_31 == _zz_decode_LEGAL_INSTRUCTION_32),{_zz_decode_LEGAL_INSTRUCTION_33,_zz_decode_LEGAL_INSTRUCTION_34}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_30 = 32'heff0707f;
  assign _zz_decode_LEGAL_INSTRUCTION_31 = (decode_INSTRUCTION & 32'hdfffffff);
  assign _zz_decode_LEGAL_INSTRUCTION_32 = 32'h10200073;
  assign _zz_decode_LEGAL_INSTRUCTION_33 = ((decode_INSTRUCTION & 32'hffefffff) == 32'h00000073);
  assign _zz_decode_LEGAL_INSTRUCTION_34 = ((decode_INSTRUCTION & 32'hffffffff) == 32'h10500073);
  assign _zz_IBusCachedPlugin_decompressor_decompressed_28 = {_zz_IBusCachedPlugin_decompressor_decompressed_13,_zz_IBusCachedPlugin_decompressor_decompressed[4 : 3]};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_29 = _zz_IBusCachedPlugin_decompressor_decompressed[5];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_30 = _zz_IBusCachedPlugin_decompressor_decompressed[2];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_32 = (_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] == 2'b01);
  assign _zz_IBusCachedPlugin_decompressor_decompressed_33 = ((_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] == 2'b11) && (_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5] == 2'b00));
  assign _zz_IBusCachedPlugin_decompressor_decompressed_34 = 7'h0;
  assign _zz_IBusCachedPlugin_decompressor_decompressed_35 = _zz_IBusCachedPlugin_decompressor_decompressed[6 : 2];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_36 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_37 = _zz_IBusCachedPlugin_decompressor_decompressed[11 : 7];
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE = (decode_INSTRUCTION & 32'h40003054);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_1 = 32'h40001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_2 = (decode_INSTRUCTION & 32'h02007054);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_3 = 32'h00001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_4 = (decode_INSTRUCTION & 32'h00001000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_5 = 32'h00001000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_6 = ((decode_INSTRUCTION & 32'h00003000) == 32'h00002000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_7 = (|_zz_decode_CfuPlugin_CFU_ENABLE_10);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_8 = (|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE_9 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_10),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_11 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_12)});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_13 = {(|{_zz_decode_CfuPlugin_CFU_ENABLE_7,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_14,_zz__zz_decode_CfuPlugin_CFU_ENABLE_17}}),{(|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_22,_zz__zz_decode_CfuPlugin_CFU_ENABLE_25}),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_40),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_49,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_58,_zz__zz_decode_CfuPlugin_CFU_ENABLE_70}}}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_9 = (decode_INSTRUCTION & 32'h00000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_10 = 32'h00000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_11 = (decode_INSTRUCTION & 32'h20002010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_12 = 32'h20002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_14 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_15 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_16);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_17 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_18,_zz__zz_decode_CfuPlugin_CFU_ENABLE_20};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_22 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_23 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_24);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_25 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_26,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_28,_zz__zz_decode_CfuPlugin_CFU_ENABLE_31}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_40 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_41,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_43,_zz__zz_decode_CfuPlugin_CFU_ENABLE_46}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_49 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_50,_zz__zz_decode_CfuPlugin_CFU_ENABLE_53});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_58 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_59);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_70 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_71,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_80,_zz__zz_decode_CfuPlugin_CFU_ENABLE_82}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_15 = (decode_INSTRUCTION & 32'h20001010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_16 = 32'h20001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_18 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_19) == 32'h08000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_20 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_21) == 32'h80000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_23 = (decode_INSTRUCTION & 32'h00001040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_24 = 32'h00001000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_26 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_27) == 32'h82000000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_28 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_29 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_30);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_31 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_32,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_34,_zz__zz_decode_CfuPlugin_CFU_ENABLE_37}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_41 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_42) == 32'h60000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_43 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_44 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_45);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_46 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_47,_zz_decode_CfuPlugin_CFU_ENABLE_13};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_50 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_51 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_52);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_53 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_54,_zz__zz_decode_CfuPlugin_CFU_ENABLE_56};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_59 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_60,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_62,_zz__zz_decode_CfuPlugin_CFU_ENABLE_65}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_71 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_72,_zz__zz_decode_CfuPlugin_CFU_ENABLE_73});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_80 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_81);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_82 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_83,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_90,_zz__zz_decode_CfuPlugin_CFU_ENABLE_94}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_19 = 32'h28000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_21 = 32'ha0100010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_27 = 32'h82000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_29 = (decode_INSTRUCTION & 32'h02000050);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_30 = 32'h02000040;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_32 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_33) == 32'h12000000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_34 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_35 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_36);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_37 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_38 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_39);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_42 = 32'h60000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_44 = (decode_INSTRUCTION & 32'h18000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_45 = 32'h18000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_47 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_48) == 32'h20000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_51 = (decode_INSTRUCTION & 32'h80000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_52 = 32'h80000000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_54 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_55) == 32'h00000040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_56 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_57) == 32'h40000000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_60 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_61) == 32'h00001010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_62 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_63 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_64);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_65 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_66,_zz__zz_decode_CfuPlugin_CFU_ENABLE_68};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_72 = _zz_decode_CfuPlugin_CFU_ENABLE_12;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_73 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_74,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_76,_zz__zz_decode_CfuPlugin_CFU_ENABLE_77}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_81 = {_zz_decode_CfuPlugin_CFU_ENABLE_12,_zz_decode_CfuPlugin_CFU_ENABLE_8};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_83 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_84,_zz__zz_decode_CfuPlugin_CFU_ENABLE_87});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_90 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_91);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_94 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_95,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_96,_zz__zz_decode_CfuPlugin_CFU_ENABLE_98}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_33 = 32'h12000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_35 = (decode_INSTRUCTION & 32'h42000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_36 = 32'h02000000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_38 = (decode_INSTRUCTION & 32'hd2000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_39 = 32'h40000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_48 = 32'ha0000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_55 = 32'h00000050;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_57 = 32'h50000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_61 = 32'h10001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_63 = (decode_INSTRUCTION & 32'h30000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_64 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_66 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_67) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_68 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_69) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_74 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_75) == 32'h90000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_76 = _zz_decode_CfuPlugin_CFU_ENABLE_13;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_77 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_78,_zz__zz_decode_CfuPlugin_CFU_ENABLE_79};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_84 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_85 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_86);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_87 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_88,_zz__zz_decode_CfuPlugin_CFU_ENABLE_89};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_91 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_92,_zz__zz_decode_CfuPlugin_CFU_ENABLE_93};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_95 = (|_zz_decode_CfuPlugin_CFU_ENABLE_11);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_96 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_97);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_98 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_99,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_102,_zz__zz_decode_CfuPlugin_CFU_ENABLE_104}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_67 = 32'h88000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_69 = 32'h50000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_75 = 32'h90000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_78 = ((decode_INSTRUCTION & 32'h58000010) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_79 = ((decode_INSTRUCTION & 32'hb0000010) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_85 = (decode_INSTRUCTION & 32'h10000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_86 = 32'h10000000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_88 = ((decode_INSTRUCTION & 32'h80000020) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_89 = ((decode_INSTRUCTION & 32'h00000030) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_92 = ((decode_INSTRUCTION & 32'h00000060) == 32'h00000040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_93 = ((decode_INSTRUCTION & 32'h0000005c) == 32'h00000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_97 = _zz_decode_CfuPlugin_CFU_ENABLE_11;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_99 = (|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_100 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_101));
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_102 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_103);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_104 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_105),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_108,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_113,_zz__zz_decode_CfuPlugin_CFU_ENABLE_116}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_100 = (decode_INSTRUCTION & 32'h02004064);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_101 = 32'h02004020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_103 = ((decode_INSTRUCTION & 32'h02004074) == 32'h02000030);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_105 = {((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_106) == 32'h00002000),((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_107) == 32'h00001000)};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_108 = (|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE_109 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_110),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_111 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_112)});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_113 = (|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_114 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_115));
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_116 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_117),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_118),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_121,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_126,_zz__zz_decode_CfuPlugin_CFU_ENABLE_129}}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_106 = 32'h00002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_107 = 32'h00005000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_109 = (decode_INSTRUCTION & 32'h00000068);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_110 = 32'h00000068;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_111 = (decode_INSTRUCTION & 32'h00002034);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_112 = 32'h00000024;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_114 = (decode_INSTRUCTION & 32'h00000078);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_115 = 32'h00000060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_117 = ((decode_INSTRUCTION & 32'h10003070) == 32'h00000070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_118 = {((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_119) == 32'h00100070),((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_120) == 32'h10000030)};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_121 = (|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE_122 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_123),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_124 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_125)});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_126 = (|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_127 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_128));
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_129 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_130),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_131),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_136,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_146,_zz__zz_decode_CfuPlugin_CFU_ENABLE_148}}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_119 = 32'h10103070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_120 = 32'h10403034;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_122 = (decode_INSTRUCTION & 32'h00001070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_123 = 32'h00001070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_124 = (decode_INSTRUCTION & 32'h00002070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_125 = 32'h00002070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_127 = (decode_INSTRUCTION & 32'h00003054);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_128 = 32'h00000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_130 = ((decode_INSTRUCTION & 32'h00004054) == 32'h00004004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_131 = {(_zz__zz_decode_CfuPlugin_CFU_ENABLE_132 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_133),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_134 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_135)};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_136 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_137,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_138,_zz__zz_decode_CfuPlugin_CFU_ENABLE_139}});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_146 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_147);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_148 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_149),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_151,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_166,_zz__zz_decode_CfuPlugin_CFU_ENABLE_175}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_132 = (decode_INSTRUCTION & 32'h00000034);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_133 = 32'h00000034;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_134 = (decode_INSTRUCTION & 32'h00000068);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_135 = 32'h00000028;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_137 = ((decode_INSTRUCTION & 32'h00000034) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_138 = _zz_decode_CfuPlugin_CFU_ENABLE_10;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_139 = {(_zz__zz_decode_CfuPlugin_CFU_ENABLE_140 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_141),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_142,_zz__zz_decode_CfuPlugin_CFU_ENABLE_144}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_147 = ((decode_INSTRUCTION & 32'h10000008) == 32'h00000008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_149 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_150) == 32'h10000008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_151 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_152,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_154,_zz__zz_decode_CfuPlugin_CFU_ENABLE_157}});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_166 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_167,_zz__zz_decode_CfuPlugin_CFU_ENABLE_170});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_175 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_176),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_189,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_202,_zz__zz_decode_CfuPlugin_CFU_ENABLE_220}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_140 = (decode_INSTRUCTION & 32'h00000064);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_141 = 32'h00000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_142 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_143) == 32'h08002008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_144 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_145) == 32'h00002008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_150 = 32'h10000008;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_152 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_153) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_154 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_155 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_156);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_157 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_158,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_160,_zz__zz_decode_CfuPlugin_CFU_ENABLE_163}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_167 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_168 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_169);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_170 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_171,_zz__zz_decode_CfuPlugin_CFU_ENABLE_173};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_176 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_177,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_179,_zz__zz_decode_CfuPlugin_CFU_ENABLE_182}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_189 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_190,_zz__zz_decode_CfuPlugin_CFU_ENABLE_191});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_202 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_203);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_220 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_221,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_226,_zz__zz_decode_CfuPlugin_CFU_ENABLE_232}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_143 = 32'h08002048;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_145 = 32'h10002048;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_153 = 32'h00000030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_155 = (decode_INSTRUCTION & 32'h00001060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_156 = 32'h00001060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_158 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_159) == 32'h00002060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_160 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_161 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_162);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_163 = {_zz_decode_CfuPlugin_CFU_ENABLE_4,_zz__zz_decode_CfuPlugin_CFU_ENABLE_164};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_168 = (decode_INSTRUCTION & 32'h08000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_169 = 32'h08000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_171 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_172) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_173 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_174) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_177 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_178) == 32'h00004020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_179 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_180 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_181);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_182 = {_zz_decode_CfuPlugin_CFU_ENABLE_9,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_183,_zz__zz_decode_CfuPlugin_CFU_ENABLE_186}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_190 = _zz_decode_CfuPlugin_CFU_ENABLE_9;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_191 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_192,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_194,_zz__zz_decode_CfuPlugin_CFU_ENABLE_197}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_203 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_204,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_206,_zz__zz_decode_CfuPlugin_CFU_ENABLE_209}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_221 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_222,_zz__zz_decode_CfuPlugin_CFU_ENABLE_223});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_226 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_227);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_232 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_233,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_236,_zz__zz_decode_CfuPlugin_CFU_ENABLE_240}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_159 = 32'h00002060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_161 = (decode_INSTRUCTION & 32'h10000060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_162 = 32'h00000060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_164 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_165) == 32'h10000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_172 = 32'h10000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_174 = 32'h00000028;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_178 = 32'h00004020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_180 = (decode_INSTRUCTION & 32'h00000060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_181 = 32'h00000060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_183 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_184 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_185);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_186 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_187 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_188);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_192 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_193) == 32'h00002010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_194 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_195 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_196);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_197 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_198,_zz__zz_decode_CfuPlugin_CFU_ENABLE_200};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_204 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_205) == 32'h00000028);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_206 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_207 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_208);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_209 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_210,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_212,_zz__zz_decode_CfuPlugin_CFU_ENABLE_215}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_222 = _zz_decode_CfuPlugin_CFU_ENABLE_7;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_223 = {_zz_decode_CfuPlugin_CFU_ENABLE_3,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_224,_zz__zz_decode_CfuPlugin_CFU_ENABLE_225}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_227 = {_zz_decode_CfuPlugin_CFU_ENABLE_7,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_228,_zz__zz_decode_CfuPlugin_CFU_ENABLE_231}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_233 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_234);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_236 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_237);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_240 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_241,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_256,_zz__zz_decode_CfuPlugin_CFU_ENABLE_258}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_165 = 32'h10400024;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_184 = (decode_INSTRUCTION & 32'h82000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_185 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_187 = (decode_INSTRUCTION & 32'h00000070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_188 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_193 = 32'h00002070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_195 = (decode_INSTRUCTION & 32'h00001070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_196 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_198 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_199) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_200 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_201) == 32'h00002020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_205 = 32'h00000028;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_207 = (decode_INSTRUCTION & 32'h00000050);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_208 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_210 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_211) == 32'h00001030);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_212 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_213 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_214);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_215 = {_zz_decode_CfuPlugin_CFU_ENABLE_8,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_216,_zz__zz_decode_CfuPlugin_CFU_ENABLE_218}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_224 = _zz_decode_CfuPlugin_CFU_ENABLE_6;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_225 = _zz_decode_CfuPlugin_CFU_ENABLE_5;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_228 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_229 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_230);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_231 = _zz_decode_CfuPlugin_CFU_ENABLE_6;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_234 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_235) == 32'h00004010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_237 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_238 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_239);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_241 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_242,_zz__zz_decode_CfuPlugin_CFU_ENABLE_244});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_256 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_257);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_258 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_259,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_268,_zz__zz_decode_CfuPlugin_CFU_ENABLE_274}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_199 = 32'h02003020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_201 = 32'h02002068;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_211 = 32'h00001030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_213 = (decode_INSTRUCTION & 32'h00002030);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_214 = 32'h00002030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_216 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_217) == 32'h00000024);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_218 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_219) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_229 = (decode_INSTRUCTION & 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_230 = 32'h0;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_235 = 32'h00004014;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_238 = (decode_INSTRUCTION & 32'h00006014);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_239 = 32'h00002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_242 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_243) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_244 = {(_zz__zz_decode_CfuPlugin_CFU_ENABLE_245 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_246),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_247,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_249,_zz__zz_decode_CfuPlugin_CFU_ENABLE_252}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_257 = {_zz_decode_CfuPlugin_CFU_ENABLE_5,_zz_decode_CfuPlugin_CFU_ENABLE_4};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_259 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_260,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_262,_zz__zz_decode_CfuPlugin_CFU_ENABLE_265}});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_268 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_269,_zz__zz_decode_CfuPlugin_CFU_ENABLE_272});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_274 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_275),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_276,_zz__zz_decode_CfuPlugin_CFU_ENABLE_277}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_217 = 32'h00002024;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_219 = 32'h00000064;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_243 = 32'h00000044;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_245 = (decode_INSTRUCTION & 32'h00000038);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_246 = 32'h00000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_247 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_248) == 32'h00004000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_249 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_250 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_251);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_252 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_253,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_254,_zz__zz_decode_CfuPlugin_CFU_ENABLE_255}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_260 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_261) == 32'h00000040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_262 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_263 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_264);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_265 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_266 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_267);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_269 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_270 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_271);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_272 = {_zz_decode_CfuPlugin_CFU_ENABLE_2,_zz__zz_decode_CfuPlugin_CFU_ENABLE_273};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_275 = {_zz_decode_CfuPlugin_CFU_ENABLE_3,_zz_decode_CfuPlugin_CFU_ENABLE_2};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_276 = (|_zz_decode_CfuPlugin_CFU_ENABLE_1);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_277 = (|_zz_decode_CfuPlugin_CFU_ENABLE_1);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_248 = 32'h00004050;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_250 = (decode_INSTRUCTION & 32'h00002050);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_251 = 32'h00002000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_253 = ((decode_INSTRUCTION & 32'h00006024) == 32'h00002020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_254 = ((decode_INSTRUCTION & 32'h00005024) == 32'h00001020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_255 = ((decode_INSTRUCTION & 32'h90000034) == 32'h90000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_261 = 32'h00000044;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_263 = (decode_INSTRUCTION & 32'h00002014);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_264 = 32'h00002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_266 = (decode_INSTRUCTION & 32'h40000034);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_267 = 32'h40000030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_270 = (decode_INSTRUCTION & 32'h00000048);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_271 = 32'h00000048;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_273 = ((decode_INSTRUCTION & 32'h00002014) == 32'h00000004);
  assign _zz_CsrPlugin_csrMapping_readDataInit_17 = 32'h0;
  assign _zz_CsrPlugin_csrMapping_readDataInit_18 = 32'h0;
  assign _zz_CsrPlugin_csrMapping_readDataInit_19 = 32'h0;
  always @(posedge io_systemClk) begin
    if(_zz_decode_RegFilePlugin_rs1Data) begin
      RegFilePlugin_regFile_spinal_port0 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress1];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_decode_RegFilePlugin_rs2Data) begin
      RegFilePlugin_regFile_spinal_port1 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress2];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      RegFilePlugin_regFile[lastStageRegFileWrite_payload_address] <= lastStageRegFileWrite_payload_data;
    end
  end

  InstructionCache IBusCachedPlugin_cache (
    .io_flush                              (IBusCachedPlugin_cache_io_flush                           ), //i
    .io_cpu_prefetch_isValid               (IBusCachedPlugin_cache_io_cpu_prefetch_isValid            ), //i
    .io_cpu_prefetch_haltIt                (IBusCachedPlugin_cache_io_cpu_prefetch_haltIt             ), //o
    .io_cpu_prefetch_pc                    (IBusCachedPlugin_iBusRsp_stages_0_input_payload[31:0]     ), //i
    .io_cpu_fetch_isValid                  (IBusCachedPlugin_cache_io_cpu_fetch_isValid               ), //i
    .io_cpu_fetch_isStuck                  (IBusCachedPlugin_cache_io_cpu_fetch_isStuck               ), //i
    .io_cpu_fetch_isRemoved                (IBusCachedPlugin_cache_io_cpu_fetch_isRemoved             ), //i
    .io_cpu_fetch_pc                       (IBusCachedPlugin_iBusRsp_stages_1_input_payload[31:0]     ), //i
    .io_cpu_fetch_data                     (IBusCachedPlugin_cache_io_cpu_fetch_data[31:0]            ), //o
    .io_cpu_fetch_mmuRsp_physicalAddress   (IBusCachedPlugin_mmuBus_rsp_physicalAddress[31:0]         ), //i
    .io_cpu_fetch_mmuRsp_isIoAccess        (IBusCachedPlugin_mmuBus_rsp_isIoAccess                    ), //i
    .io_cpu_fetch_mmuRsp_isPaging          (IBusCachedPlugin_mmuBus_rsp_isPaging                      ), //i
    .io_cpu_fetch_mmuRsp_allowRead         (IBusCachedPlugin_mmuBus_rsp_allowRead                     ), //i
    .io_cpu_fetch_mmuRsp_allowWrite        (IBusCachedPlugin_mmuBus_rsp_allowWrite                    ), //i
    .io_cpu_fetch_mmuRsp_allowExecute      (IBusCachedPlugin_mmuBus_rsp_allowExecute                  ), //i
    .io_cpu_fetch_mmuRsp_exception         (IBusCachedPlugin_mmuBus_rsp_exception                     ), //i
    .io_cpu_fetch_mmuRsp_refilling         (IBusCachedPlugin_mmuBus_rsp_refilling                     ), //i
    .io_cpu_fetch_mmuRsp_bypassTranslation (IBusCachedPlugin_mmuBus_rsp_bypassTranslation             ), //i
    .io_cpu_fetch_physicalAddress          (IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress[31:0] ), //o
    .io_cpu_decode_isValid                 (IBusCachedPlugin_cache_io_cpu_decode_isValid              ), //i
    .io_cpu_decode_isStuck                 (IBusCachedPlugin_cache_io_cpu_decode_isStuck              ), //i
    .io_cpu_decode_pc                      (IBusCachedPlugin_iBusRsp_stages_2_input_payload[31:0]     ), //i
    .io_cpu_decode_physicalAddress         (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31:0]), //o
    .io_cpu_decode_data                    (IBusCachedPlugin_cache_io_cpu_decode_data[31:0]           ), //o
    .io_cpu_decode_cacheMiss               (IBusCachedPlugin_cache_io_cpu_decode_cacheMiss            ), //o
    .io_cpu_decode_error                   (IBusCachedPlugin_cache_io_cpu_decode_error                ), //o
    .io_cpu_decode_mmuRefilling            (IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling         ), //o
    .io_cpu_decode_mmuException            (IBusCachedPlugin_cache_io_cpu_decode_mmuException         ), //o
    .io_cpu_decode_isUser                  (IBusCachedPlugin_cache_io_cpu_decode_isUser               ), //i
    .io_cpu_fill_valid                     (IBusCachedPlugin_cache_io_cpu_fill_valid                  ), //i
    .io_cpu_fill_payload                   (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31:0]), //i
    .io_mem_cmd_valid                      (IBusCachedPlugin_cache_io_mem_cmd_valid                   ), //o
    .io_mem_cmd_ready                      (iBus_cmd_ready                                            ), //i
    .io_mem_cmd_payload_address            (IBusCachedPlugin_cache_io_mem_cmd_payload_address[31:0]   ), //o
    .io_mem_cmd_payload_size               (IBusCachedPlugin_cache_io_mem_cmd_payload_size[2:0]       ), //o
    .io_mem_rsp_valid                      (iBus_rsp_valid                                            ), //i
    .io_mem_rsp_payload_data               (iBus_rsp_payload_data[63:0]                               ), //i
    .io_mem_rsp_payload_error              (iBus_rsp_payload_error                                    ), //i
    .io_systemClk                          (io_systemClk                                              ), //i
    .systemCd_logic_outputReset            (systemCd_logic_outputReset                                )  //i
  );
  DataCache dataCache_2 (
    .io_cpu_execute_isValid                 (dataCache_2_io_cpu_execute_isValid               ), //i
    .io_cpu_execute_address                 (dataCache_2_io_cpu_execute_address[31:0]         ), //i
    .io_cpu_execute_haltIt                  (dataCache_2_io_cpu_execute_haltIt                ), //o
    .io_cpu_execute_args_wr                 (execute_MEMORY_WR                                ), //i
    .io_cpu_execute_args_size               (execute_DBusCachedPlugin_size[1:0]               ), //i
    .io_cpu_execute_args_isLrsc             (dataCache_2_io_cpu_execute_args_isLrsc           ), //i
    .io_cpu_execute_args_isAmo              (execute_MEMORY_AMO                               ), //i
    .io_cpu_execute_args_amoCtrl_swap       (dataCache_2_io_cpu_execute_args_amoCtrl_swap     ), //i
    .io_cpu_execute_args_amoCtrl_alu        (dataCache_2_io_cpu_execute_args_amoCtrl_alu[2:0] ), //i
    .io_cpu_execute_args_totalyConsistent   (execute_MEMORY_FORCE_CONSTISTENCY                ), //i
    .io_cpu_execute_refilling               (dataCache_2_io_cpu_execute_refilling             ), //o
    .io_cpu_memory_isValid                  (dataCache_2_io_cpu_memory_isValid                ), //i
    .io_cpu_memory_isStuck                  (memory_arbitration_isStuck                       ), //i
    .io_cpu_memory_isWrite                  (dataCache_2_io_cpu_memory_isWrite                ), //o
    .io_cpu_memory_address                  (memory_MEMORY_VIRTUAL_ADDRESS[31:0]              ), //i
    .io_cpu_memory_mmuRsp_physicalAddress   (DBusCachedPlugin_mmuBus_rsp_physicalAddress[31:0]), //i
    .io_cpu_memory_mmuRsp_isIoAccess        (dataCache_2_io_cpu_memory_mmuRsp_isIoAccess      ), //i
    .io_cpu_memory_mmuRsp_isPaging          (DBusCachedPlugin_mmuBus_rsp_isPaging             ), //i
    .io_cpu_memory_mmuRsp_allowRead         (DBusCachedPlugin_mmuBus_rsp_allowRead            ), //i
    .io_cpu_memory_mmuRsp_allowWrite        (DBusCachedPlugin_mmuBus_rsp_allowWrite           ), //i
    .io_cpu_memory_mmuRsp_allowExecute      (DBusCachedPlugin_mmuBus_rsp_allowExecute         ), //i
    .io_cpu_memory_mmuRsp_exception         (DBusCachedPlugin_mmuBus_rsp_exception            ), //i
    .io_cpu_memory_mmuRsp_refilling         (DBusCachedPlugin_mmuBus_rsp_refilling            ), //i
    .io_cpu_memory_mmuRsp_bypassTranslation (DBusCachedPlugin_mmuBus_rsp_bypassTranslation    ), //i
    .io_cpu_writeBack_isValid               (dataCache_2_io_cpu_writeBack_isValid             ), //i
    .io_cpu_writeBack_isStuck               (writeBack_arbitration_isStuck                    ), //i
    .io_cpu_writeBack_isFiring              (writeBack_arbitration_isFiring                   ), //i
    .io_cpu_writeBack_isUser                (dataCache_2_io_cpu_writeBack_isUser              ), //i
    .io_cpu_writeBack_haltIt                (dataCache_2_io_cpu_writeBack_haltIt              ), //o
    .io_cpu_writeBack_isWrite               (dataCache_2_io_cpu_writeBack_isWrite             ), //o
    .io_cpu_writeBack_storeData             (dataCache_2_io_cpu_writeBack_storeData[63:0]     ), //i
    .io_cpu_writeBack_data                  (dataCache_2_io_cpu_writeBack_data[63:0]          ), //o
    .io_cpu_writeBack_address               (dataCache_2_io_cpu_writeBack_address[31:0]       ), //i
    .io_cpu_writeBack_mmuException          (dataCache_2_io_cpu_writeBack_mmuException        ), //o
    .io_cpu_writeBack_unalignedAccess       (dataCache_2_io_cpu_writeBack_unalignedAccess     ), //o
    .io_cpu_writeBack_accessError           (dataCache_2_io_cpu_writeBack_accessError         ), //o
    .io_cpu_writeBack_keepMemRspData        (dataCache_2_io_cpu_writeBack_keepMemRspData      ), //o
    .io_cpu_writeBack_fence_SW              (dataCache_2_io_cpu_writeBack_fence_SW            ), //i
    .io_cpu_writeBack_fence_SR              (dataCache_2_io_cpu_writeBack_fence_SR            ), //i
    .io_cpu_writeBack_fence_SO              (dataCache_2_io_cpu_writeBack_fence_SO            ), //i
    .io_cpu_writeBack_fence_SI              (dataCache_2_io_cpu_writeBack_fence_SI            ), //i
    .io_cpu_writeBack_fence_PW              (dataCache_2_io_cpu_writeBack_fence_PW            ), //i
    .io_cpu_writeBack_fence_PR              (dataCache_2_io_cpu_writeBack_fence_PR            ), //i
    .io_cpu_writeBack_fence_PO              (dataCache_2_io_cpu_writeBack_fence_PO            ), //i
    .io_cpu_writeBack_fence_PI              (dataCache_2_io_cpu_writeBack_fence_PI            ), //i
    .io_cpu_writeBack_fence_FM              (dataCache_2_io_cpu_writeBack_fence_FM[3:0]       ), //i
    .io_cpu_writeBack_exclusiveOk           (dataCache_2_io_cpu_writeBack_exclusiveOk         ), //o
    .io_cpu_redo                            (dataCache_2_io_cpu_redo                          ), //o
    .io_cpu_flush_valid                     (dataCache_2_io_cpu_flush_valid                   ), //i
    .io_cpu_flush_ready                     (dataCache_2_io_cpu_flush_ready                   ), //o
    .io_cpu_flush_payload_singleLine        (dataCache_2_io_cpu_flush_payload_singleLine      ), //i
    .io_cpu_flush_payload_lineId            (dataCache_2_io_cpu_flush_payload_lineId[5:0]     ), //i
    .io_cpu_writesPending                   (dataCache_2_io_cpu_writesPending                 ), //o
    .io_mem_cmd_valid                       (dataCache_2_io_mem_cmd_valid                     ), //o
    .io_mem_cmd_ready                       (dataCache_2_io_mem_cmd_rValidN                   ), //i
    .io_mem_cmd_payload_wr                  (dataCache_2_io_mem_cmd_payload_wr                ), //o
    .io_mem_cmd_payload_uncached            (dataCache_2_io_mem_cmd_payload_uncached          ), //o
    .io_mem_cmd_payload_address             (dataCache_2_io_mem_cmd_payload_address[31:0]     ), //o
    .io_mem_cmd_payload_data                (dataCache_2_io_mem_cmd_payload_data[63:0]        ), //o
    .io_mem_cmd_payload_mask                (dataCache_2_io_mem_cmd_payload_mask[7:0]         ), //o
    .io_mem_cmd_payload_size                (dataCache_2_io_mem_cmd_payload_size[2:0]         ), //o
    .io_mem_cmd_payload_exclusive           (dataCache_2_io_mem_cmd_payload_exclusive         ), //o
    .io_mem_cmd_payload_last                (dataCache_2_io_mem_cmd_payload_last              ), //o
    .io_mem_rsp_valid                       (dBus_rsp_valid_regNext                           ), //i
    .io_mem_rsp_payload_aggregated          (dBus_rsp_payload_aggregated_regNext[3:0]         ), //i
    .io_mem_rsp_payload_last                (dBus_rsp_payload_last_regNext                    ), //i
    .io_mem_rsp_payload_data                (dBus_rsp_payload_data_regNextWhen[63:0]          ), //i
    .io_mem_rsp_payload_error               (dBus_rsp_payload_error_regNext                   ), //i
    .io_mem_rsp_payload_exclusive           (dBus_rsp_payload_exclusive_regNext               ), //i
    .io_mem_inv_valid                       (dBus_inv_valid                                   ), //i
    .io_mem_inv_ready                       (dataCache_2_io_mem_inv_ready                     ), //o
    .io_mem_inv_payload_last                (dBus_inv_payload_last                            ), //i
    .io_mem_inv_payload_fragment_enable     (dBus_inv_payload_fragment_enable                 ), //i
    .io_mem_inv_payload_fragment_address    (dBus_inv_payload_fragment_address[31:0]          ), //i
    .io_mem_ack_valid                       (dataCache_2_io_mem_ack_valid                     ), //o
    .io_mem_ack_ready                       (dBus_ack_ready                                   ), //i
    .io_mem_ack_payload_last                (dataCache_2_io_mem_ack_payload_last              ), //o
    .io_mem_ack_payload_fragment_hit        (dataCache_2_io_mem_ack_payload_fragment_hit      ), //o
    .io_mem_sync_valid                      (dBus_sync_valid                                  ), //i
    .io_mem_sync_ready                      (dataCache_2_io_mem_sync_ready                    ), //o
    .io_mem_sync_payload_aggregated         (dBus_sync_payload_aggregated[3:0]                ), //i
    .io_systemClk                           (io_systemClk                                     ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                       )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC systemCd_logic_outputReset_buffercc (
    .io_dataIn                  (systemCd_logic_outputReset                    ), //i
    .io_dataOut                 (systemCd_logic_outputReset_buffercc_io_dataOut), //o
    .io_systemClk               (io_systemClk                                  ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                    )  //i
  );
  EfxCPUSp1 EfxCPUSp1_inst (
    .src1    (execute_SRC1[31:0]           ), //i
    .src2    (execute_SRC2[31:0]           ), //i
    .bitCtrl (execute_ALU_BITWISE_CTRL[1:0]), //i
    .ctrl    (execute_ALU_CTRL[1:0]        ), //i
    .less    (execute_SRC_LESS             ), //i
    .addSub  (execute_SRC_ADD_SUB[31:0]    ), //i
    .result  (EfxCPUSp1_inst_result[31:0]  )  //o
  );
  EfxCPUSp2 EfxCPUSp2_inst (
    .ctrl   (execute_SHIFT_CTRL[1:0]    ), //i
    .src1   (execute_SRC1[31:0]         ), //i
    .src2   (execute_SRC2[31:0]         ), //i
    .result (EfxCPUSp2_inst_result[31:0])  //o
  );
  always @(*) begin
    case(_zz_IBusCachedPlugin_jump_pcLoad_payload_5)
      2'b00 : _zz_IBusCachedPlugin_jump_pcLoad_payload_4 = DBusCachedPlugin_redoBranch_payload;
      2'b01 : _zz_IBusCachedPlugin_jump_pcLoad_payload_4 = CsrPlugin_jumpInterface_payload;
      default : _zz_IBusCachedPlugin_jump_pcLoad_payload_4 = BranchPlugin_jumpInterface_payload;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_1)
      3'b000 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_0;
      3'b001 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_1;
      3'b010 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_2;
      3'b011 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_3;
      3'b100 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_4;
      3'b101 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_5;
      3'b110 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_6;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_7;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_3)
      2'b00 : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_1;
      2'b01 : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_3;
      2'b10 : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_5;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_7;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_5)
      1'b0 : _zz_writeBack_DBusCachedPlugin_rspShifted_4 = writeBack_DBusCachedPlugin_rspSplits_2;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted_4 = writeBack_DBusCachedPlugin_rspSplits_6;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_7)
      1'b0 : _zz_writeBack_DBusCachedPlugin_rspShifted_6 = writeBack_DBusCachedPlugin_rspSplits_3;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted_6 = writeBack_DBusCachedPlugin_rspSplits_7;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(_zz_execute_to_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_execute_to_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_execute_to_memory_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : decode_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : decode_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : decode_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : decode_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : decode_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL_1)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : decode_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : decode_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : decode_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1)
      Input2Kind_RS : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string = "IMM_I";
      default : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(memory_FPU_OPCODE)
      FpuOpcode_LOAD : memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : memory_FPU_OPCODE_string = "FCVT_X_X";
      default : memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_memory_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_memory_to_writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_memory_to_writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_memory_to_writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_memory_to_writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_memory_to_writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_memory_to_writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_memory_to_writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_memory_to_writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_memory_to_writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_memory_to_writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_memory_to_writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_memory_to_writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_memory_to_writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_memory_to_writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_memory_to_writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_memory_to_writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_memory_to_writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_FPU_OPCODE)
      FpuOpcode_LOAD : execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : execute_FPU_OPCODE_string = "FCVT_X_X";
      default : execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_execute_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_execute_to_memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_execute_to_memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_execute_to_memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_execute_to_memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_execute_to_memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_execute_to_memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_execute_to_memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_execute_to_memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_execute_to_memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_execute_to_memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_execute_to_memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_execute_to_memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_execute_to_memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_execute_to_memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_execute_to_memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_execute_to_memory_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_execute_to_memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_execute_to_memory_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_execute_to_memory_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_execute_to_memory_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_execute_to_memory_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_execute_to_memory_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_execute_to_memory_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_execute_to_memory_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_execute_to_memory_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_execute_to_memory_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_execute_to_memory_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_execute_to_memory_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_execute_to_memory_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_execute_to_memory_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_execute_to_memory_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_execute_to_memory_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_execute_to_memory_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_execute_to_memory_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_decode_to_execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_to_execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_to_execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_to_execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_to_execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_to_execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_to_execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_to_execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_to_execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_to_execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_to_execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_to_execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_to_execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_to_execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_to_execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_to_execute_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_decode_to_execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_decode_to_execute_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_to_execute_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_to_execute_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_to_execute_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_to_execute_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_to_execute_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_to_execute_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_to_execute_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_to_execute_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_to_execute_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_to_execute_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_to_execute_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_to_execute_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_to_execute_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_to_execute_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_to_execute_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_decode_to_execute_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_BRANCH_CTRL)
      BranchCtrlEnum_INC : decode_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : decode_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : decode_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : decode_BRANCH_CTRL_string = "JALR";
      default : decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_decode_to_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_to_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_to_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL_1)
      BranchCtrlEnum_INC : _zz_decode_to_execute_BRANCH_CTRL_1_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_to_execute_BRANCH_CTRL_1_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_memory_to_writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_memory_to_writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_memory_to_writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_memory_to_writeBack_ENV_CTRL_string = "EBREAK";
      default : _zz_memory_to_writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_memory_to_writeBack_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_memory_to_writeBack_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_memory_to_writeBack_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_memory_to_writeBack_ENV_CTRL_1_string = "EBREAK";
      default : _zz_memory_to_writeBack_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_execute_to_memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_execute_to_memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_execute_to_memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_execute_to_memory_ENV_CTRL_string = "EBREAK";
      default : _zz_execute_to_memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_execute_to_memory_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_execute_to_memory_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_execute_to_memory_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_execute_to_memory_ENV_CTRL_1_string = "EBREAK";
      default : _zz_execute_to_memory_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_ENV_CTRL)
      EnvCtrlEnum_NONE : decode_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : decode_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : decode_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : decode_ENV_CTRL_string = "EBREAK";
      default : decode_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_ENV_CTRL_string = "EBREAK";
      default : _zz_decode_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_decode_to_execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_to_execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_to_execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_to_execute_ENV_CTRL_string = "EBREAK";
      default : _zz_decode_to_execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_decode_to_execute_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_to_execute_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_to_execute_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_to_execute_ENV_CTRL_1_string = "EBREAK";
      default : _zz_decode_to_execute_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : decode_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : decode_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : decode_ALU_CTRL_string = "BITWISE ";
      default : decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL_1)
      AluCtrlEnum_ADD_SUB : _zz_decode_to_execute_ALU_CTRL_1_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_to_execute_ALU_CTRL_1_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_to_execute_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : memory_SHIFT_CTRL_string = "SRA_1    ";
      default : memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : execute_SHIFT_CTRL_string = "SRA_1    ";
      default : execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : execute_ALU_CTRL_string = "BITWISE ";
      default : execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_FPU_FORMAT)
      FpuFormat_FLOAT : decode_FPU_FORMAT_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_FPU_FORMAT_string = "DOUBLE";
      default : decode_FPU_FORMAT_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_FORMAT)
      FpuFormat_FLOAT : _zz_decode_FPU_FORMAT_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_decode_FPU_FORMAT_string = "DOUBLE";
      default : _zz_decode_FPU_FORMAT_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_FPU_OPCODE)
      FpuOpcode_LOAD : decode_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : decode_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : decode_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : decode_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : decode_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : decode_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : decode_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : decode_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : decode_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : decode_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : decode_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : decode_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : decode_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : decode_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : decode_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : decode_FPU_OPCODE_string = "FCVT_X_X";
      default : decode_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_decode_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_decode_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : execute_BRANCH_CTRL_string = "JALR";
      default : execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(memory_ENV_CTRL)
      EnvCtrlEnum_NONE : memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : memory_ENV_CTRL_string = "EBREAK";
      default : memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_memory_ENV_CTRL_string = "EBREAK";
      default : _zz_memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ENV_CTRL)
      EnvCtrlEnum_NONE : execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : execute_ENV_CTRL_string = "EBREAK";
      default : execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_execute_ENV_CTRL_string = "EBREAK";
      default : _zz_execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : writeBack_ENV_CTRL_string = "EBREAK";
      default : writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_writeBack_ENV_CTRL_string = "EBREAK";
      default : _zz_writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_SRC2_CTRL)
      Src2CtrlEnum_RS : decode_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : decode_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : decode_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : decode_SRC2_CTRL_string = "PC ";
      default : decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_string = "PC ";
      default : _zz_decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_SRC1_CTRL)
      Src1CtrlEnum_RS : decode_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : decode_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : decode_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : decode_SRC1_CTRL_string = "URS1        ";
      default : decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_1)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1)
      Input2Kind_RS : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string = "IMM_I";
      default : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_FORMAT_1)
      FpuFormat_FLOAT : _zz_decode_FPU_FORMAT_1_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_decode_FPU_FORMAT_1_string = "DOUBLE";
      default : _zz_decode_FPU_FORMAT_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_decode_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_decode_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_1)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_1_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_1_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_1_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_ENV_CTRL_1_string = "EBREAK";
      default : _zz_decode_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_1)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_1_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_1_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_1_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_1_string = "PC ";
      default : _zz_decode_SRC2_CTRL_1_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_1)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_1_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_1_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_1)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_1_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_1_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_1_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_1_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_1_string = "????????????";
    endcase
  end
  always @(*) begin
    case(debugBus_dmToHart_payload_op)
      DebugDmToHartOp_DATA : debugBus_dmToHart_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : debugBus_dmToHart_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : debugBus_dmToHart_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : debugBus_dmToHart_payload_op_string = "REG_READ ";
      default : debugBus_dmToHart_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_cmd_payload_opcode)
      FpuOpcode_LOAD : FpuPlugin_port_cmd_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_cmd_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_cmd_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_cmd_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_cmd_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_cmd_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_cmd_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_cmd_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_cmd_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_cmd_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_cmd_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_cmd_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_cmd_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_cmd_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_cmd_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_cmd_payload_opcode_string = "FCVT_X_X";
      default : FpuPlugin_port_cmd_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_cmd_payload_format)
      FpuFormat_FLOAT : FpuPlugin_port_cmd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : FpuPlugin_port_cmd_payload_format_string = "DOUBLE";
      default : FpuPlugin_port_cmd_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_cmd_payload_roundMode)
      FpuRoundMode_RNE : FpuPlugin_port_cmd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuPlugin_port_cmd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuPlugin_port_cmd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuPlugin_port_cmd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuPlugin_port_cmd_payload_roundMode_string = "RMM";
      default : FpuPlugin_port_cmd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_commit_payload_opcode)
      FpuOpcode_LOAD : FpuPlugin_port_commit_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_commit_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_commit_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_commit_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_commit_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_commit_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_commit_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_commit_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_commit_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_commit_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_commit_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_commit_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_commit_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_commit_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_commit_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_commit_payload_opcode_string = "FCVT_X_X";
      default : FpuPlugin_port_commit_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_2)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_2_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_2_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_2_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_2_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_2_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_2)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_2_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_2_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_2_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_2)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_2_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_2_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_2_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_2_string = "PC ";
      default : _zz_decode_SRC2_CTRL_2_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_2)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_2_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_2_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_2_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_ENV_CTRL_2_string = "EBREAK";
      default : _zz_decode_ENV_CTRL_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_2)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_2_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_2_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_2_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_2_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_OPCODE_2)
      FpuOpcode_LOAD : _zz_decode_FPU_OPCODE_2_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_FPU_OPCODE_2_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_FPU_OPCODE_2_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_FPU_OPCODE_2_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_FPU_OPCODE_2_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_FPU_OPCODE_2_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_FPU_OPCODE_2_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_FPU_OPCODE_2_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_FPU_OPCODE_2_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_FPU_OPCODE_2_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_FPU_OPCODE_2_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_FPU_OPCODE_2_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_FPU_OPCODE_2_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_FPU_OPCODE_2_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_FPU_OPCODE_2_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_FPU_OPCODE_2_string = "FCVT_X_X";
      default : _zz_decode_FPU_OPCODE_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_FORMAT_2)
      FpuFormat_FLOAT : _zz_decode_FPU_FORMAT_2_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_decode_FPU_FORMAT_2_string = "DOUBLE";
      default : _zz_decode_FPU_FORMAT_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2)
      Input2Kind_RS : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string = "IMM_I";
      default : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_2)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_2)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_2_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_2_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_2_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_2_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_2_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_cmd_payload_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_cmd_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_cmd_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_cmd_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_cmd_payload_op_string = "REG_READ ";
      default : CsrPlugin_inject_cmd_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_cmd_toStream_payload_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_cmd_toStream_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_cmd_toStream_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_cmd_toStream_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_cmd_toStream_payload_op_string = "REG_READ ";
      default : CsrPlugin_inject_cmd_toStream_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_buffer_payload_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_buffer_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_buffer_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_buffer_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_buffer_payload_op_string = "REG_READ ";
      default : CsrPlugin_inject_buffer_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_cmd_toStream_rData_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_cmd_toStream_rData_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_cmd_toStream_rData_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_cmd_toStream_rData_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_cmd_toStream_rData_op_string = "REG_READ ";
      default : CsrPlugin_inject_cmd_toStream_rData_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_BOOT : CsrPlugin_dcsr_stepLogic_stateReg_string = "BOOT  ";
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : CsrPlugin_dcsr_stepLogic_stateReg_string = "IDLE  ";
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : CsrPlugin_dcsr_stepLogic_stateReg_string = "SINGLE";
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : CsrPlugin_dcsr_stepLogic_stateReg_string = "WAIT_1";
      default : CsrPlugin_dcsr_stepLogic_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_dcsr_stepLogic_stateNext)
      CsrPlugin_dcsr_stepLogic_enumDef_BOOT : CsrPlugin_dcsr_stepLogic_stateNext_string = "BOOT  ";
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : CsrPlugin_dcsr_stepLogic_stateNext_string = "IDLE  ";
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : CsrPlugin_dcsr_stepLogic_stateNext_string = "SINGLE";
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : CsrPlugin_dcsr_stepLogic_stateNext_string = "WAIT_1";
      default : CsrPlugin_dcsr_stepLogic_stateNext_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPlugin_port_cmd_payload_roundMode)
      FpuRoundMode_RNE : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RMM";
      default : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPlugin_port_cmd_payload_roundMode_1)
      FpuRoundMode_RNE : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RMM";
      default : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "???";
    endcase
  end
  always @(*) begin
    case(writeBack_FpuPlugin_commit_payload_opcode)
      FpuOpcode_LOAD : writeBack_FpuPlugin_commit_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FpuPlugin_commit_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FpuPlugin_commit_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FpuPlugin_commit_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FpuPlugin_commit_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FpuPlugin_commit_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FpuPlugin_commit_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FpuPlugin_commit_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FpuPlugin_commit_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FpuPlugin_commit_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FpuPlugin_commit_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FpuPlugin_commit_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FpuPlugin_commit_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FpuPlugin_commit_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FpuPlugin_commit_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FpuPlugin_commit_payload_opcode_string = "FCVT_X_X";
      default : writeBack_FpuPlugin_commit_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(writeBack_FpuPlugin_commit_s2mPipe_payload_opcode)
      FpuOpcode_LOAD : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCVT_X_X";
      default : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(writeBack_FpuPlugin_commit_rData_opcode)
      FpuOpcode_LOAD : writeBack_FpuPlugin_commit_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FpuPlugin_commit_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FpuPlugin_commit_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FpuPlugin_commit_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FpuPlugin_commit_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FpuPlugin_commit_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FpuPlugin_commit_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FpuPlugin_commit_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FpuPlugin_commit_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FpuPlugin_commit_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FpuPlugin_commit_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FpuPlugin_commit_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FpuPlugin_commit_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FpuPlugin_commit_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FpuPlugin_commit_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FpuPlugin_commit_rData_opcode_string = "FCVT_X_X";
      default : writeBack_FpuPlugin_commit_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode)
      FpuOpcode_LOAD : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCVT_X_X";
      default : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : decode_to_execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : decode_to_execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : decode_to_execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : decode_to_execute_ENV_CTRL_string = "EBREAK";
      default : decode_to_execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : execute_to_memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : execute_to_memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : execute_to_memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : execute_to_memory_ENV_CTRL_string = "EBREAK";
      default : execute_to_memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(memory_to_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : memory_to_writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : memory_to_writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : memory_to_writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : memory_to_writeBack_ENV_CTRL_string = "EBREAK";
      default : memory_to_writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : decode_to_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : decode_to_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : decode_to_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_FPU_OPCODE)
      FpuOpcode_LOAD : decode_to_execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : decode_to_execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : decode_to_execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : decode_to_execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : decode_to_execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : decode_to_execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : decode_to_execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : decode_to_execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : decode_to_execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : decode_to_execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : decode_to_execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : decode_to_execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : decode_to_execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : decode_to_execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : decode_to_execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : decode_to_execute_FPU_OPCODE_string = "FCVT_X_X";
      default : decode_to_execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_FPU_OPCODE)
      FpuOpcode_LOAD : execute_to_memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : execute_to_memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : execute_to_memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : execute_to_memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : execute_to_memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : execute_to_memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : execute_to_memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : execute_to_memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : execute_to_memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : execute_to_memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : execute_to_memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : execute_to_memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : execute_to_memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : execute_to_memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : execute_to_memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : execute_to_memory_FPU_OPCODE_string = "FCVT_X_X";
      default : execute_to_memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(memory_to_writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : memory_to_writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : memory_to_writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : memory_to_writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : memory_to_writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : memory_to_writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : memory_to_writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : memory_to_writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : memory_to_writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : memory_to_writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : memory_to_writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : memory_to_writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : memory_to_writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : memory_to_writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : memory_to_writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : memory_to_writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : memory_to_writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : memory_to_writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : execute_to_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : execute_to_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : execute_to_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : execute_to_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : execute_to_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_BOOT : FpuPlugin_stateReg_string = "BOOT  ";
      FpuPlugin_enumDef_IDLE : FpuPlugin_stateReg_string = "IDLE  ";
      FpuPlugin_enumDef_CMD : FpuPlugin_stateReg_string = "CMD   ";
      FpuPlugin_enumDef_RSP : FpuPlugin_stateReg_string = "RSP   ";
      FpuPlugin_enumDef_RSP_0 : FpuPlugin_stateReg_string = "RSP_0 ";
      FpuPlugin_enumDef_RSP_1 : FpuPlugin_stateReg_string = "RSP_1 ";
      FpuPlugin_enumDef_COMMIT : FpuPlugin_stateReg_string = "COMMIT";
      FpuPlugin_enumDef_DONE : FpuPlugin_stateReg_string = "DONE  ";
      default : FpuPlugin_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_stateNext)
      FpuPlugin_enumDef_BOOT : FpuPlugin_stateNext_string = "BOOT  ";
      FpuPlugin_enumDef_IDLE : FpuPlugin_stateNext_string = "IDLE  ";
      FpuPlugin_enumDef_CMD : FpuPlugin_stateNext_string = "CMD   ";
      FpuPlugin_enumDef_RSP : FpuPlugin_stateNext_string = "RSP   ";
      FpuPlugin_enumDef_RSP_0 : FpuPlugin_stateNext_string = "RSP_0 ";
      FpuPlugin_enumDef_RSP_1 : FpuPlugin_stateNext_string = "RSP_1 ";
      FpuPlugin_enumDef_COMMIT : FpuPlugin_stateNext_string = "COMMIT";
      FpuPlugin_enumDef_DONE : FpuPlugin_stateNext_string = "DONE  ";
      default : FpuPlugin_stateNext_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPlugin_port_cmd_payload_format)
      FpuFormat_FLOAT : _zz_FpuPlugin_port_cmd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_FpuPlugin_port_cmd_payload_format_string = "DOUBLE";
      default : _zz_FpuPlugin_port_cmd_payload_format_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    CsrPlugin_running_aheadValue = CsrPlugin_running;
    if(when_CsrPlugin_l1534) begin
      if(!when_CsrPlugin_l1542) begin
        CsrPlugin_running_aheadValue = 1'b0;
      end
    end
    if(CsrPlugin_doResume) begin
      CsrPlugin_running_aheadValue = 1'b1;
    end
  end

  assign writeBack_MEMORY_LOAD_DATA = writeBack_DBusCachedPlugin_rspShifted;
  assign memory_MUL_LOW = ($signed(_zz_memory_MUL_LOW) + $signed(_zz_memory_MUL_LOW_6));
  assign execute_SHIFT_RIGHT = EfxCPUSp2_inst_result;
  assign execute_REGFILE_WRITE_DATA = EfxCPUSp1_inst_result;
  assign memory_CfuPlugin_CFU_IN_FLIGHT = execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
  assign execute_CfuPlugin_CFU_IN_FLIGHT = ((execute_CfuPlugin_schedule || execute_CfuPlugin_hold) || execute_CfuPlugin_fired);
  assign memory_MUL_HH = execute_to_memory_MUL_HH;
  assign execute_MUL_HH = execute_MulPlugin_withOuputBuffer_mul_hh;
  assign execute_MUL_HL = execute_MulPlugin_withOuputBuffer_mul_hl;
  assign execute_MUL_LH = execute_MulPlugin_withOuputBuffer_mul_lh;
  assign execute_MUL_LL = execute_MulPlugin_withOuputBuffer_mul_ll;
  assign execute_BRANCH_CALC = {execute_BranchPlugin_branchAdder[31 : 1],1'b0};
  assign execute_BRANCH_DO = _zz_execute_BRANCH_DO_1;
  assign execute_MEMORY_VIRTUAL_ADDRESS = dataCache_2_io_cpu_execute_address;
  assign execute_MEMORY_STORE_DATA_RF = _zz_execute_MEMORY_STORE_DATA_RF;
  assign memory_FPU_COMMIT_LOAD = execute_to_memory_FPU_COMMIT_LOAD;
  assign execute_FPU_COMMIT_LOAD = decode_to_execute_FPU_COMMIT_LOAD;
  assign decode_FPU_COMMIT_LOAD = (decode_FPU_OPCODE == FpuOpcode_LOAD);
  assign memory_FPU_FORKED = execute_to_memory_FPU_FORKED;
  assign execute_FPU_FORKED = decode_to_execute_FPU_FORKED;
  assign decode_FPU_FORKED = (decode_FpuPlugin_forked || (FpuPlugin_port_cmd_fire && (! _zz_decode_FPU_FORKED)));
  assign decode_CSR_READ_OPCODE = (decode_INSTRUCTION[13 : 7] != 7'h20);
  assign decode_CSR_WRITE_OPCODE = (! (((decode_INSTRUCTION[14 : 13] == 2'b01) && (decode_INSTRUCTION[19 : 15] == 5'h0)) || ((decode_INSTRUCTION[14 : 13] == 2'b11) && (decode_INSTRUCTION[19 : 15] == 5'h0))));
  assign decode_SRC2 = _zz_decode_SRC2_4;
  assign decode_SRC1 = _zz_decode_SRC1;
  assign decode_SRC2_FORCE_ZERO = (decode_SRC_ADD_ZERO && (! decode_SRC_USE_SUB_LESS));
  assign memory_RS1 = execute_to_memory_RS1;
  assign _zz_execute_to_memory_SHIFT_CTRL = _zz_execute_to_memory_SHIFT_CTRL_1;
  assign decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL = _zz_decode_to_execute_SHIFT_CTRL_1;
  assign decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL = _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  assign decode_CfuPlugin_CFU_INPUT_2_KIND = _zz_decode_CfuPlugin_CFU_INPUT_2_KIND;
  assign _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND = _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1;
  assign decode_CfuPlugin_CFU_ENABLE = _zz_decode_CfuPlugin_CFU_ENABLE[42];
  assign memory_FPU_OPCODE = _zz_memory_FPU_OPCODE;
  assign _zz_memory_to_writeBack_FPU_OPCODE = _zz_memory_to_writeBack_FPU_OPCODE_1;
  assign execute_FPU_OPCODE = _zz_execute_FPU_OPCODE;
  assign _zz_execute_to_memory_FPU_OPCODE = _zz_execute_to_memory_FPU_OPCODE_1;
  assign _zz_decode_to_execute_FPU_OPCODE = _zz_decode_to_execute_FPU_OPCODE_1;
  assign memory_FPU_RSP = execute_to_memory_FPU_RSP;
  assign execute_FPU_RSP = decode_to_execute_FPU_RSP;
  assign decode_FPU_RSP = _zz_decode_CfuPlugin_CFU_ENABLE[34];
  assign memory_FPU_COMMIT = execute_to_memory_FPU_COMMIT;
  assign execute_FPU_COMMIT = decode_to_execute_FPU_COMMIT;
  assign decode_FPU_COMMIT = _zz_decode_CfuPlugin_CFU_ENABLE[33];
  assign decode_IS_RS2_SIGNED = _zz_decode_CfuPlugin_CFU_ENABLE[31];
  assign decode_IS_RS1_SIGNED = _zz_decode_CfuPlugin_CFU_ENABLE[30];
  assign decode_IS_DIV = _zz_decode_CfuPlugin_CFU_ENABLE[29];
  assign memory_IS_MUL = execute_to_memory_IS_MUL;
  assign decode_IS_MUL = _zz_decode_CfuPlugin_CFU_ENABLE[28];
  assign decode_SRC_LESS_UNSIGNED = _zz_decode_CfuPlugin_CFU_ENABLE[27];
  assign decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL = _zz_decode_to_execute_BRANCH_CTRL_1;
  assign _zz_memory_to_writeBack_ENV_CTRL = _zz_memory_to_writeBack_ENV_CTRL_1;
  assign _zz_execute_to_memory_ENV_CTRL = _zz_execute_to_memory_ENV_CTRL_1;
  assign decode_ENV_CTRL = _zz_decode_ENV_CTRL;
  assign _zz_decode_to_execute_ENV_CTRL = _zz_decode_to_execute_ENV_CTRL_1;
  assign decode_IS_CSR = _zz_decode_CfuPlugin_CFU_ENABLE[22];
  assign memory_MEMORY_FENCE = execute_to_memory_MEMORY_FENCE;
  assign execute_MEMORY_FENCE = decode_to_execute_MEMORY_FENCE;
  assign decode_MEMORY_FENCE = _zz_decode_CfuPlugin_CFU_ENABLE[21];
  assign decode_MEMORY_MANAGMENT = _zz_decode_CfuPlugin_CFU_ENABLE[20];
  assign memory_MEMORY_AMO = execute_to_memory_MEMORY_AMO;
  assign memory_MEMORY_LRSC = execute_to_memory_MEMORY_LRSC;
  assign execute_HAS_SIDE_EFFECT = decode_to_execute_HAS_SIDE_EFFECT;
  assign decode_HAS_SIDE_EFFECT = _zz_decode_CfuPlugin_CFU_ENABLE[15];
  assign decode_MEMORY_WR = _zz_decode_CfuPlugin_CFU_ENABLE[14];
  assign execute_BYPASSABLE_MEMORY_STAGE = decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  assign decode_BYPASSABLE_MEMORY_STAGE = _zz_decode_CfuPlugin_CFU_ENABLE[13];
  assign decode_BYPASSABLE_EXECUTE_STAGE = _zz_decode_CfuPlugin_CFU_ENABLE[12];
  assign decode_ALU_CTRL = _zz_decode_ALU_CTRL;
  assign _zz_decode_to_execute_ALU_CTRL = _zz_decode_to_execute_ALU_CTRL_1;
  assign decode_MEMORY_FENCE_WR = _zz_decode_CfuPlugin_CFU_ENABLE[1];
  assign decode_MEMORY_FORCE_CONSTISTENCY = _zz_decode_MEMORY_FORCE_CONSTISTENCY;
  assign writeBack_FORMAL_PC_NEXT = memory_to_writeBack_FORMAL_PC_NEXT;
  assign memory_FORMAL_PC_NEXT = execute_to_memory_FORMAL_PC_NEXT;
  assign execute_FORMAL_PC_NEXT = decode_to_execute_FORMAL_PC_NEXT;
  assign decode_FORMAL_PC_NEXT = (decode_PC + _zz_decode_FORMAL_PC_NEXT);
  assign memory_SHIFT_RIGHT = execute_to_memory_SHIFT_RIGHT;
  assign memory_SHIFT_CTRL = _zz_memory_SHIFT_CTRL;
  assign execute_SHIFT_CTRL = _zz_execute_SHIFT_CTRL;
  assign execute_SRC_ADD_SUB = execute_SrcPlugin_addSub;
  assign execute_ALU_CTRL = _zz_execute_ALU_CTRL;
  assign execute_ALU_BITWISE_CTRL = _zz_execute_ALU_BITWISE_CTRL;
  always @(*) begin
    _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT = memory_CfuPlugin_CFU_IN_FLIGHT;
    if(memory_arbitration_isStuck) begin
      _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT = 1'b0;
    end
  end

  always @(*) begin
    _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT = execute_CfuPlugin_CFU_IN_FLIGHT;
    if(execute_arbitration_isStuck) begin
      _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT = 1'b0;
    end
  end

  assign writeBack_CfuPlugin_CFU_IN_FLIGHT = memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
  assign execute_CfuPlugin_CFU_INPUT_2_KIND = _zz_execute_CfuPlugin_CFU_INPUT_2_KIND;
  assign writeBack_HAS_SIDE_EFFECT = memory_to_writeBack_HAS_SIDE_EFFECT;
  assign memory_HAS_SIDE_EFFECT = execute_to_memory_HAS_SIDE_EFFECT;
  assign execute_LEGAL_INSTRUCTION = decode_to_execute_LEGAL_INSTRUCTION;
  always @(*) begin
    execute_CfuPlugin_CFU_ENABLE = decode_to_execute_CfuPlugin_CFU_ENABLE;
    if(when_CfuPlugin_l192) begin
      execute_CfuPlugin_CFU_ENABLE = 1'b0;
    end
  end

  always @(*) begin
    _zz_memory_to_writeBack_FPU_FORKED = memory_FPU_FORKED;
    if(memory_arbitration_isStuck) begin
      _zz_memory_to_writeBack_FPU_FORKED = 1'b0;
    end
  end

  always @(*) begin
    _zz_execute_to_memory_FPU_FORKED = execute_FPU_FORKED;
    if(execute_arbitration_isStuck) begin
      _zz_execute_to_memory_FPU_FORKED = 1'b0;
    end
  end

  always @(*) begin
    _zz_decode_to_execute_FPU_FORKED = decode_FPU_FORKED;
    if(decode_arbitration_isStuck) begin
      _zz_decode_to_execute_FPU_FORKED = 1'b0;
    end
  end

  assign writeBack_FPU_OPCODE = _zz_writeBack_FPU_OPCODE;
  assign writeBack_RS1 = memory_to_writeBack_RS1;
  assign _zz_writeBack_FpuPlugin_commit_payload_value = writeBack_MEMORY_LOAD_DATA;
  assign writeBack_FPU_COMMIT_LOAD = memory_to_writeBack_FPU_COMMIT_LOAD;
  always @(*) begin
    DBusBypass0_cond = 1'b0;
    if(writeBack_FpuPlugin_isRsp) begin
      if(writeBack_arbitration_isValid) begin
        DBusBypass0_cond = 1'b1;
      end
    end
  end

  assign writeBack_FPU_COMMIT = memory_to_writeBack_FPU_COMMIT;
  assign writeBack_FPU_RSP = memory_to_writeBack_FPU_RSP;
  assign writeBack_FPU_FORKED = memory_to_writeBack_FPU_FORKED;
  assign decode_FPU_FORMAT = _zz_decode_FPU_FORMAT;
  assign decode_FPU_ARG = _zz_decode_CfuPlugin_CFU_ENABLE[41 : 40];
  assign decode_FPU_OPCODE = _zz_decode_FPU_OPCODE;
  always @(*) begin
    decode_FPU_ENABLE = _zz_decode_FPU_ENABLE;
    if(when_FpuPlugin_l272) begin
      decode_FPU_ENABLE = 1'b0;
    end
  end

  assign execute_IS_RS1_SIGNED = decode_to_execute_IS_RS1_SIGNED;
  assign execute_IS_DIV = decode_to_execute_IS_DIV;
  assign execute_IS_RS2_SIGNED = decode_to_execute_IS_RS2_SIGNED;
  assign memory_IS_DIV = execute_to_memory_IS_DIV;
  assign writeBack_IS_MUL = memory_to_writeBack_IS_MUL;
  assign writeBack_MUL_HH = memory_to_writeBack_MUL_HH;
  assign writeBack_MUL_LOW = memory_to_writeBack_MUL_LOW;
  assign memory_MUL_HL = execute_to_memory_MUL_HL;
  assign memory_MUL_LH = execute_to_memory_MUL_LH;
  assign memory_MUL_LL = execute_to_memory_MUL_LL;
  assign execute_IS_MUL = decode_to_execute_IS_MUL;
  assign memory_BRANCH_CALC = execute_to_memory_BRANCH_CALC;
  assign memory_BRANCH_DO = execute_to_memory_BRANCH_DO;
  assign execute_PC = decode_to_execute_PC;
  assign execute_BRANCH_CTRL = _zz_execute_BRANCH_CTRL;
  assign execute_SRC_LESS = execute_SrcPlugin_less;
  assign execute_CSR_READ_OPCODE = decode_to_execute_CSR_READ_OPCODE;
  assign execute_CSR_WRITE_OPCODE = decode_to_execute_CSR_WRITE_OPCODE;
  assign execute_IS_CSR = decode_to_execute_IS_CSR;
  assign memory_ENV_CTRL = _zz_memory_ENV_CTRL;
  assign execute_ENV_CTRL = _zz_execute_ENV_CTRL;
  assign writeBack_ENV_CTRL = _zz_writeBack_ENV_CTRL;
  assign decode_RS2_USE = _zz_decode_CfuPlugin_CFU_ENABLE[18];
  assign decode_RS1_USE = _zz_decode_CfuPlugin_CFU_ENABLE[6];
  always @(*) begin
    _zz_decode_RS2 = execute_REGFILE_WRITE_DATA;
    if(when_CsrPlugin_l1731) begin
      _zz_decode_RS2 = CsrPlugin_csrMapping_readDataSignal;
    end
  end

  assign execute_REGFILE_WRITE_VALID = decode_to_execute_REGFILE_WRITE_VALID;
  assign execute_BYPASSABLE_EXECUTE_STAGE = decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  always @(*) begin
    _zz_decode_RS2_1 = memory_REGFILE_WRITE_DATA;
    if(when_MulDivIterativePlugin_l128) begin
      _zz_decode_RS2_1 = memory_MulDivIterativePlugin_div_result;
    end
    if(memory_arbitration_isValid) begin
      case(memory_SHIFT_CTRL)
        ShiftCtrlEnum_SLL_1 : begin
          _zz_decode_RS2_1 = _zz_decode_RS2_3;
        end
        ShiftCtrlEnum_SRL_1, ShiftCtrlEnum_SRA_1 : begin
          _zz_decode_RS2_1 = memory_SHIFT_RIGHT;
        end
        default : begin
        end
      endcase
    end
  end

  assign memory_REGFILE_WRITE_VALID = execute_to_memory_REGFILE_WRITE_VALID;
  assign memory_BYPASSABLE_MEMORY_STAGE = execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  assign writeBack_REGFILE_WRITE_VALID = memory_to_writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    decode_RS2 = decode_RegFilePlugin_rs2Data;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr1Match) begin
        decode_RS2 = HazardSimplePlugin_writeBackBuffer_payload_data;
      end
    end
    if(when_HazardSimplePlugin_l45) begin
      if(when_HazardSimplePlugin_l47) begin
        if(when_HazardSimplePlugin_l51) begin
          decode_RS2 = _zz_decode_RS2_2;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_1) begin
      if(memory_BYPASSABLE_MEMORY_STAGE) begin
        if(when_HazardSimplePlugin_l51_1) begin
          decode_RS2 = _zz_decode_RS2_1;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_2) begin
      if(execute_BYPASSABLE_EXECUTE_STAGE) begin
        if(when_HazardSimplePlugin_l51_2) begin
          decode_RS2 = _zz_decode_RS2;
        end
      end
    end
  end

  always @(*) begin
    decode_RS1 = decode_RegFilePlugin_rs1Data;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr0Match) begin
        decode_RS1 = HazardSimplePlugin_writeBackBuffer_payload_data;
      end
    end
    if(when_HazardSimplePlugin_l45) begin
      if(when_HazardSimplePlugin_l47) begin
        if(when_HazardSimplePlugin_l48) begin
          decode_RS1 = _zz_decode_RS2_2;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_1) begin
      if(memory_BYPASSABLE_MEMORY_STAGE) begin
        if(when_HazardSimplePlugin_l48_1) begin
          decode_RS1 = _zz_decode_RS2_1;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_2) begin
      if(execute_BYPASSABLE_EXECUTE_STAGE) begin
        if(when_HazardSimplePlugin_l48_2) begin
          decode_RS1 = _zz_decode_RS2;
        end
      end
    end
  end

  assign execute_SRC_LESS_UNSIGNED = decode_to_execute_SRC_LESS_UNSIGNED;
  assign execute_SRC2_FORCE_ZERO = decode_to_execute_SRC2_FORCE_ZERO;
  assign execute_SRC2 = decode_to_execute_SRC2;
  assign execute_SRC_USE_SUB_LESS = decode_to_execute_SRC_USE_SUB_LESS;
  assign execute_SRC1 = decode_to_execute_SRC1;
  assign _zz_decode_to_execute_PC = decode_PC;
  assign _zz_decode_to_execute_RS2 = decode_RS2;
  assign decode_SRC2_CTRL = _zz_decode_SRC2_CTRL;
  assign _zz_decode_to_execute_RS1 = decode_RS1;
  assign decode_SRC1_CTRL = _zz_decode_SRC1_CTRL;
  assign decode_SRC_USE_SUB_LESS = _zz_decode_CfuPlugin_CFU_ENABLE[4];
  assign decode_SRC_ADD_ZERO = _zz_decode_CfuPlugin_CFU_ENABLE[19];
  assign _zz_lastStageRegFileWrite_payload_address = writeBack_INSTRUCTION;
  assign _zz_lastStageRegFileWrite_valid = writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    _zz_1 = 1'b0;
    if(lastStageRegFileWrite_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign decode_INSTRUCTION_ANTICIPATED = (decode_arbitration_isStuck ? decode_INSTRUCTION : IBusCachedPlugin_decompressor_output_payload_rsp_inst);
  always @(*) begin
    decode_REGFILE_WRITE_VALID = _zz_decode_CfuPlugin_CFU_ENABLE[11];
    if(when_RegFilePlugin_l63) begin
      decode_REGFILE_WRITE_VALID = 1'b0;
    end
  end

  always @(*) begin
    decode_LEGAL_INSTRUCTION = (|{((decode_INSTRUCTION & 32'h0000005f) == 32'h00000017),{((decode_INSTRUCTION & 32'h04000073) == 32'h00000043),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION) == 32'h0000006f),{(_zz_decode_LEGAL_INSTRUCTION_1 == _zz_decode_LEGAL_INSTRUCTION_2),{_zz_decode_LEGAL_INSTRUCTION_3,{_zz_decode_LEGAL_INSTRUCTION_4,_zz_decode_LEGAL_INSTRUCTION_5}}}}}});
    if(decode_FpuPlugin_trap) begin
      decode_LEGAL_INSTRUCTION = 1'b0;
    end
  end

  always @(*) begin
    _zz_decode_RS2_2 = writeBack_REGFILE_WRITE_DATA;
    if(when_DBusCachedPlugin_l599) begin
      _zz_decode_RS2_2 = writeBack_DBusCachedPlugin_rspFormated;
    end
    if(when_MulPlugin_l147) begin
      case(switch_MulPlugin_l148)
        2'b00 : begin
          _zz_decode_RS2_2 = _zz__zz_decode_RS2_2;
        end
        default : begin
          _zz_decode_RS2_2 = _zz__zz_decode_RS2_2_1;
        end
      endcase
    end
    if(writeBack_FpuPlugin_isRsp) begin
      if(writeBack_arbitration_isValid) begin
        _zz_decode_RS2_2 = FpuPlugin_port_rsp_payload_value[31 : 0];
      end
    end
    if(writeBack_CfuPlugin_CFU_IN_FLIGHT) begin
      _zz_decode_RS2_2 = writeBack_CfuPlugin_rsp_payload_outputs_0;
    end
  end

  assign writeBack_MEMORY_WR = memory_to_writeBack_MEMORY_WR;
  assign writeBack_MEMORY_FENCE = memory_to_writeBack_MEMORY_FENCE;
  assign writeBack_MEMORY_AMO = memory_to_writeBack_MEMORY_AMO;
  assign writeBack_MEMORY_LRSC = memory_to_writeBack_MEMORY_LRSC;
  assign writeBack_MEMORY_STORE_DATA_RF = memory_to_writeBack_MEMORY_STORE_DATA_RF;
  assign writeBack_REGFILE_WRITE_DATA = memory_to_writeBack_REGFILE_WRITE_DATA;
  assign writeBack_MEMORY_ENABLE = memory_to_writeBack_MEMORY_ENABLE;
  assign memory_PC = execute_to_memory_PC;
  assign memory_MEMORY_STORE_DATA_RF = execute_to_memory_MEMORY_STORE_DATA_RF;
  assign memory_REGFILE_WRITE_DATA = execute_to_memory_REGFILE_WRITE_DATA;
  assign memory_INSTRUCTION = execute_to_memory_INSTRUCTION;
  assign memory_MEMORY_WR = execute_to_memory_MEMORY_WR;
  assign memory_MEMORY_ENABLE = execute_to_memory_MEMORY_ENABLE;
  assign execute_MEMORY_FENCE_WR = decode_to_execute_MEMORY_FENCE_WR;
  assign memory_MEMORY_VIRTUAL_ADDRESS = execute_to_memory_MEMORY_VIRTUAL_ADDRESS;
  assign execute_MEMORY_AMO = decode_to_execute_MEMORY_AMO;
  assign execute_MEMORY_LRSC = decode_to_execute_MEMORY_LRSC;
  assign execute_MEMORY_FORCE_CONSTISTENCY = decode_to_execute_MEMORY_FORCE_CONSTISTENCY;
  assign execute_RS1 = decode_to_execute_RS1;
  assign execute_MEMORY_MANAGMENT = decode_to_execute_MEMORY_MANAGMENT;
  assign execute_RS2 = decode_to_execute_RS2;
  assign execute_MEMORY_WR = decode_to_execute_MEMORY_WR;
  assign execute_SRC_ADD = execute_SrcPlugin_addSub;
  assign execute_MEMORY_ENABLE = decode_to_execute_MEMORY_ENABLE;
  assign execute_INSTRUCTION = decode_to_execute_INSTRUCTION;
  assign decode_MEMORY_AMO = _zz_decode_CfuPlugin_CFU_ENABLE[17];
  assign decode_MEMORY_LRSC = _zz_decode_CfuPlugin_CFU_ENABLE[16];
  assign decode_MEMORY_ENABLE = _zz_decode_CfuPlugin_CFU_ENABLE[5];
  assign decode_FLUSH_ALL = _zz_decode_CfuPlugin_CFU_ENABLE[0];
  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_4 = IBusCachedPlugin_rsp_issueDetected_3;
    if(when_IBusCachedPlugin_l262) begin
      IBusCachedPlugin_rsp_issueDetected_4 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_3 = IBusCachedPlugin_rsp_issueDetected_2;
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_rsp_issueDetected_3 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_2 = IBusCachedPlugin_rsp_issueDetected_1;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_issueDetected_2 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_1 = IBusCachedPlugin_rsp_issueDetected;
    if(when_IBusCachedPlugin_l245) begin
      IBusCachedPlugin_rsp_issueDetected_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_memory_to_writeBack_FORMAL_PC_NEXT = memory_FORMAL_PC_NEXT;
    if(BranchPlugin_jumpInterface_valid) begin
      _zz_memory_to_writeBack_FORMAL_PC_NEXT = BranchPlugin_jumpInterface_payload;
    end
  end

  assign decode_PC = IBusCachedPlugin_decodePc_pcReg;
  assign decode_INSTRUCTION = IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  assign decode_IS_RVC = IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  assign writeBack_PC = memory_to_writeBack_PC;
  assign writeBack_INSTRUCTION = memory_to_writeBack_INSTRUCTION;
  always @(*) begin
    decode_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l356) begin
      decode_arbitration_haltItself = 1'b1;
    end
    if(when_FpuPlugin_l273) begin
      decode_arbitration_haltItself = 1'b1;
    end
    if(FpuPlugin_port_cmd_isStall) begin
      decode_arbitration_haltItself = 1'b1;
    end
    case(IBusCachedPlugin_injector_port_state)
      3'b010 : begin
        decode_arbitration_haltItself = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    decode_arbitration_haltByOther = 1'b0;
    if(when_HazardSimplePlugin_l113) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
        if(decode_arbitration_isValid) begin
          decode_arbitration_haltByOther = 1'b1;
        end
      end
      default : begin
      end
    endcase
    if(CsrPlugin_pipelineLiberator_active) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(when_CsrPlugin_l1671) begin
      decode_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    decode_arbitration_removeIt = 1'b0;
    if(_zz_when) begin
      decode_arbitration_removeIt = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      decode_arbitration_removeIt = 1'b1;
    end
  end

  assign decode_arbitration_flushIt = 1'b0;
  always @(*) begin
    decode_arbitration_flushNext = 1'b0;
    if(_zz_when) begin
      decode_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l398) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_DBusCachedPlugin_l427) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_CsrPlugin_l1735) begin
      if(execute_CsrPlugin_blockedBySideEffects) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
    if(when_MulPlugin_l65) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_CfuPlugin_l196) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_CfuPlugin_l203) begin
      execute_arbitration_haltItself = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_haltByOther = 1'b0;
    if(when_DBusCachedPlugin_l414) begin
      execute_arbitration_haltByOther = 1'b1;
    end
    if(when_FpuPlugin_l229) begin
      execute_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_removeIt = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_removeIt = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      execute_arbitration_removeIt = 1'b1;
    end
  end

  assign execute_arbitration_flushIt = 1'b0;
  always @(*) begin
    execute_arbitration_flushNext = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    memory_arbitration_haltItself = 1'b0;
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l129) begin
        memory_arbitration_haltItself = 1'b1;
      end
    end
  end

  always @(*) begin
    memory_arbitration_haltByOther = 1'b0;
    if(when_DBusCachedPlugin_l535) begin
      memory_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    memory_arbitration_removeIt = 1'b0;
    if(DBusCachedPlugin_trigger_hitBefore) begin
      memory_arbitration_removeIt = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      memory_arbitration_removeIt = 1'b1;
    end
  end

  assign memory_arbitration_flushIt = 1'b0;
  always @(*) begin
    memory_arbitration_flushNext = 1'b0;
    if(DBusCachedPlugin_trigger_hitBefore) begin
      memory_arbitration_flushNext = 1'b1;
    end
    if(BranchPlugin_jumpInterface_valid) begin
      memory_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l572) begin
      writeBack_arbitration_haltItself = 1'b1;
    end
    if(writeBack_CfuPlugin_CFU_IN_FLIGHT) begin
      if(when_CfuPlugin_l239) begin
        writeBack_arbitration_haltItself = 1'b1;
      end
    end
  end

  always @(*) begin
    writeBack_arbitration_haltByOther = 1'b0;
    if(writeBack_FpuPlugin_isRsp) begin
      if(when_FpuPlugin_l323) begin
        writeBack_arbitration_haltByOther = 1'b1;
      end
    end
    if(when_FpuPlugin_l339) begin
      writeBack_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_removeIt = 1'b0;
    if(DBusCachedPlugin_exceptionBus_valid) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
    if(writeBack_arbitration_isFlushed) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_flushIt = 1'b0;
    if(DBusCachedPlugin_redoBranch_valid) begin
      writeBack_arbitration_flushIt = 1'b1;
    end
    if(CsrPlugin_doResume) begin
      writeBack_arbitration_flushIt = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_flushNext = 1'b0;
    if(DBusCachedPlugin_redoBranch_valid) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(DBusCachedPlugin_exceptionBus_valid) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1534) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1600) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
  end

  assign lastStageInstruction = writeBack_INSTRUCTION;
  assign lastStagePc = writeBack_PC;
  assign lastStageIsValid = writeBack_arbitration_isValid;
  assign lastStageIsFiring = writeBack_arbitration_isFiring;
  always @(*) begin
    IBusCachedPlugin_fetcherHalt = 1'b0;
    if(when_CsrPlugin_l729) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1416) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1534) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1600) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
  end

  assign IBusCachedPlugin_forceNoDecodeCond = 1'b0;
  always @(*) begin
    IBusCachedPlugin_incomingInstruction = 1'b0;
    if(when_Fetcher_l242) begin
      IBusCachedPlugin_incomingInstruction = 1'b1;
    end
    if(IBusCachedPlugin_injector_decodeInput_valid) begin
      IBusCachedPlugin_incomingInstruction = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_csrMapping_allowCsrSignal = 1'b0;
    if(when_CsrPlugin_l1846) begin
      CsrPlugin_csrMapping_allowCsrSignal = 1'b1;
    end
    if(when_CsrPlugin_l1853) begin
      CsrPlugin_csrMapping_allowCsrSignal = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_csrMapping_doForceFailCsr = 1'b0;
    if(when_FpuPlugin_l253) begin
      CsrPlugin_csrMapping_doForceFailCsr = 1'b1;
    end
  end

  assign CsrPlugin_csrMapping_readDataSignal = CsrPlugin_csrMapping_readDataInit;
  assign CsrPlugin_inWfi = 1'b0;
  always @(*) begin
    CsrPlugin_thirdPartyWake = 1'b0;
    if(when_CsrPlugin_l880) begin
      CsrPlugin_thirdPartyWake = 1'b1;
    end
    if(decode_FpuPlugin_forked) begin
      CsrPlugin_thirdPartyWake = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_valid = 1'b0;
    if(when_CsrPlugin_l1534) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
    if(when_CsrPlugin_l1600) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
    if(CsrPlugin_doResume) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CsrPlugin_l1534) begin
      CsrPlugin_jumpInterface_payload = {CsrPlugin_xtvec_base,2'b00};
    end
    if(when_CsrPlugin_l1600) begin
      case(switch_CsrPlugin_l1604)
        2'b11 : begin
          CsrPlugin_jumpInterface_payload = CsrPlugin_mepc;
        end
        default : begin
        end
      endcase
    end
    if(CsrPlugin_doResume) begin
      CsrPlugin_jumpInterface_payload = CsrPlugin_dpc;
    end
  end

  assign CsrPlugin_forceMachineWire = 1'b0;
  always @(*) begin
    CsrPlugin_allowInterrupts = 1'b1;
    if(debugMode) begin
      CsrPlugin_allowInterrupts = 1'b0;
    end
  end

  assign CsrPlugin_allowException = 1'b1;
  assign CsrPlugin_allowEbreakException = 1'b1;
  always @(*) begin
    CsrPlugin_xretAwayFromMachine = 1'b0;
    if(when_CsrPlugin_l1600) begin
      case(switch_CsrPlugin_l1604)
        2'b11 : begin
          if(when_CsrPlugin_l1612) begin
            CsrPlugin_xretAwayFromMachine = 1'b1;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    BranchPlugin_inDebugNoFetchFlag = 1'b0;
    if(debugMode) begin
      BranchPlugin_inDebugNoFetchFlag = 1'b1;
    end
  end

  assign IBusCachedPlugin_mmuBus_rsp_physicalAddress = IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign IBusCachedPlugin_mmuBus_rsp_allowRead = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowWrite = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowExecute = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_isIoAccess = (((IBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'hf8000000) || ((IBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'he1000000));
  assign IBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign IBusCachedPlugin_mmuBus_busy = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_physicalAddress = DBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign DBusCachedPlugin_mmuBus_rsp_allowRead = 1'b1;
  assign DBusCachedPlugin_mmuBus_rsp_allowWrite = 1'b1;
  assign DBusCachedPlugin_mmuBus_rsp_allowExecute = 1'b1;
  assign DBusCachedPlugin_mmuBus_rsp_isIoAccess = (((DBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'hf8000000) || ((DBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'he1000000));
  assign DBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign DBusCachedPlugin_mmuBus_busy = 1'b0;
  assign IBusCachedPlugin_externalFlush = (|{writeBack_arbitration_flushNext,{memory_arbitration_flushNext,{execute_arbitration_flushNext,decode_arbitration_flushNext}}});
  assign IBusCachedPlugin_jump_pcLoad_valid = (|{BranchPlugin_jumpInterface_valid,{CsrPlugin_jumpInterface_valid,DBusCachedPlugin_redoBranch_valid}});
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload = {BranchPlugin_jumpInterface_valid,{CsrPlugin_jumpInterface_valid,DBusCachedPlugin_redoBranch_valid}};
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload & (~ _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1));
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_2 = _zz_IBusCachedPlugin_jump_pcLoad_payload_1[1];
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_3 = _zz_IBusCachedPlugin_jump_pcLoad_payload_1[2];
  assign IBusCachedPlugin_jump_pcLoad_payload = _zz_IBusCachedPlugin_jump_pcLoad_payload_4;
  always @(*) begin
    IBusCachedPlugin_fetchPc_correction = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
  end

  assign IBusCachedPlugin_fetchPc_output_fire = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign IBusCachedPlugin_fetchPc_corrected = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_correctionReg);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b0;
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b1;
    end
  end

  assign when_Fetcher_l133 = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_pcRegPropagate);
  assign when_Fetcher_l133_1 = ((! IBusCachedPlugin_fetchPc_output_valid) && IBusCachedPlugin_fetchPc_output_ready);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pc = (IBusCachedPlugin_fetchPc_pcReg + _zz_IBusCachedPlugin_fetchPc_pc);
    if(IBusCachedPlugin_fetchPc_inc) begin
      IBusCachedPlugin_fetchPc_pc[1] = 1'b0;
    end
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_fetchPc_redo_payload;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_jump_pcLoad_payload;
    end
    IBusCachedPlugin_fetchPc_pc[0] = 1'b0;
  end

  always @(*) begin
    IBusCachedPlugin_fetchPc_flushed = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
  end

  assign when_Fetcher_l160 = (IBusCachedPlugin_fetchPc_booted && ((IBusCachedPlugin_fetchPc_output_ready || IBusCachedPlugin_fetchPc_correction) || IBusCachedPlugin_fetchPc_pcRegPropagate));
  assign IBusCachedPlugin_fetchPc_output_valid = ((! IBusCachedPlugin_fetcherHalt) && IBusCachedPlugin_fetchPc_booted);
  assign IBusCachedPlugin_fetchPc_output_payload = IBusCachedPlugin_fetchPc_pc;
  always @(*) begin
    IBusCachedPlugin_decodePc_flushed = 1'b0;
    if(when_Fetcher_l194) begin
      IBusCachedPlugin_decodePc_flushed = 1'b1;
    end
  end

  assign IBusCachedPlugin_decodePc_pcPlus = (IBusCachedPlugin_decodePc_pcReg + _zz_IBusCachedPlugin_decodePc_pcPlus);
  always @(*) begin
    IBusCachedPlugin_decodePc_injectedDecode = 1'b0;
    if(when_Fetcher_l373) begin
      IBusCachedPlugin_decodePc_injectedDecode = 1'b1;
    end
  end

  assign when_Fetcher_l182 = (decode_arbitration_isFiring && (! IBusCachedPlugin_decodePc_injectedDecode));
  assign when_Fetcher_l194 = (IBusCachedPlugin_jump_pcLoad_valid && ((! decode_arbitration_isStuck) || decode_arbitration_removeIt));
  always @(*) begin
    IBusCachedPlugin_iBusRsp_redoFetch = 1'b0;
    if(IBusCachedPlugin_rsp_redoFetch) begin
      IBusCachedPlugin_iBusRsp_redoFetch = 1'b1;
    end
  end

  assign IBusCachedPlugin_iBusRsp_stages_0_input_valid = IBusCachedPlugin_fetchPc_output_valid;
  assign IBusCachedPlugin_fetchPc_output_ready = IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_0_input_payload = IBusCachedPlugin_fetchPc_output_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b0;
    if(IBusCachedPlugin_cache_io_cpu_prefetch_haltIt) begin
      IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready = (! IBusCachedPlugin_iBusRsp_stages_0_halt);
  assign IBusCachedPlugin_iBusRsp_stages_0_input_ready = (IBusCachedPlugin_iBusRsp_stages_0_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_valid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_payload = IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b0;
    if(IBusCachedPlugin_mmuBus_busy) begin
      IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready = (! IBusCachedPlugin_iBusRsp_stages_1_halt);
  assign IBusCachedPlugin_iBusRsp_stages_1_input_ready = (IBusCachedPlugin_iBusRsp_stages_1_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_valid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_payload = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b0;
    if(when_IBusCachedPlugin_l273) begin
      IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready = (! IBusCachedPlugin_iBusRsp_stages_2_halt);
  assign IBusCachedPlugin_iBusRsp_stages_2_input_ready = (IBusCachedPlugin_iBusRsp_stages_2_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_valid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_fetchPc_redo_valid = IBusCachedPlugin_iBusRsp_redoFetch;
  always @(*) begin
    IBusCachedPlugin_fetchPc_redo_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
    if(IBusCachedPlugin_decompressor_throw2BytesReg) begin
      IBusCachedPlugin_fetchPc_redo_payload[1] = 1'b1;
    end
  end

  assign IBusCachedPlugin_iBusRsp_flush = (IBusCachedPlugin_externalFlush || IBusCachedPlugin_iBusRsp_redoFetch);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_ready = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready = ((1'b0 && (! _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid)) || IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_payload = IBusCachedPlugin_fetchPc_pcReg;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_ready = ((1'b0 && (! IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid)) || IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_valid = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready = IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_payload = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_readyForError = 1'b1;
    if(IBusCachedPlugin_injector_decodeInput_valid) begin
      IBusCachedPlugin_iBusRsp_readyForError = 1'b0;
    end
  end

  assign when_Fetcher_l242 = (IBusCachedPlugin_iBusRsp_stages_1_input_valid || IBusCachedPlugin_iBusRsp_stages_2_input_valid);
  assign IBusCachedPlugin_decompressor_input_valid = (IBusCachedPlugin_iBusRsp_output_valid && (! IBusCachedPlugin_iBusRsp_redoFetch));
  assign IBusCachedPlugin_decompressor_input_payload_pc = IBusCachedPlugin_iBusRsp_output_payload_pc;
  assign IBusCachedPlugin_decompressor_input_payload_rsp_error = IBusCachedPlugin_iBusRsp_output_payload_rsp_error;
  assign IBusCachedPlugin_decompressor_input_payload_rsp_inst = IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  assign IBusCachedPlugin_decompressor_input_payload_isRvc = IBusCachedPlugin_iBusRsp_output_payload_isRvc;
  assign IBusCachedPlugin_iBusRsp_output_ready = IBusCachedPlugin_decompressor_input_ready;
  assign IBusCachedPlugin_decompressor_flushNext = 1'b0;
  assign IBusCachedPlugin_decompressor_consumeCurrent = 1'b0;
  assign IBusCachedPlugin_decompressor_isInputLowRvc = (IBusCachedPlugin_decompressor_input_payload_rsp_inst[1 : 0] != 2'b11);
  assign IBusCachedPlugin_decompressor_isInputHighRvc = (IBusCachedPlugin_decompressor_input_payload_rsp_inst[17 : 16] != 2'b11);
  assign IBusCachedPlugin_decompressor_throw2Bytes = (IBusCachedPlugin_decompressor_throw2BytesReg || IBusCachedPlugin_decompressor_input_payload_pc[1]);
  assign IBusCachedPlugin_decompressor_unaligned = (IBusCachedPlugin_decompressor_throw2Bytes || IBusCachedPlugin_decompressor_bufferValid);
  assign IBusCachedPlugin_decompressor_bufferValidPatched = (IBusCachedPlugin_decompressor_input_valid ? IBusCachedPlugin_decompressor_bufferValid : IBusCachedPlugin_decompressor_bufferValidLatch);
  assign IBusCachedPlugin_decompressor_throw2BytesPatched = (IBusCachedPlugin_decompressor_input_valid ? IBusCachedPlugin_decompressor_throw2Bytes : IBusCachedPlugin_decompressor_throw2BytesLatch);
  assign IBusCachedPlugin_decompressor_raw = (IBusCachedPlugin_decompressor_bufferValidPatched ? {IBusCachedPlugin_decompressor_input_payload_rsp_inst[15 : 0],IBusCachedPlugin_decompressor_bufferData} : {IBusCachedPlugin_decompressor_input_payload_rsp_inst[31 : 16],(IBusCachedPlugin_decompressor_throw2BytesPatched ? IBusCachedPlugin_decompressor_input_payload_rsp_inst[31 : 16] : IBusCachedPlugin_decompressor_input_payload_rsp_inst[15 : 0])});
  assign IBusCachedPlugin_decompressor_isRvc = (IBusCachedPlugin_decompressor_raw[1 : 0] != 2'b11);
  assign _zz_IBusCachedPlugin_decompressor_decompressed = IBusCachedPlugin_decompressor_raw[15 : 0];
  always @(*) begin
    IBusCachedPlugin_decompressor_decompressed = 32'h0;
    case(switch_Misc_l44)
      5'h0 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{{2'b00,_zz_IBusCachedPlugin_decompressor_decompressed[10 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 11]},_zz_IBusCachedPlugin_decompressor_decompressed[5]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},2'b00},5'h02},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h13};
        if(when_Misc_l47) begin
          IBusCachedPlugin_decompressor_decompressed = 32'h0;
        end
      end
      5'h01 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_4,_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h07};
      end
      5'h02 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_3,_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h03};
      end
      5'h03 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_3,_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h07};
      end
      5'h05 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_4[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed_2},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed_4[4 : 0]},7'h27};
      end
      5'h06 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_3[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed_2},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_3[4 : 0]},7'h23};
      end
      5'h07 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_3[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed_2},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_3[4 : 0]},7'h27};
      end
      5'h08 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_6,_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13};
      end
      5'h09 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_9[20],_zz_IBusCachedPlugin_decompressor_decompressed_9[10 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_9[11]},_zz_IBusCachedPlugin_decompressor_decompressed_9[19 : 12]},_zz_IBusCachedPlugin_decompressor_decompressed_21},7'h6f};
      end
      5'h0a : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_6,5'h0},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13};
      end
      5'h0b : begin
        IBusCachedPlugin_decompressor_decompressed = ((_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7] == 5'h02) ? {{{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_28,_zz_IBusCachedPlugin_decompressor_decompressed_29},_zz_IBusCachedPlugin_decompressor_decompressed_30},_zz_IBusCachedPlugin_decompressor_decompressed[6]},4'b0000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13} : {{_zz_IBusCachedPlugin_decompressor_decompressed_31[31 : 12],_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h37});
      end
      5'h0c : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{((_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] == 2'b10) ? _zz_IBusCachedPlugin_decompressor_decompressed_27 : {{1'b0,(_zz_IBusCachedPlugin_decompressor_decompressed_32 || _zz_IBusCachedPlugin_decompressor_decompressed_33)},5'h0}),(((! _zz_IBusCachedPlugin_decompressor_decompressed[11]) || _zz_IBusCachedPlugin_decompressor_decompressed_23) ? _zz_IBusCachedPlugin_decompressor_decompressed[6 : 2] : _zz_IBusCachedPlugin_decompressor_decompressed_2)},_zz_IBusCachedPlugin_decompressor_decompressed_1},_zz_IBusCachedPlugin_decompressor_decompressed_25},_zz_IBusCachedPlugin_decompressor_decompressed_1},(_zz_IBusCachedPlugin_decompressor_decompressed_23 ? 7'h13 : 7'h33)};
      end
      5'h0d : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_16[20],_zz_IBusCachedPlugin_decompressor_decompressed_16[10 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_16[11]},_zz_IBusCachedPlugin_decompressor_decompressed_16[19 : 12]},_zz_IBusCachedPlugin_decompressor_decompressed_20},7'h6f};
      end
      5'h0e : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_19[12],_zz_IBusCachedPlugin_decompressor_decompressed_19[10 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed_20},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed_19[4 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_19[11]},7'h63};
      end
      5'h0f : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_19[12],_zz_IBusCachedPlugin_decompressor_decompressed_19[10 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed_20},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b001},_zz_IBusCachedPlugin_decompressor_decompressed_19[4 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_19[11]},7'h63};
      end
      5'h10 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{7'h0,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b001},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13};
      end
      5'h11 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{3'b000,_zz_IBusCachedPlugin_decompressor_decompressed[4 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[12]},_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5]},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h07};
      end
      5'h12 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[3 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[12]},_zz_IBusCachedPlugin_decompressor_decompressed[6 : 4]},2'b00},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h03};
      end
      5'h13 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[3 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[12]},_zz_IBusCachedPlugin_decompressor_decompressed[6 : 4]},2'b00},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h07};
      end
      5'h14 : begin
        IBusCachedPlugin_decompressor_decompressed = ((_zz_IBusCachedPlugin_decompressor_decompressed[12 : 2] == 11'h400) ? 32'h00100073 : ((_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2] == 5'h0) ? {{{{12'h0,_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b000},(_zz_IBusCachedPlugin_decompressor_decompressed[12] ? _zz_IBusCachedPlugin_decompressor_decompressed_21 : _zz_IBusCachedPlugin_decompressor_decompressed_20)},7'h67} : {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_34,_zz_IBusCachedPlugin_decompressor_decompressed_35},(_zz_IBusCachedPlugin_decompressor_decompressed_36 ? _zz_IBusCachedPlugin_decompressor_decompressed_37 : _zz_IBusCachedPlugin_decompressor_decompressed_20)},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h33}));
      end
      5'h15 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_38[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed_39[4 : 0]},7'h27};
      end
      5'h16 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_40[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_41[4 : 0]},7'h23};
      end
      5'h17 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_42[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_43[4 : 0]},7'h27};
      end
      default : begin
      end
    endcase
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_1 = {2'b01,_zz_IBusCachedPlugin_decompressor_decompressed[9 : 7]};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_2 = {2'b01,_zz_IBusCachedPlugin_decompressor_decompressed[4 : 2]};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_3 = {{{{5'h0,_zz_IBusCachedPlugin_decompressor_decompressed[5]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_4 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},3'b000};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_5 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_6[11] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[10] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[9] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[8] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[7] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[6] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[5] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[4 : 0] = _zz_IBusCachedPlugin_decompressor_decompressed[6 : 2];
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_7 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_8[9] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[8] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[7] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[6] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[5] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[4] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[3] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[2] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[1] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[0] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_9 = {{{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_8,_zz_IBusCachedPlugin_decompressor_decompressed[8]},_zz_IBusCachedPlugin_decompressor_decompressed[10 : 9]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},_zz_IBusCachedPlugin_decompressor_decompressed[7]},_zz_IBusCachedPlugin_decompressor_decompressed[2]},_zz_IBusCachedPlugin_decompressor_decompressed[11]},_zz_IBusCachedPlugin_decompressor_decompressed[5 : 3]},1'b0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_10 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_11[14] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[13] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[12] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[11] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[10] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[9] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[8] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[7] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[6] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[5] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[4] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[3] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[2] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[1] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[0] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_12 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_13[2] = _zz_IBusCachedPlugin_decompressor_decompressed_12;
    _zz_IBusCachedPlugin_decompressor_decompressed_13[1] = _zz_IBusCachedPlugin_decompressor_decompressed_12;
    _zz_IBusCachedPlugin_decompressor_decompressed_13[0] = _zz_IBusCachedPlugin_decompressor_decompressed_12;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_14 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_15[9] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[8] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[7] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[6] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[5] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[4] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[3] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[2] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[1] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[0] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_16 = {{{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_15,_zz_IBusCachedPlugin_decompressor_decompressed[8]},_zz_IBusCachedPlugin_decompressor_decompressed[10 : 9]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},_zz_IBusCachedPlugin_decompressor_decompressed[7]},_zz_IBusCachedPlugin_decompressor_decompressed[2]},_zz_IBusCachedPlugin_decompressor_decompressed[11]},_zz_IBusCachedPlugin_decompressor_decompressed[5 : 3]},1'b0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_17 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_18[4] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[3] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[2] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[1] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[0] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_19 = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_18,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed[2]},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10]},_zz_IBusCachedPlugin_decompressor_decompressed[4 : 3]},1'b0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_20 = 5'h0;
  assign _zz_IBusCachedPlugin_decompressor_decompressed_21 = 5'h01;
  assign _zz_IBusCachedPlugin_decompressor_decompressed_22 = 5'h02;
  assign switch_Misc_l44 = {_zz_IBusCachedPlugin_decompressor_decompressed[1 : 0],_zz_IBusCachedPlugin_decompressor_decompressed[15 : 13]};
  assign when_Misc_l47 = (_zz_IBusCachedPlugin_decompressor_decompressed[12 : 2] == 11'h0);
  assign _zz_IBusCachedPlugin_decompressor_decompressed_23 = (_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] != 2'b11);
  assign switch_Misc_l241 = _zz_IBusCachedPlugin_decompressor_decompressed[11 : 10];
  assign switch_Misc_l241_1 = _zz_IBusCachedPlugin_decompressor_decompressed[6 : 5];
  always @(*) begin
    case(switch_Misc_l241_1)
      2'b00 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b000;
      end
      2'b01 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b100;
      end
      2'b10 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b110;
      end
      default : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b111;
      end
    endcase
  end

  always @(*) begin
    case(switch_Misc_l241)
      2'b00 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = 3'b101;
      end
      2'b01 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = 3'b101;
      end
      2'b10 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = 3'b111;
      end
      default : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = _zz_IBusCachedPlugin_decompressor_decompressed_24;
      end
    endcase
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_26 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_27[6] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[5] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[4] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[3] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[2] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[1] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[0] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
  end

  assign IBusCachedPlugin_decompressor_output_valid = (IBusCachedPlugin_decompressor_input_valid && (! ((IBusCachedPlugin_decompressor_throw2Bytes && (! IBusCachedPlugin_decompressor_bufferValid)) && (! IBusCachedPlugin_decompressor_isInputHighRvc))));
  assign IBusCachedPlugin_decompressor_output_payload_pc = IBusCachedPlugin_decompressor_input_payload_pc;
  assign IBusCachedPlugin_decompressor_output_payload_isRvc = IBusCachedPlugin_decompressor_isRvc;
  assign IBusCachedPlugin_decompressor_output_payload_rsp_inst = (IBusCachedPlugin_decompressor_isRvc ? IBusCachedPlugin_decompressor_decompressed : IBusCachedPlugin_decompressor_raw);
  assign IBusCachedPlugin_decompressor_input_ready = (IBusCachedPlugin_decompressor_output_ready && (((! IBusCachedPlugin_iBusRsp_stages_2_input_valid) || IBusCachedPlugin_decompressor_flushNext) || ((! (IBusCachedPlugin_decompressor_bufferValid && IBusCachedPlugin_decompressor_isInputHighRvc)) && (! (((! IBusCachedPlugin_decompressor_unaligned) && IBusCachedPlugin_decompressor_isInputLowRvc) && IBusCachedPlugin_decompressor_isInputHighRvc)))));
  assign IBusCachedPlugin_decompressor_output_fire = (IBusCachedPlugin_decompressor_output_valid && IBusCachedPlugin_decompressor_output_ready);
  assign IBusCachedPlugin_decompressor_bufferFill = (((((! IBusCachedPlugin_decompressor_unaligned) && IBusCachedPlugin_decompressor_isInputLowRvc) && (! IBusCachedPlugin_decompressor_isInputHighRvc)) || (IBusCachedPlugin_decompressor_bufferValid && (! IBusCachedPlugin_decompressor_isInputHighRvc))) || ((IBusCachedPlugin_decompressor_throw2Bytes && (! IBusCachedPlugin_decompressor_isRvc)) && (! IBusCachedPlugin_decompressor_isInputHighRvc)));
  assign when_Fetcher_l285 = (IBusCachedPlugin_decompressor_output_ready && IBusCachedPlugin_decompressor_input_valid);
  assign when_Fetcher_l288 = (IBusCachedPlugin_decompressor_output_ready && IBusCachedPlugin_decompressor_input_valid);
  assign when_Fetcher_l293 = (IBusCachedPlugin_externalFlush || IBusCachedPlugin_decompressor_consumeCurrent);
  assign IBusCachedPlugin_decompressor_output_ready = ((1'b0 && (! IBusCachedPlugin_injector_decodeInput_valid)) || IBusCachedPlugin_injector_decodeInput_ready);
  assign IBusCachedPlugin_injector_decodeInput_valid = _zz_IBusCachedPlugin_injector_decodeInput_valid;
  assign IBusCachedPlugin_injector_decodeInput_payload_pc = _zz_IBusCachedPlugin_injector_decodeInput_payload_pc;
  assign IBusCachedPlugin_injector_decodeInput_payload_rsp_error = _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_error;
  assign IBusCachedPlugin_injector_decodeInput_payload_rsp_inst = _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  assign IBusCachedPlugin_injector_decodeInput_payload_isRvc = _zz_IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  assign when_Fetcher_l331 = (! 1'b0);
  assign when_Fetcher_l331_1 = (! execute_arbitration_isStuck);
  assign when_Fetcher_l331_2 = (! memory_arbitration_isStuck);
  assign when_Fetcher_l331_3 = (! writeBack_arbitration_isStuck);
  assign IBusCachedPlugin_pcValids_0 = IBusCachedPlugin_injector_nextPcCalc_valids_0;
  assign IBusCachedPlugin_pcValids_1 = IBusCachedPlugin_injector_nextPcCalc_valids_1;
  assign IBusCachedPlugin_pcValids_2 = IBusCachedPlugin_injector_nextPcCalc_valids_2;
  assign IBusCachedPlugin_pcValids_3 = IBusCachedPlugin_injector_nextPcCalc_valids_3;
  assign IBusCachedPlugin_injector_decodeInput_ready = (! decode_arbitration_isStuck);
  always @(*) begin
    decode_arbitration_isValid = IBusCachedPlugin_injector_decodeInput_valid;
    case(IBusCachedPlugin_injector_port_state)
      3'b010 : begin
        decode_arbitration_isValid = 1'b1;
      end
      3'b011 : begin
        decode_arbitration_isValid = 1'b1;
      end
      default : begin
      end
    endcase
    if(IBusCachedPlugin_forceNoDecodeCond) begin
      decode_arbitration_isValid = 1'b0;
    end
  end

  assign iBus_cmd_valid = IBusCachedPlugin_cache_io_mem_cmd_valid;
  always @(*) begin
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  end

  assign iBus_cmd_payload_size = IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  assign IBusCachedPlugin_s0_tightlyCoupledHit = 1'b0;
  assign IBusCachedPlugin_cache_io_cpu_prefetch_isValid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && (! IBusCachedPlugin_s0_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isValid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && (! IBusCachedPlugin_s1_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_isValid = IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  assign IBusCachedPlugin_mmuBus_cmd_0_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_virtualAddress = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  assign IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign IBusCachedPlugin_mmuBus_end = (IBusCachedPlugin_iBusRsp_stages_1_input_ready || IBusCachedPlugin_externalFlush);
  assign IBusCachedPlugin_cache_io_cpu_decode_isValid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && (! IBusCachedPlugin_s2_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_decode_isStuck = (! IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_cache_io_cpu_decode_isUser = (CsrPlugin_privilege == 2'b00);
  assign IBusCachedPlugin_rsp_iBusRspOutputHalt = 1'b0;
  assign IBusCachedPlugin_rsp_issueDetected = 1'b0;
  always @(*) begin
    IBusCachedPlugin_rsp_redoFetch = 1'b0;
    if(when_IBusCachedPlugin_l245) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_cache_io_cpu_fill_valid = (IBusCachedPlugin_rsp_redoFetch && (! IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling));
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_cache_io_cpu_fill_valid = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_valid = 1'b0;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
    if(when_IBusCachedPlugin_l262) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_payload_code = 4'bxxxx;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b1100;
    end
    if(when_IBusCachedPlugin_l262) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b0001;
    end
  end

  assign IBusCachedPlugin_decodeExceptionPort_payload_badAddr = {IBusCachedPlugin_iBusRsp_stages_2_input_payload[31 : 2],2'b00};
  assign when_IBusCachedPlugin_l245 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling) && (! IBusCachedPlugin_rsp_issueDetected));
  assign when_IBusCachedPlugin_l250 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuException) && (! IBusCachedPlugin_rsp_issueDetected_1));
  assign when_IBusCachedPlugin_l256 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_cacheMiss) && (! IBusCachedPlugin_rsp_issueDetected_2));
  assign when_IBusCachedPlugin_l262 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_error) && (! IBusCachedPlugin_rsp_issueDetected_3));
  assign when_IBusCachedPlugin_l273 = (IBusCachedPlugin_rsp_issueDetected_4 || IBusCachedPlugin_rsp_iBusRspOutputHalt);
  assign IBusCachedPlugin_iBusRsp_output_valid = IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  assign IBusCachedPlugin_iBusRsp_stages_2_output_ready = IBusCachedPlugin_iBusRsp_output_ready;
  assign IBusCachedPlugin_iBusRsp_output_payload_rsp_inst = IBusCachedPlugin_cache_io_cpu_decode_data;
  assign IBusCachedPlugin_iBusRsp_output_payload_pc = IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  assign IBusCachedPlugin_cache_io_flush = (decode_arbitration_isValid && decode_FLUSH_ALL);
  assign dataCache_2_io_mem_cmd_s2mPipe_valid = (dataCache_2_io_mem_cmd_valid || (! dataCache_2_io_mem_cmd_rValidN));
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_wr = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_wr : dataCache_2_io_mem_cmd_rData_wr);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_uncached = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_uncached : dataCache_2_io_mem_cmd_rData_uncached);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_address = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_address : dataCache_2_io_mem_cmd_rData_address);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_data = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_data : dataCache_2_io_mem_cmd_rData_data);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_mask = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_mask : dataCache_2_io_mem_cmd_rData_mask);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_size = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_size : dataCache_2_io_mem_cmd_rData_size);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_exclusive = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_exclusive : dataCache_2_io_mem_cmd_rData_exclusive);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_last = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_last : dataCache_2_io_mem_cmd_rData_last);
  always @(*) begin
    dataCache_2_io_mem_cmd_s2mPipe_ready = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375) begin
      dataCache_2_io_mem_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid);
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid = dataCache_2_io_mem_cmd_s2mPipe_rValid;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_wr = dataCache_2_io_mem_cmd_s2mPipe_rData_wr;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached = dataCache_2_io_mem_cmd_s2mPipe_rData_uncached;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_address = dataCache_2_io_mem_cmd_s2mPipe_rData_address;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_data = dataCache_2_io_mem_cmd_s2mPipe_rData_data;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_mask = dataCache_2_io_mem_cmd_s2mPipe_rData_mask;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_size = dataCache_2_io_mem_cmd_s2mPipe_rData_size;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_exclusive = dataCache_2_io_mem_cmd_s2mPipe_rData_exclusive;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_last = dataCache_2_io_mem_cmd_s2mPipe_rData_last;
  assign dBus_cmd_valid = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_ready = dBus_cmd_ready;
  assign dBus_cmd_payload_wr = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_wr;
  assign dBus_cmd_payload_uncached = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached;
  assign dBus_cmd_payload_address = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_address;
  assign dBus_cmd_payload_data = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_data;
  assign dBus_cmd_payload_mask = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_mask;
  assign dBus_cmd_payload_size = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_size;
  assign dBus_cmd_payload_exclusive = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_exclusive;
  assign dBus_cmd_payload_last = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_last;
  assign when_DBusCachedPlugin_l334 = (dBus_rsp_valid && (! dataCache_2_io_cpu_writeBack_keepMemRspData));
  assign dBus_inv_ready = dataCache_2_io_mem_inv_ready;
  assign dBus_ack_valid = dataCache_2_io_mem_ack_valid;
  assign dBus_ack_payload_last = dataCache_2_io_mem_ack_payload_last;
  assign dBus_ack_payload_fragment_hit = dataCache_2_io_mem_ack_payload_fragment_hit;
  assign dBus_sync_ready = dataCache_2_io_mem_sync_ready;
  assign when_DBusCachedPlugin_l356 = ((DBusCachedPlugin_mmuBus_busy && decode_arbitration_isValid) && decode_MEMORY_ENABLE);
  always @(*) begin
    _zz_decode_MEMORY_FORCE_CONSTISTENCY = 1'b0;
    if(when_DBusCachedPlugin_l364) begin
      if(decode_MEMORY_LRSC) begin
        _zz_decode_MEMORY_FORCE_CONSTISTENCY = 1'b1;
      end
      if(decode_MEMORY_AMO) begin
        _zz_decode_MEMORY_FORCE_CONSTISTENCY = 1'b1;
      end
    end
  end

  assign when_DBusCachedPlugin_l364 = decode_INSTRUCTION[25];
  assign execute_DBusCachedPlugin_size = execute_INSTRUCTION[13 : 12];
  assign dataCache_2_io_cpu_execute_isValid = (execute_arbitration_isValid && execute_MEMORY_ENABLE);
  assign dataCache_2_io_cpu_execute_address = execute_SRC_ADD;
  always @(*) begin
    case(execute_DBusCachedPlugin_size)
      2'b00 : begin
        _zz_execute_MEMORY_STORE_DATA_RF = {{{execute_RS2[7 : 0],execute_RS2[7 : 0]},execute_RS2[7 : 0]},execute_RS2[7 : 0]};
      end
      2'b01 : begin
        _zz_execute_MEMORY_STORE_DATA_RF = {execute_RS2[15 : 0],execute_RS2[15 : 0]};
      end
      default : begin
        _zz_execute_MEMORY_STORE_DATA_RF = execute_RS2[31 : 0];
      end
    endcase
  end

  assign dataCache_2_io_cpu_flush_valid = (execute_arbitration_isValid && execute_MEMORY_MANAGMENT);
  assign dataCache_2_io_cpu_flush_payload_singleLine = (execute_INSTRUCTION[19 : 15] != 5'h0);
  assign dataCache_2_io_cpu_flush_payload_lineId = _zz_io_cpu_flush_payload_lineId[5:0];
  assign dataCache_2_io_cpu_flush_isStall = (dataCache_2_io_cpu_flush_valid && (! dataCache_2_io_cpu_flush_ready));
  assign when_DBusCachedPlugin_l398 = (dataCache_2_io_cpu_flush_isStall || dataCache_2_io_cpu_execute_haltIt);
  always @(*) begin
    dataCache_2_io_cpu_execute_args_isLrsc = 1'b0;
    if(execute_MEMORY_LRSC) begin
      dataCache_2_io_cpu_execute_args_isLrsc = 1'b1;
    end
  end

  assign dataCache_2_io_cpu_execute_args_amoCtrl_alu = execute_INSTRUCTION[31 : 29];
  assign dataCache_2_io_cpu_execute_args_amoCtrl_swap = execute_INSTRUCTION[27];
  assign when_DBusCachedPlugin_l414 = (dataCache_2_io_cpu_execute_refilling && execute_arbitration_isValid);
  assign when_DBusCachedPlugin_l427 = ((execute_arbitration_isValid && execute_MEMORY_FENCE_WR) && dataCache_2_io_cpu_writesPending);
  assign DBusCachedPlugin_writesPending = dataCache_2_io_cpu_writesPending;
  assign dataCache_2_io_cpu_memory_isValid = (memory_arbitration_isValid && memory_MEMORY_ENABLE);
  assign DBusCachedPlugin_mmuBus_cmd_0_isValid = dataCache_2_io_cpu_memory_isValid;
  assign DBusCachedPlugin_mmuBus_cmd_0_isStuck = memory_arbitration_isStuck;
  assign DBusCachedPlugin_mmuBus_cmd_0_virtualAddress = memory_MEMORY_VIRTUAL_ADDRESS;
  assign DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign DBusCachedPlugin_mmuBus_end = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  always @(*) begin
    dataCache_2_io_cpu_memory_mmuRsp_isIoAccess = DBusCachedPlugin_mmuBus_rsp_isIoAccess;
    if(when_DBusCachedPlugin_l476) begin
      dataCache_2_io_cpu_memory_mmuRsp_isIoAccess = 1'b1;
    end
  end

  assign when_DBusCachedPlugin_l476 = (1'b0 && (! dataCache_2_io_cpu_memory_isWrite));
  assign DBusCachedPlugin_trigger_valid = (((memory_arbitration_isValid && (! memory_arbitration_isStuck)) && (! memory_arbitration_isFlushed)) && memory_MEMORY_ENABLE);
  assign DBusCachedPlugin_trigger_load = (! memory_MEMORY_WR);
  assign DBusCachedPlugin_trigger_store = memory_MEMORY_WR;
  assign DBusCachedPlugin_trigger_size = memory_INSTRUCTION[13 : 12];
  assign DBusCachedPlugin_trigger_virtual = memory_REGFILE_WRITE_DATA;
  assign DBusCachedPlugin_trigger_writeData = memory_MEMORY_STORE_DATA_RF;
  assign DBusCachedPlugin_trigger_readData = 32'h0;
  assign DBusCachedPlugin_trigger_readDataValid = 1'b0;
  assign DBusCachedPlugin_trigger_dpc = memory_PC;
  always @(*) begin
    dataCache_2_io_cpu_writeBack_isValid = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
    if(writeBack_arbitration_haltByOther) begin
      dataCache_2_io_cpu_writeBack_isValid = 1'b0;
    end
  end

  assign dataCache_2_io_cpu_writeBack_isUser = (CsrPlugin_privilege == 2'b00);
  assign dataCache_2_io_cpu_writeBack_address = writeBack_REGFILE_WRITE_DATA;
  always @(*) begin
    dataCache_2_io_cpu_writeBack_storeData[31 : 0] = writeBack_MEMORY_STORE_DATA_RF;
    dataCache_2_io_cpu_writeBack_storeData[63 : 32] = writeBack_MEMORY_STORE_DATA_RF;
    if(DBusBypass0_cond) begin
      dataCache_2_io_cpu_writeBack_storeData[63 : 0] = DBusBypass0_value;
    end
  end

  assign _zz_io_cpu_writeBack_fence_SW = writeBack_INSTRUCTION[31 : 20];
  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SW = _zz_io_cpu_writeBack_fence_SW[0];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SW = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SW = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SR = _zz_io_cpu_writeBack_fence_SW[1];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SR = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SR = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SO = _zz_io_cpu_writeBack_fence_SW[2];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SO = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SO = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SI = _zz_io_cpu_writeBack_fence_SW[3];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SI = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SI = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PW = _zz_io_cpu_writeBack_fence_SW[4];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PW = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PW = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PR = _zz_io_cpu_writeBack_fence_SW[5];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PR = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PR = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PO = _zz_io_cpu_writeBack_fence_SW[6];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PO = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PO = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PI = _zz_io_cpu_writeBack_fence_SW[7];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PI = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PI = 1'b0;
    end
  end

  assign dataCache_2_io_cpu_writeBack_fence_FM = _zz_io_cpu_writeBack_fence_SW[11 : 8];
  always @(*) begin
    writeBack_DBusCachedPlugin_fence_aquire = 1'b0;
    if(when_DBusCachedPlugin_l518) begin
      if(writeBack_MEMORY_LRSC) begin
        writeBack_DBusCachedPlugin_fence_aquire = 1'b1;
      end
      if(writeBack_MEMORY_AMO) begin
        writeBack_DBusCachedPlugin_fence_aquire = 1'b1;
      end
    end
  end

  assign when_DBusCachedPlugin_l518 = (writeBack_MEMORY_ENABLE && writeBack_INSTRUCTION[26]);
  assign when_DBusCachedPlugin_l531 = ((! writeBack_MEMORY_FENCE) || (! writeBack_arbitration_isFiring));
  assign when_DBusCachedPlugin_l535 = (writeBack_arbitration_isValid && (writeBack_MEMORY_FENCE || writeBack_DBusCachedPlugin_fence_aquire));
  always @(*) begin
    DBusCachedPlugin_redoBranch_valid = 1'b0;
    if(when_DBusCachedPlugin_l552) begin
      if(dataCache_2_io_cpu_redo) begin
        DBusCachedPlugin_redoBranch_valid = 1'b1;
      end
    end
  end

  assign DBusCachedPlugin_redoBranch_payload = writeBack_PC;
  always @(*) begin
    DBusCachedPlugin_exceptionBus_valid = 1'b0;
    if(when_DBusCachedPlugin_l552) begin
      if(dataCache_2_io_cpu_writeBack_accessError) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_2_io_cpu_writeBack_mmuException) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_2_io_cpu_writeBack_unalignedAccess) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_2_io_cpu_redo) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b0;
      end
    end
  end

  assign DBusCachedPlugin_exceptionBus_payload_badAddr = writeBack_REGFILE_WRITE_DATA;
  always @(*) begin
    DBusCachedPlugin_exceptionBus_payload_code = 4'bxxxx;
    if(when_DBusCachedPlugin_l552) begin
      if(dataCache_2_io_cpu_writeBack_accessError) begin
        DBusCachedPlugin_exceptionBus_payload_code = {1'd0, _zz_DBusCachedPlugin_exceptionBus_payload_code};
      end
      if(dataCache_2_io_cpu_writeBack_mmuException) begin
        DBusCachedPlugin_exceptionBus_payload_code = (writeBack_MEMORY_WR ? 4'b1111 : 4'b1101);
      end
      if(dataCache_2_io_cpu_writeBack_unalignedAccess) begin
        DBusCachedPlugin_exceptionBus_payload_code = {1'd0, _zz_DBusCachedPlugin_exceptionBus_payload_code_1};
      end
    end
  end

  assign when_DBusCachedPlugin_l552 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign when_DBusCachedPlugin_l572 = (dataCache_2_io_cpu_writeBack_isValid && dataCache_2_io_cpu_writeBack_haltIt);
  assign writeBack_DBusCachedPlugin_rspData = dataCache_2_io_cpu_writeBack_data;
  assign writeBack_DBusCachedPlugin_rspSplits_0 = writeBack_DBusCachedPlugin_rspData[7 : 0];
  assign writeBack_DBusCachedPlugin_rspSplits_1 = writeBack_DBusCachedPlugin_rspData[15 : 8];
  assign writeBack_DBusCachedPlugin_rspSplits_2 = writeBack_DBusCachedPlugin_rspData[23 : 16];
  assign writeBack_DBusCachedPlugin_rspSplits_3 = writeBack_DBusCachedPlugin_rspData[31 : 24];
  assign writeBack_DBusCachedPlugin_rspSplits_4 = writeBack_DBusCachedPlugin_rspData[39 : 32];
  assign writeBack_DBusCachedPlugin_rspSplits_5 = writeBack_DBusCachedPlugin_rspData[47 : 40];
  assign writeBack_DBusCachedPlugin_rspSplits_6 = writeBack_DBusCachedPlugin_rspData[55 : 48];
  assign writeBack_DBusCachedPlugin_rspSplits_7 = writeBack_DBusCachedPlugin_rspData[63 : 56];
  always @(*) begin
    writeBack_DBusCachedPlugin_rspShifted[7 : 0] = _zz_writeBack_DBusCachedPlugin_rspShifted;
    writeBack_DBusCachedPlugin_rspShifted[15 : 8] = _zz_writeBack_DBusCachedPlugin_rspShifted_2;
    writeBack_DBusCachedPlugin_rspShifted[23 : 16] = _zz_writeBack_DBusCachedPlugin_rspShifted_4;
    writeBack_DBusCachedPlugin_rspShifted[31 : 24] = _zz_writeBack_DBusCachedPlugin_rspShifted_6;
    writeBack_DBusCachedPlugin_rspShifted[39 : 32] = writeBack_DBusCachedPlugin_rspSplits_4;
    writeBack_DBusCachedPlugin_rspShifted[47 : 40] = writeBack_DBusCachedPlugin_rspSplits_5;
    writeBack_DBusCachedPlugin_rspShifted[55 : 48] = writeBack_DBusCachedPlugin_rspSplits_6;
    writeBack_DBusCachedPlugin_rspShifted[63 : 56] = writeBack_DBusCachedPlugin_rspSplits_7;
  end

  always @(*) begin
    writeBack_DBusCachedPlugin_rspRf = writeBack_DBusCachedPlugin_rspShifted[31 : 0];
    if(when_DBusCachedPlugin_l589) begin
      writeBack_DBusCachedPlugin_rspRf = {31'd0, _zz_writeBack_DBusCachedPlugin_rspRf};
    end
  end

  assign when_DBusCachedPlugin_l589 = (writeBack_MEMORY_LRSC && writeBack_MEMORY_WR);
  assign switch_Misc_l241_2 = writeBack_INSTRUCTION[13 : 12];
  assign _zz_writeBack_DBusCachedPlugin_rspFormated = (writeBack_DBusCachedPlugin_rspRf[7] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[31] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[30] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[29] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[28] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[27] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[26] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[25] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[24] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[23] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[22] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[21] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[20] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[19] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[18] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[17] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[16] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[15] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[14] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[13] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[12] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[11] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[10] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[9] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[8] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[7 : 0] = writeBack_DBusCachedPlugin_rspRf[7 : 0];
  end

  assign _zz_writeBack_DBusCachedPlugin_rspFormated_2 = (writeBack_DBusCachedPlugin_rspRf[15] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[31] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[30] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[29] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[28] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[27] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[26] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[25] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[24] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[23] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[22] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[21] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[20] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[19] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[18] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[17] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[16] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[15 : 0] = writeBack_DBusCachedPlugin_rspRf[15 : 0];
  end

  always @(*) begin
    case(switch_Misc_l241_2)
      2'b00 : begin
        writeBack_DBusCachedPlugin_rspFormated = _zz_writeBack_DBusCachedPlugin_rspFormated_1;
      end
      2'b01 : begin
        writeBack_DBusCachedPlugin_rspFormated = _zz_writeBack_DBusCachedPlugin_rspFormated_3;
      end
      default : begin
        writeBack_DBusCachedPlugin_rspFormated = writeBack_DBusCachedPlugin_rspRf;
      end
    endcase
  end

  assign when_DBusCachedPlugin_l599 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_1 = ((decode_INSTRUCTION & 32'h00007054) == 32'h00001004);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_2 = ((decode_INSTRUCTION & 32'h00004050) == 32'h00004050);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_3 = ((decode_INSTRUCTION & 32'h00000014) == 32'h00000014);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_4 = ((decode_INSTRUCTION & 32'h00000058) == 32'h0);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_5 = ((decode_INSTRUCTION & 32'h00000070) == 32'h00000020);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_6 = ((decode_INSTRUCTION & 32'h00002004) == 32'h00000004);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_7 = ((decode_INSTRUCTION & 32'h00000008) == 32'h00000008);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_8 = ((decode_INSTRUCTION & 32'h90000010) == 32'h80000010);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_9 = ((decode_INSTRUCTION & 32'h0000000c) == 32'h00000004);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_10 = ((decode_INSTRUCTION & 32'h0000004c) == 32'h00000008);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_11 = ((decode_INSTRUCTION & 32'h00001000) == 32'h0);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_12 = ((decode_INSTRUCTION & 32'h00000020) == 32'h00000020);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_13 = ((decode_INSTRUCTION & 32'hc0000010) == 32'h40000010);
  assign _zz_decode_CfuPlugin_CFU_ENABLE = {(|((decode_INSTRUCTION & 32'h02007054) == 32'h00005010)),{(|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE == _zz__zz_decode_CfuPlugin_CFU_ENABLE_1),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_2 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_3)}),{(|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_4 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_5)),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_6),{1'b0,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_7,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_8,_zz__zz_decode_CfuPlugin_CFU_ENABLE_13}}}}}}};
  assign _zz_decode_SRC1_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[3 : 2];
  assign _zz_decode_SRC1_CTRL_1 = _zz_decode_SRC1_CTRL_2;
  assign _zz_decode_ALU_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[8 : 7];
  assign _zz_decode_ALU_CTRL_1 = _zz_decode_ALU_CTRL_2;
  assign _zz_decode_SRC2_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[10 : 9];
  assign _zz_decode_SRC2_CTRL_1 = _zz_decode_SRC2_CTRL_2;
  assign _zz_decode_ENV_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[24 : 23];
  assign _zz_decode_ENV_CTRL_1 = _zz_decode_ENV_CTRL_2;
  assign _zz_decode_BRANCH_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[26 : 25];
  assign _zz_decode_BRANCH_CTRL_1 = _zz_decode_BRANCH_CTRL_2;
  assign _zz_decode_FPU_ENABLE = _zz_decode_CfuPlugin_CFU_ENABLE[32];
  assign _zz_decode_FPU_OPCODE_2 = _zz_decode_CfuPlugin_CFU_ENABLE[38 : 35];
  assign _zz_decode_FPU_OPCODE_1 = _zz_decode_FPU_OPCODE_2;
  assign _zz_decode_FPU_FORMAT_2 = _zz_decode_CfuPlugin_CFU_ENABLE[39 : 39];
  assign _zz_decode_FPU_FORMAT_1 = _zz_decode_FPU_FORMAT_2;
  assign _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2 = _zz_decode_CfuPlugin_CFU_ENABLE[43 : 43];
  assign _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1 = _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2;
  assign _zz_decode_ALU_BITWISE_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[45 : 44];
  assign _zz_decode_ALU_BITWISE_CTRL_1 = _zz_decode_ALU_BITWISE_CTRL_2;
  assign _zz_decode_SHIFT_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[47 : 46];
  assign _zz_decode_SHIFT_CTRL_1 = _zz_decode_SHIFT_CTRL_2;
  assign decodeExceptionPort_valid = (decode_arbitration_isValid && (! decode_LEGAL_INSTRUCTION));
  assign decodeExceptionPort_payload_code = 4'b0010;
  assign decodeExceptionPort_payload_badAddr = decode_INSTRUCTION;
  assign when_RegFilePlugin_l63 = (decode_INSTRUCTION[11 : 7] == 5'h0);
  assign decode_RegFilePlugin_regFileReadAddress1 = decode_INSTRUCTION_ANTICIPATED[19 : 15];
  assign decode_RegFilePlugin_regFileReadAddress2 = decode_INSTRUCTION_ANTICIPATED[24 : 20];
  assign decode_RegFilePlugin_rs1Data = RegFilePlugin_regFile_spinal_port0;
  assign decode_RegFilePlugin_rs2Data = RegFilePlugin_regFile_spinal_port1;
  always @(*) begin
    lastStageRegFileWrite_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
    if(_zz_5) begin
      lastStageRegFileWrite_valid = 1'b1;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
    if(_zz_5) begin
      lastStageRegFileWrite_payload_address = 5'h0;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_data = _zz_decode_RS2_2;
    if(_zz_5) begin
      lastStageRegFileWrite_payload_data = 32'h0;
    end
  end

  always @(*) begin
    case(decode_SRC1_CTRL)
      Src1CtrlEnum_RS : begin
        _zz_decode_SRC1 = _zz_decode_to_execute_RS1;
      end
      Src1CtrlEnum_PC_INCREMENT : begin
        _zz_decode_SRC1 = {29'd0, _zz__zz_decode_SRC1};
      end
      Src1CtrlEnum_IMU : begin
        _zz_decode_SRC1 = {decode_INSTRUCTION[31 : 12],12'h0};
      end
      default : begin
        _zz_decode_SRC1 = {27'd0, _zz__zz_decode_SRC1_1};
      end
    endcase
  end

  assign _zz_decode_SRC2 = decode_INSTRUCTION[31];
  always @(*) begin
    _zz_decode_SRC2_1[19] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[18] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[17] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[16] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[15] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[14] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[13] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[12] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[11] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[10] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[9] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[8] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[7] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[6] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[5] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[4] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[3] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[2] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[1] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[0] = _zz_decode_SRC2;
  end

  assign _zz_decode_SRC2_2 = _zz__zz_decode_SRC2_2[11];
  always @(*) begin
    _zz_decode_SRC2_3[19] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[18] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[17] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[16] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[15] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[14] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[13] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[12] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[11] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[10] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[9] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[8] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[7] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[6] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[5] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[4] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[3] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[2] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[1] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[0] = _zz_decode_SRC2_2;
  end

  always @(*) begin
    case(decode_SRC2_CTRL)
      Src2CtrlEnum_RS : begin
        _zz_decode_SRC2_4 = _zz_decode_to_execute_RS2;
      end
      Src2CtrlEnum_IMI : begin
        _zz_decode_SRC2_4 = {_zz_decode_SRC2_1,decode_INSTRUCTION[31 : 20]};
      end
      Src2CtrlEnum_IMS : begin
        _zz_decode_SRC2_4 = {_zz_decode_SRC2_3,{decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]}};
      end
      default : begin
        _zz_decode_SRC2_4 = _zz_decode_to_execute_PC;
      end
    endcase
  end

  always @(*) begin
    execute_SrcPlugin_addSub = _zz_execute_SrcPlugin_addSub;
    if(execute_SRC2_FORCE_ZERO) begin
      execute_SrcPlugin_addSub = execute_SRC1;
    end
  end

  assign execute_SrcPlugin_less = ((execute_SRC1[31] == execute_SRC2[31]) ? execute_SrcPlugin_addSub[31] : (execute_SRC_LESS_UNSIGNED ? execute_SRC2[31] : execute_SRC1[31]));
  always @(*) begin
    HazardSimplePlugin_src0Hazard = 1'b0;
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l48) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l48_1) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l48_2) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l105) begin
      HazardSimplePlugin_src0Hazard = 1'b0;
    end
  end

  always @(*) begin
    HazardSimplePlugin_src1Hazard = 1'b0;
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l51) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l51_1) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l51_2) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l108) begin
      HazardSimplePlugin_src1Hazard = 1'b0;
    end
  end

  assign HazardSimplePlugin_writeBackWrites_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
  assign HazardSimplePlugin_writeBackWrites_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
  assign HazardSimplePlugin_writeBackWrites_payload_data = _zz_decode_RS2_2;
  assign HazardSimplePlugin_addr0Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[19 : 15]);
  assign HazardSimplePlugin_addr1Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l47 = 1'b1;
  assign when_HazardSimplePlugin_l48 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58 = (1'b0 || (! when_HazardSimplePlugin_l47));
  assign when_HazardSimplePlugin_l48_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_1 = (1'b0 || (! memory_BYPASSABLE_MEMORY_STAGE));
  assign when_HazardSimplePlugin_l48_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_2 = (1'b0 || (! execute_BYPASSABLE_EXECUTE_STAGE));
  assign when_HazardSimplePlugin_l105 = (! decode_RS1_USE);
  assign when_HazardSimplePlugin_l108 = (! decode_RS2_USE);
  assign when_HazardSimplePlugin_l113 = (decode_arbitration_isValid && (HazardSimplePlugin_src0Hazard || HazardSimplePlugin_src1Hazard));
  always @(*) begin
    when_CsrPlugin_l836 = 1'b0;
    if(when_CsrPlugin_l1534) begin
      when_CsrPlugin_l836 = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_privilege = _zz_CsrPlugin_privilege;
    if(CsrPlugin_forceMachineWire) begin
      CsrPlugin_privilege = 2'b11;
    end
  end

  assign debugMode = (! CsrPlugin_running);
  assign when_CsrPlugin_l729 = (! CsrPlugin_running);
  always @(*) begin
    debugBus_resume_rsp_valid = 1'b0;
    if(CsrPlugin_doResume) begin
      debugBus_resume_rsp_valid = 1'b1;
    end
  end

  assign debugBus_running = CsrPlugin_running;
  assign debugBus_halted = (! CsrPlugin_running);
  assign debugBus_unavailable = systemCd_logic_outputReset_buffercc_io_dataOut;
  assign debugBus_haveReset = _zz_debugBus_haveReset;
  assign CsrPlugin_enterHalt = ((! CsrPlugin_running_aheadValue) && CsrPlugin_running_aheadValue_regNext);
  assign when_CsrPlugin_l747 = ((debugBus_haltReq && debugBus_running) && (! debugMode));
  assign CsrPlugin_forceResume = 1'b0;
  assign CsrPlugin_doResume = (CsrPlugin_forceResume || _zz_CsrPlugin_doResume);
  always @(*) begin
    CsrPlugin_timeout_stateRise = 1'b0;
    if(CsrPlugin_timeout_counter_willOverflow) begin
      CsrPlugin_timeout_stateRise = (! CsrPlugin_timeout_state);
    end
    if(when_CsrPlugin_l753) begin
      CsrPlugin_timeout_stateRise = 1'b0;
    end
    if(CsrPlugin_inject_cmd_valid) begin
      CsrPlugin_timeout_stateRise = 1'b0;
    end
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
        CsrPlugin_timeout_stateRise = 1'b0;
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_timeout_counter_willClear = 1'b0;
    if(when_CsrPlugin_l753) begin
      CsrPlugin_timeout_counter_willClear = 1'b1;
    end
    if(CsrPlugin_inject_cmd_valid) begin
      CsrPlugin_timeout_counter_willClear = 1'b1;
    end
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
        CsrPlugin_timeout_counter_willClear = 1'b1;
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrPlugin_timeout_counter_willOverflowIfInc = (CsrPlugin_timeout_counter_value == 3'b110);
  assign CsrPlugin_timeout_counter_willOverflow = (CsrPlugin_timeout_counter_willOverflowIfInc && CsrPlugin_timeout_counter_willIncrement);
  always @(*) begin
    if(CsrPlugin_timeout_counter_willOverflow) begin
      CsrPlugin_timeout_counter_valueNext = 3'b000;
    end else begin
      CsrPlugin_timeout_counter_valueNext = (CsrPlugin_timeout_counter_value + _zz_CsrPlugin_timeout_counter_valueNext);
    end
    if(CsrPlugin_timeout_counter_willClear) begin
      CsrPlugin_timeout_counter_valueNext = 3'b000;
    end
  end

  assign CsrPlugin_timeout_counter_willIncrement = 1'b1;
  assign when_CsrPlugin_l753 = (|{writeBack_arbitration_isValid,{memory_arbitration_isValid,execute_arbitration_isValid}});
  always @(*) begin
    _zz_debugBus_hartToDm_valid = 1'b0;
    if(execute_CsrPlugin_csr_1972) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_debugBus_hartToDm_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    debugBus_hartToDm_valid = _zz_debugBus_hartToDm_valid;
    if(fpuAccess_readDataValid) begin
      debugBus_hartToDm_valid = 1'b1;
    end
  end

  always @(*) begin
    debugBus_hartToDm_payload_address = 4'b0000;
    if(fpuAccess_readDataValid) begin
      debugBus_hartToDm_payload_address = {3'd0, fpuAccess_readDataChunk};
    end
  end

  always @(*) begin
    debugBus_hartToDm_payload_data = execute_SRC1;
    if(fpuAccess_readDataValid) begin
      debugBus_hartToDm_payload_data = fpuAccess_readData;
    end
  end

  assign when_CsrPlugin_l768 = (debugBus_dmToHart_valid && (debugBus_dmToHart_payload_op == DebugDmToHartOp_DATA));
  assign _zz_6 = ({1'd0,1'b1} <<< _zz__zz_6);
  assign CsrPlugin_inject_cmd_valid = (debugBus_dmToHart_valid && (((debugBus_dmToHart_payload_op == DebugDmToHartOp_EXECUTE) || (debugBus_dmToHart_payload_op == DebugDmToHartOp_REG_READ)) || (debugBus_dmToHart_payload_op == DebugDmToHartOp_REG_WRITE)));
  assign CsrPlugin_inject_cmd_payload_op = debugBus_dmToHart_payload_op;
  assign CsrPlugin_inject_cmd_payload_address = debugBus_dmToHart_payload_address;
  assign CsrPlugin_inject_cmd_payload_data = debugBus_dmToHart_payload_data;
  assign CsrPlugin_inject_cmd_payload_size = debugBus_dmToHart_payload_size;
  assign CsrPlugin_inject_cmd_toStream_valid = CsrPlugin_inject_cmd_valid;
  assign CsrPlugin_inject_cmd_toStream_payload_op = CsrPlugin_inject_cmd_payload_op;
  assign CsrPlugin_inject_cmd_toStream_payload_address = CsrPlugin_inject_cmd_payload_address;
  assign CsrPlugin_inject_cmd_toStream_payload_data = CsrPlugin_inject_cmd_payload_data;
  assign CsrPlugin_inject_cmd_toStream_payload_size = CsrPlugin_inject_cmd_payload_size;
  always @(*) begin
    CsrPlugin_inject_cmd_toStream_ready = CsrPlugin_inject_buffer_ready;
    if(when_Stream_l375_1) begin
      CsrPlugin_inject_cmd_toStream_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! CsrPlugin_inject_buffer_valid);
  assign CsrPlugin_inject_buffer_valid = CsrPlugin_inject_cmd_toStream_rValid;
  assign CsrPlugin_inject_buffer_payload_op = CsrPlugin_inject_cmd_toStream_rData_op;
  assign CsrPlugin_inject_buffer_payload_address = CsrPlugin_inject_cmd_toStream_rData_address;
  assign CsrPlugin_inject_buffer_payload_data = CsrPlugin_inject_cmd_toStream_rData_data;
  assign CsrPlugin_inject_buffer_payload_size = CsrPlugin_inject_cmd_toStream_rData_size;
  assign CsrPlugin_injectionPort_valid = (CsrPlugin_inject_buffer_valid && (CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_EXECUTE));
  assign CsrPlugin_injectionPort_payload = CsrPlugin_inject_buffer_payload_data;
  assign CsrPlugin_injectionPort_fire = (CsrPlugin_injectionPort_valid && CsrPlugin_injectionPort_ready);
  always @(*) begin
    CsrPlugin_inject_buffer_ready = CsrPlugin_injectionPort_fire;
    if(fpuAccess_done) begin
      CsrPlugin_inject_buffer_ready = 1'b1;
    end
  end

  assign fpuAccess_start = (CsrPlugin_inject_buffer_valid && ((CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_REG_READ) || (CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_REG_WRITE)));
  assign fpuAccess_regId = CsrPlugin_inject_buffer_payload_address;
  assign fpuAccess_write = (CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_REG_WRITE);
  assign fpuAccess_writeData = {CsrPlugin_dataCsrw_value_1,CsrPlugin_dataCsrw_value_0};
  assign fpuAccess_size = CsrPlugin_inject_buffer_payload_size;
  assign debugBus_regSuccess = fpuAccess_done;
  assign when_CsrPlugin_l804 = (CsrPlugin_inject_cmd_valid && (debugBus_dmToHart_payload_op == DebugDmToHartOp_EXECUTE));
  assign when_CsrPlugin_l804_1 = (((debugBus_exception || debugBus_commit) || debugBus_ebreak) || debugBus_redo);
  assign debugBus_redo = (CsrPlugin_inject_pending && CsrPlugin_timeout_state);
  assign CsrPlugin_dcsr_nmip = 1'b0;
  assign CsrPlugin_dcsr_mprven = 1'b1;
  assign CsrPlugin_dcsr_xdebugver = 4'b0100;
  assign CsrPlugin_dcsr_stepLogic_wantExit = 1'b0;
  always @(*) begin
    CsrPlugin_dcsr_stepLogic_wantStart = 1'b0;
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
      end
      default : begin
        CsrPlugin_dcsr_stepLogic_wantStart = 1'b1;
      end
    endcase
  end

  assign CsrPlugin_dcsr_stepLogic_wantKill = 1'b0;
  always @(*) begin
    CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_stateReg;
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
        if(when_CsrPlugin_l830) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_SINGLE;
        end
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
        if(when_CsrPlugin_l836) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1;
        end
        if(decode_arbitration_isFiring) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1;
        end
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
        if(when_CsrPlugin_l848) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_SINGLE;
        end
      end
      default : begin
      end
    endcase
    if(CsrPlugin_enterHalt) begin
      CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_IDLE;
    end
    if(CsrPlugin_dcsr_stepLogic_wantStart) begin
      CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_IDLE;
    end
    if(CsrPlugin_dcsr_stepLogic_wantKill) begin
      CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_BOOT;
    end
  end

  assign when_CsrPlugin_l830 = (CsrPlugin_dcsr_step && debugBus_resume_rsp_valid);
  assign when_CsrPlugin_l848 = ((! CsrPlugin_doHalt) && CsrPlugin_timeout_state);
  assign when_CsrPlugin_l880 = ((debugMode || CsrPlugin_dcsr_step) || debugBus_haltReq);
  assign CsrPlugin_misa_base = 2'b01;
  assign CsrPlugin_misa_extensions = 26'h000112d;
  assign _zz_when_CsrPlugin_l1446 = (CsrPlugin_mip_MTIP && CsrPlugin_mie_MTIE);
  assign _zz_when_CsrPlugin_l1446_1 = (CsrPlugin_mip_MSIP && CsrPlugin_mie_MSIE);
  assign _zz_when_CsrPlugin_l1446_2 = (CsrPlugin_mip_MEIP && CsrPlugin_mie_MEIE);
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped = 2'b11;
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege = ((CsrPlugin_privilege < CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped) ? CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped : CsrPlugin_privilege);
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code = {decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid};
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1[0];
  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_decode = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_execute = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_memory = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
    if(memory_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
    if(DBusCachedPlugin_exceptionBus_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b1;
    end
    if(writeBack_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b0;
    end
  end

  assign when_CsrPlugin_l1403 = (! decode_arbitration_isStuck);
  assign when_CsrPlugin_l1403_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1403_2 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l1403_3 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l1416 = (|{CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValids_memory,{CsrPlugin_exceptionPortCtrl_exceptionValids_execute,CsrPlugin_exceptionPortCtrl_exceptionValids_decode}}});
  assign CsrPlugin_exceptionPendings_0 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  assign CsrPlugin_exceptionPendings_1 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  assign CsrPlugin_exceptionPendings_2 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  assign CsrPlugin_exceptionPendings_3 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  assign when_CsrPlugin_l1440 = (CsrPlugin_mstatus_MIE || (CsrPlugin_privilege < 2'b11));
  assign when_CsrPlugin_l1446 = ((_zz_when_CsrPlugin_l1446 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l1446_1 = ((_zz_when_CsrPlugin_l1446_1 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l1446_2 = ((_zz_when_CsrPlugin_l1446_2 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l1459 = (CsrPlugin_dcsr_step && (! CsrPlugin_dcsr_stepie));
  assign CsrPlugin_exception = (CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack && CsrPlugin_allowException);
  assign CsrPlugin_lastStageWasWfi = 1'b0;
  assign CsrPlugin_pipelineLiberator_active = ((CsrPlugin_interrupt_valid && CsrPlugin_allowInterrupts) && decode_arbitration_isValid);
  assign when_CsrPlugin_l1479 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1479_1 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l1479_2 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l1484 = ((! CsrPlugin_pipelineLiberator_active) || decode_arbitration_removeIt);
  always @(*) begin
    CsrPlugin_pipelineLiberator_done = CsrPlugin_pipelineLiberator_pcValids_2;
    if(when_CsrPlugin_l1490) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
    if(CsrPlugin_hadException) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
  end

  assign when_CsrPlugin_l1490 = (|{CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory,CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute}});
  assign CsrPlugin_interruptJump = ((CsrPlugin_interrupt_valid && CsrPlugin_pipelineLiberator_done) && CsrPlugin_allowInterrupts);
  assign debugBus_commit = (debugMode && writeBack_arbitration_isFiring);
  always @(*) begin
    debugBus_exception = (debugMode && CsrPlugin_hadException);
    if(when_CsrPlugin_l1534) begin
      if(!when_CsrPlugin_l1542) begin
        if(!when_CsrPlugin_l1572) begin
          debugBus_exception = (! CsrPlugin_trapCauseEbreakDebug);
        end
      end
    end
  end

  always @(*) begin
    debugBus_ebreak = 1'b0;
    if(when_CsrPlugin_l1534) begin
      if(!when_CsrPlugin_l1542) begin
        if(!when_CsrPlugin_l1572) begin
          debugBus_ebreak = CsrPlugin_trapCauseEbreakDebug;
        end
      end
    end
  end

  always @(*) begin
    CsrPlugin_targetPrivilege = CsrPlugin_interrupt_targetPrivilege;
    if(CsrPlugin_hadException) begin
      CsrPlugin_targetPrivilege = CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
    end
  end

  always @(*) begin
    CsrPlugin_trapCause = CsrPlugin_interrupt_code;
    if(CsrPlugin_hadException) begin
      CsrPlugin_trapCause = CsrPlugin_exceptionPortCtrl_exceptionContext_code;
    end
  end

  always @(*) begin
    CsrPlugin_trapCauseEbreakDebug = 1'b0;
    if(CsrPlugin_hadException) begin
      if(when_CsrPlugin_l1517) begin
        if(debugMode) begin
          CsrPlugin_trapCauseEbreakDebug = 1'b1;
        end
        if(when_CsrPlugin_l1519) begin
          CsrPlugin_trapCauseEbreakDebug = 1'b1;
        end
      end
    end
  end

  assign when_CsrPlugin_l1517 = (CsrPlugin_exceptionPortCtrl_exceptionContext_code == 4'b0011);
  assign when_CsrPlugin_l1519 = ((CsrPlugin_privilege == 2'b11) && CsrPlugin_dcsr_ebreakm);
  always @(*) begin
    CsrPlugin_xtvec_mode = 2'bxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_mode = CsrPlugin_mtvec_mode;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_xtvec_base = 30'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_base = CsrPlugin_mtvec_base;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_trapEnterDebug = 1'b0;
    if(when_CsrPlugin_l1533) begin
      CsrPlugin_trapEnterDebug = 1'b1;
    end
  end

  assign when_CsrPlugin_l1533 = (((CsrPlugin_doHalt || CsrPlugin_trapCauseEbreakDebug) || ((! CsrPlugin_hadException) && CsrPlugin_doHalt)) || (! CsrPlugin_running));
  assign when_CsrPlugin_l1534 = (CsrPlugin_hadException || CsrPlugin_interruptJump);
  assign when_CsrPlugin_l1542 = (! CsrPlugin_trapEnterDebug);
  assign when_CsrPlugin_l1572 = (! debugMode);
  assign when_CsrPlugin_l1600 = (writeBack_arbitration_isValid && (writeBack_ENV_CTRL == EnvCtrlEnum_XRET));
  assign switch_CsrPlugin_l1604 = writeBack_INSTRUCTION[29 : 28];
  assign when_CsrPlugin_l1612 = (CsrPlugin_mstatus_MPP < 2'b11);
  assign contextSwitching = CsrPlugin_jumpInterface_valid;
  assign when_CsrPlugin_l1671 = (|{(writeBack_arbitration_isValid && (writeBack_ENV_CTRL == EnvCtrlEnum_XRET)),{(memory_arbitration_isValid && (memory_ENV_CTRL == EnvCtrlEnum_XRET)),(execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_XRET))}});
  assign execute_CsrPlugin_blockedBySideEffects = ((|{writeBack_arbitration_isValid,memory_arbitration_isValid}) || 1'b0);
  always @(*) begin
    execute_CsrPlugin_illegalAccess = 1'b1;
    if(execute_CsrPlugin_csr_1972) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_1969) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_1968) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_3857) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3858) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3859) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3860) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_769) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_768) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_836) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_772) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_773) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_833) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_832) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_834) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_835) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_2) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_1) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_256) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(CsrPlugin_csrMapping_allowCsrSignal) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(when_CsrPlugin_l1863) begin
      execute_CsrPlugin_illegalAccess = 1'b1;
    end
    if(when_CsrPlugin_l1869) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_illegalInstruction = 1'b0;
    if(when_CsrPlugin_l1691) begin
      if(when_CsrPlugin_l1692) begin
        execute_CsrPlugin_illegalInstruction = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrPlugin_selfException_valid = 1'b0;
    if(when_CsrPlugin_l1684) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
    if(when_CsrPlugin_l1699) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
    if(when_CsrPlugin_l1709) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_selfException_payload_code = 4'bxxxx;
    if(when_CsrPlugin_l1684) begin
      CsrPlugin_selfException_payload_code = 4'b0010;
    end
    if(when_CsrPlugin_l1699) begin
      case(CsrPlugin_privilege)
        2'b00 : begin
          CsrPlugin_selfException_payload_code = 4'b1000;
        end
        default : begin
          CsrPlugin_selfException_payload_code = 4'b1011;
        end
      endcase
    end
    if(when_CsrPlugin_l1709) begin
      CsrPlugin_selfException_payload_code = 4'b0011;
    end
  end

  assign CsrPlugin_selfException_payload_badAddr = execute_INSTRUCTION;
  assign when_CsrPlugin_l1684 = (execute_CsrPlugin_illegalAccess || execute_CsrPlugin_illegalInstruction);
  assign when_CsrPlugin_l1691 = (execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_XRET));
  assign when_CsrPlugin_l1692 = (CsrPlugin_privilege < execute_INSTRUCTION[29 : 28]);
  assign when_CsrPlugin_l1699 = (execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_ECALL));
  assign when_CsrPlugin_l1709 = ((execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_EBREAK)) && CsrPlugin_allowEbreakException);
  always @(*) begin
    execute_CsrPlugin_writeInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_WRITE_OPCODE);
    if(when_CsrPlugin_l1863) begin
      execute_CsrPlugin_writeInstruction = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_readInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_READ_OPCODE);
    if(when_CsrPlugin_l1863) begin
      execute_CsrPlugin_readInstruction = 1'b0;
    end
  end

  assign execute_CsrPlugin_writeEnable = (execute_CsrPlugin_writeInstruction && (! execute_arbitration_isStuck));
  assign execute_CsrPlugin_readEnable = (execute_CsrPlugin_readInstruction && (! execute_arbitration_isStuck));
  assign CsrPlugin_csrMapping_hazardFree = (! execute_CsrPlugin_blockedBySideEffects);
  assign execute_CsrPlugin_readToWriteData = CsrPlugin_csrMapping_readDataSignal;
  assign switch_Misc_l241_3 = execute_INSTRUCTION[13];
  always @(*) begin
    case(switch_Misc_l241_3)
      1'b0 : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = execute_SRC1;
      end
      default : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = (execute_INSTRUCTION[12] ? (execute_CsrPlugin_readToWriteData & (~ execute_SRC1)) : (execute_CsrPlugin_readToWriteData | execute_SRC1));
      end
    endcase
  end

  assign CsrPlugin_csrMapping_writeDataSignal = _zz_CsrPlugin_csrMapping_writeDataSignal;
  assign when_CsrPlugin_l1731 = (execute_arbitration_isValid && execute_IS_CSR);
  assign when_CsrPlugin_l1735 = (execute_arbitration_isValid && (execute_IS_CSR || 1'b0));
  assign execute_CsrPlugin_csrAddress = execute_INSTRUCTION[31 : 20];
  assign execute_BranchPlugin_eq = (execute_SRC1 == execute_SRC2);
  assign switch_Misc_l241_4 = execute_INSTRUCTION[14 : 12];
  always @(*) begin
    case(switch_Misc_l241_4)
      3'b000 : begin
        _zz_execute_BRANCH_DO = execute_BranchPlugin_eq;
      end
      3'b001 : begin
        _zz_execute_BRANCH_DO = (! execute_BranchPlugin_eq);
      end
      3'b101 : begin
        _zz_execute_BRANCH_DO = (! execute_SRC_LESS);
      end
      3'b111 : begin
        _zz_execute_BRANCH_DO = (! execute_SRC_LESS);
      end
      default : begin
        _zz_execute_BRANCH_DO = execute_SRC_LESS;
      end
    endcase
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : begin
        _zz_execute_BRANCH_DO_1 = 1'b0;
      end
      BranchCtrlEnum_JAL : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      BranchCtrlEnum_JALR : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      default : begin
        _zz_execute_BRANCH_DO_1 = _zz_execute_BRANCH_DO;
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src1 = ((execute_BRANCH_CTRL == BranchCtrlEnum_JALR) ? execute_RS1 : execute_PC);
  assign _zz_execute_BranchPlugin_branch_src2 = _zz__zz_execute_BranchPlugin_branch_src2[19];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_1[10] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[9] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[8] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[7] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[6] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[5] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[4] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[3] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[2] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[1] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[0] = _zz_execute_BranchPlugin_branch_src2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_2 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_3[19] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[18] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[17] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[16] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[15] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[14] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[13] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[12] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[11] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[10] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[9] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[8] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[7] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[6] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[5] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[4] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[3] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[2] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[1] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[0] = _zz_execute_BranchPlugin_branch_src2_2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_4 = _zz__zz_execute_BranchPlugin_branch_src2_4[11];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_5[18] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[17] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[16] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[15] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[14] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[13] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[12] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[11] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[10] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[9] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[8] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[7] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[6] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[5] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[4] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[3] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[2] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[1] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[0] = _zz_execute_BranchPlugin_branch_src2_4;
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_JAL : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_1,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]}},1'b0};
      end
      BranchCtrlEnum_JALR : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {_zz_execute_BranchPlugin_branch_src2_3,execute_INSTRUCTION[31 : 20]};
      end
      default : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_5,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]}},1'b0};
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src2 = _zz_execute_BranchPlugin_branch_src2_6;
  assign execute_BranchPlugin_branchAdder = (execute_BranchPlugin_branch_src1 + execute_BranchPlugin_branch_src2);
  assign BranchPlugin_jumpInterface_valid = ((memory_arbitration_isValid && memory_BRANCH_DO) && (! 1'b0));
  assign BranchPlugin_jumpInterface_payload = memory_BRANCH_CALC;
  assign when_MulPlugin_l65 = ((execute_arbitration_isValid && execute_IS_MUL) && (execute_MulPlugin_delayLogic_counter != 1'b1));
  assign when_MulPlugin_l70 = ((! execute_arbitration_isStuck) || execute_arbitration_isStuckByOthers);
  assign execute_MulPlugin_a = execute_RS1;
  assign execute_MulPlugin_b = execute_RS2;
  assign switch_MulPlugin_l87 = execute_INSTRUCTION[13 : 12];
  always @(*) begin
    case(switch_MulPlugin_l87)
      2'b01 : begin
        execute_MulPlugin_aSigned = 1'b1;
      end
      2'b10 : begin
        execute_MulPlugin_aSigned = 1'b1;
      end
      default : begin
        execute_MulPlugin_aSigned = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(switch_MulPlugin_l87)
      2'b01 : begin
        execute_MulPlugin_bSigned = 1'b1;
      end
      2'b10 : begin
        execute_MulPlugin_bSigned = 1'b0;
      end
      default : begin
        execute_MulPlugin_bSigned = 1'b0;
      end
    endcase
  end

  assign execute_MulPlugin_aULow = execute_MulPlugin_a[15 : 0];
  assign execute_MulPlugin_bULow = execute_MulPlugin_b[15 : 0];
  assign execute_MulPlugin_aSLow = {1'b0,execute_MulPlugin_a[15 : 0]};
  assign execute_MulPlugin_bSLow = {1'b0,execute_MulPlugin_b[15 : 0]};
  assign execute_MulPlugin_aHigh = {(execute_MulPlugin_aSigned && execute_MulPlugin_a[31]),execute_MulPlugin_a[31 : 16]};
  assign execute_MulPlugin_bHigh = {(execute_MulPlugin_bSigned && execute_MulPlugin_b[31]),execute_MulPlugin_b[31 : 16]};
  assign writeBack_MulPlugin_result = ($signed(_zz_writeBack_MulPlugin_result) + $signed(_zz_writeBack_MulPlugin_result_1));
  assign when_MulPlugin_l147 = (writeBack_arbitration_isValid && writeBack_IS_MUL);
  assign switch_MulPlugin_l148 = writeBack_INSTRUCTION[13 : 12];
  assign memory_MulDivIterativePlugin_frontendOk = 1'b1;
  always @(*) begin
    memory_MulDivIterativePlugin_div_counter_willIncrement = 1'b0;
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l132) begin
        memory_MulDivIterativePlugin_div_counter_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    memory_MulDivIterativePlugin_div_counter_willClear = 1'b0;
    if(when_MulDivIterativePlugin_l162) begin
      memory_MulDivIterativePlugin_div_counter_willClear = 1'b1;
    end
  end

  assign memory_MulDivIterativePlugin_div_counter_willOverflowIfInc = (memory_MulDivIterativePlugin_div_counter_value == 6'h21);
  assign memory_MulDivIterativePlugin_div_counter_willOverflow = (memory_MulDivIterativePlugin_div_counter_willOverflowIfInc && memory_MulDivIterativePlugin_div_counter_willIncrement);
  always @(*) begin
    if(memory_MulDivIterativePlugin_div_counter_willOverflow) begin
      memory_MulDivIterativePlugin_div_counter_valueNext = 6'h0;
    end else begin
      memory_MulDivIterativePlugin_div_counter_valueNext = (memory_MulDivIterativePlugin_div_counter_value + _zz_memory_MulDivIterativePlugin_div_counter_valueNext);
    end
    if(memory_MulDivIterativePlugin_div_counter_willClear) begin
      memory_MulDivIterativePlugin_div_counter_valueNext = 6'h0;
    end
  end

  assign when_MulDivIterativePlugin_l126 = (memory_MulDivIterativePlugin_div_counter_value == 6'h20);
  assign when_MulDivIterativePlugin_l126_1 = (! memory_arbitration_isStuck);
  assign when_MulDivIterativePlugin_l128 = (memory_arbitration_isValid && memory_IS_DIV);
  assign when_MulDivIterativePlugin_l129 = ((! memory_MulDivIterativePlugin_frontendOk) || (! memory_MulDivIterativePlugin_div_done));
  assign when_MulDivIterativePlugin_l132 = (memory_MulDivIterativePlugin_frontendOk && (! memory_MulDivIterativePlugin_div_done));
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted = memory_MulDivIterativePlugin_rs1[31 : 0];
  assign memory_MulDivIterativePlugin_div_stage_0_remainderShifted = {memory_MulDivIterativePlugin_accumulator[31 : 0],_zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted[31]};
  assign memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator = (memory_MulDivIterativePlugin_div_stage_0_remainderShifted - _zz_memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator);
  assign memory_MulDivIterativePlugin_div_stage_0_outRemainder = ((! memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator[32]) ? _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder : _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder_1);
  assign memory_MulDivIterativePlugin_div_stage_0_outNumerator = _zz_memory_MulDivIterativePlugin_div_stage_0_outNumerator[31:0];
  assign when_MulDivIterativePlugin_l151 = (memory_MulDivIterativePlugin_div_counter_value == 6'h20);
  assign _zz_memory_MulDivIterativePlugin_div_result = (memory_INSTRUCTION[13] ? memory_MulDivIterativePlugin_accumulator[31 : 0] : memory_MulDivIterativePlugin_rs1[31 : 0]);
  assign when_MulDivIterativePlugin_l162 = (! memory_arbitration_isStuck);
  assign _zz_memory_MulDivIterativePlugin_rs2 = (execute_RS2[31] && execute_IS_RS2_SIGNED);
  assign _zz_memory_MulDivIterativePlugin_rs1 = (1'b0 || ((execute_IS_DIV && execute_RS1[31]) && execute_IS_RS1_SIGNED));
  always @(*) begin
    _zz_memory_MulDivIterativePlugin_rs1_1[32] = (execute_IS_RS1_SIGNED && execute_RS1[31]);
    _zz_memory_MulDivIterativePlugin_rs1_1[31 : 0] = execute_RS1;
  end

  assign FpuPlugin_port_cmd_fire = (FpuPlugin_port_cmd_valid && FpuPlugin_port_cmd_ready);
  assign FpuPlugin_port_rsp_fire = (FpuPlugin_port_rsp_valid && FpuPlugin_port_rsp_ready);
  assign FpuPlugin_hasPending = (FpuPlugin_pendings != 6'h0);
  assign when_FpuPlugin_l215 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_NV);
  assign when_FpuPlugin_l216 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_DZ);
  assign when_FpuPlugin_l217 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_OF);
  assign when_FpuPlugin_l218 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_UF);
  assign when_FpuPlugin_l219 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_NX);
  assign FpuPlugin_csrActive = (execute_arbitration_isValid && execute_IS_CSR);
  assign when_FpuPlugin_l229 = (FpuPlugin_csrActive && FpuPlugin_hasPending);
  assign FpuPlugin_sd = (FpuPlugin_fs == 2'b11);
  assign when_FpuPlugin_l234 = (FpuPlugin_port_completion_valid && (FpuPlugin_port_completion_payload_written || (|{FpuPlugin_port_completion_payload_flags_NV,{FpuPlugin_port_completion_payload_flags_DZ,{FpuPlugin_port_completion_payload_flags_OF,{FpuPlugin_port_completion_payload_flags_UF,FpuPlugin_port_completion_payload_flags_NX}}}})));
  always @(*) begin
    _zz_when_FpuPlugin_l237 = 1'b0;
    if(execute_CsrPlugin_csr_2) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_when_FpuPlugin_l237 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_when_FpuPlugin_l237_1 = 1'b0;
    if(execute_CsrPlugin_csr_3) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_when_FpuPlugin_l237_1 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_when_FpuPlugin_l237_2 = 1'b0;
    if(execute_CsrPlugin_csr_1) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_when_FpuPlugin_l237_2 = 1'b1;
      end
    end
  end

  assign when_FpuPlugin_l237 = (|{_zz_when_FpuPlugin_l237_2,{_zz_when_FpuPlugin_l237_1,_zz_when_FpuPlugin_l237}});
  always @(*) begin
    FpuPlugin_accessFpuCsr = 1'b0;
    if(execute_CsrPlugin_csr_3) begin
      FpuPlugin_accessFpuCsr = 1'b1;
    end
    if(execute_CsrPlugin_csr_2) begin
      FpuPlugin_accessFpuCsr = 1'b1;
    end
    if(execute_CsrPlugin_csr_1) begin
      FpuPlugin_accessFpuCsr = 1'b1;
    end
  end

  assign when_FpuPlugin_l253 = ((FpuPlugin_accessFpuCsr && (FpuPlugin_fs == 2'b00)) && (! debugMode));
  always @(*) begin
    _zz_decode_FPU_FORKED = 1'b0;
    if(when_FpuPlugin_l350) begin
      _zz_decode_FPU_FORKED = 1'b1;
    end
  end

  assign decode_FpuPlugin_trap = (((_zz_decode_FPU_ENABLE && (FpuPlugin_fs == 2'b00)) && (! debugMode)) && (! (|{writeBack_arbitration_isValid,{memory_arbitration_isValid,execute_arbitration_isValid}})));
  assign when_FpuPlugin_l268 = (FpuPlugin_port_cmd_fire && (! _zz_decode_FPU_FORKED));
  assign when_FpuPlugin_l268_1 = (! decode_arbitration_isStuck);
  assign decode_FpuPlugin_hazard = ((FpuPlugin_pendings[5] || FpuPlugin_csrActive) || ((FpuPlugin_fs == 2'b00) && (! debugMode)));
  assign when_FpuPlugin_l272 = (! decode_LEGAL_INSTRUCTION);
  assign when_FpuPlugin_l273 = ((decode_arbitration_isValid && decode_FPU_ENABLE) && decode_FpuPlugin_hazard);
  assign FpuPlugin_port_cmd_isStall = (FpuPlugin_port_cmd_valid && (! FpuPlugin_port_cmd_ready));
  assign decode_FpuPlugin_iRoundMode = decode_INSTRUCTION[14 : 12];
  assign decode_FpuPlugin_roundMode = ((decode_INSTRUCTION[14 : 12] == 3'b111) ? FpuPlugin_rm : decode_INSTRUCTION[14 : 12]);
  always @(*) begin
    FpuPlugin_port_cmd_valid = (((decode_arbitration_isValid && decode_FPU_ENABLE) && (! decode_FpuPlugin_forked)) && (! decode_FpuPlugin_hazard));
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_valid = 1'b1;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_cmd_payload_opcode = decode_FPU_OPCODE;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        if(fpuAccess_write) begin
          FpuPlugin_port_cmd_payload_opcode = FpuOpcode_LOAD;
        end else begin
          FpuPlugin_port_cmd_payload_opcode = FpuOpcode_STORE;
        end
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign FpuPlugin_port_cmd_payload_arg = decode_FPU_ARG;
  assign FpuPlugin_port_cmd_payload_rs1 = decode_INSTRUCTION[19 : 15];
  always @(*) begin
    FpuPlugin_port_cmd_payload_rs2 = decode_INSTRUCTION[24 : 20];
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_payload_rs2 = fpuAccess_regId;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign FpuPlugin_port_cmd_payload_rs3 = decode_INSTRUCTION[31 : 27];
  always @(*) begin
    FpuPlugin_port_cmd_payload_rd = decode_INSTRUCTION[11 : 7];
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_payload_rd = fpuAccess_regId;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_cmd_payload_format = decode_FPU_FORMAT;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_payload_format = _zz_FpuPlugin_port_cmd_payload_format;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign _zz_FpuPlugin_port_cmd_payload_roundMode_1 = decode_FpuPlugin_roundMode;
  assign _zz_FpuPlugin_port_cmd_payload_roundMode = _zz_FpuPlugin_port_cmd_payload_roundMode_1;
  assign FpuPlugin_port_cmd_payload_roundMode = _zz_FpuPlugin_port_cmd_payload_roundMode;
  assign writeBack_FpuPlugin_isRsp = (writeBack_FPU_FORKED && writeBack_FPU_RSP);
  assign writeBack_FpuPlugin_isCommit = (writeBack_FPU_FORKED && writeBack_FPU_COMMIT);
  always @(*) begin
    writeBack_FpuPlugin_storeFormated = FpuPlugin_port_rsp_payload_value;
    if(when_FpuPlugin_l306) begin
      writeBack_FpuPlugin_storeFormated[63 : 32] = FpuPlugin_port_rsp_payload_value[31 : 0];
    end
  end

  assign when_FpuPlugin_l306 = (! writeBack_INSTRUCTION[12]);
  always @(*) begin
    FpuPlugin_port_rsp_ready = 1'b0;
    if(writeBack_FpuPlugin_isRsp) begin
      if(!when_FpuPlugin_l323) begin
        if(when_FpuPlugin_l325) begin
          FpuPlugin_port_rsp_ready = 1'b1;
        end
      end
    end
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
        FpuPlugin_port_rsp_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign DBusBypass0_value = writeBack_FpuPlugin_storeFormated;
  assign when_FpuPlugin_l315 = ((! writeBack_arbitration_isStuck) && (! writeBack_arbitration_removeIt));
  assign when_FpuPlugin_l318 = (FpuPlugin_port_rsp_payload_NV || FpuPlugin_port_rsp_payload_NX);
  assign when_FpuPlugin_l323 = (! FpuPlugin_port_rsp_valid);
  assign when_FpuPlugin_l325 = (! writeBack_arbitration_haltItself);
  assign writeBack_FpuPlugin_commit_valid = (writeBack_FpuPlugin_isCommit && (! writeBack_arbitration_isStuck));
  always @(*) begin
    writeBack_FpuPlugin_commit_payload_value[31 : 0] = (writeBack_FPU_COMMIT_LOAD ? _zz_writeBack_FpuPlugin_commit_payload_value[31 : 0] : writeBack_RS1);
    writeBack_FpuPlugin_commit_payload_value[63 : 32] = _zz_writeBack_FpuPlugin_commit_payload_value[63 : 32];
  end

  assign writeBack_FpuPlugin_commit_payload_write = (writeBack_arbitration_isValid && (! writeBack_arbitration_removeIt));
  assign writeBack_FpuPlugin_commit_payload_opcode = writeBack_FPU_OPCODE;
  assign writeBack_FpuPlugin_commit_payload_rd = writeBack_INSTRUCTION[11 : 7];
  assign when_FpuPlugin_l339 = (writeBack_FpuPlugin_isCommit && (! writeBack_FpuPlugin_commit_ready));
  assign writeBack_FpuPlugin_commit_ready = writeBack_FpuPlugin_commit_rValidN;
  assign writeBack_FpuPlugin_commit_s2mPipe_valid = (writeBack_FpuPlugin_commit_valid || (! writeBack_FpuPlugin_commit_rValidN));
  assign _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_opcode : writeBack_FpuPlugin_commit_rData_opcode);
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_opcode = _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_rd = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_rd : writeBack_FpuPlugin_commit_rData_rd);
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_write = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_write : writeBack_FpuPlugin_commit_rData_write);
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_value = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_value : writeBack_FpuPlugin_commit_rData_value);
  always @(*) begin
    FpuPlugin_port_commit_valid = writeBack_FpuPlugin_commit_s2mPipe_valid;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_valid = 1'b1;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign writeBack_FpuPlugin_commit_s2mPipe_ready = FpuPlugin_port_commit_ready;
  always @(*) begin
    FpuPlugin_port_commit_payload_opcode = writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_opcode = FpuOpcode_LOAD;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_commit_payload_rd = writeBack_FpuPlugin_commit_s2mPipe_payload_rd;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_rd = fpuAccess_regId;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_commit_payload_write = writeBack_FpuPlugin_commit_s2mPipe_payload_write;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_write = 1'b1;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_commit_payload_value = writeBack_FpuPlugin_commit_s2mPipe_payload_value;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_value = fpuAccess_writeData;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign FpuPlugin_wantExit = 1'b0;
  always @(*) begin
    FpuPlugin_wantStart = 1'b0;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
        FpuPlugin_wantStart = 1'b1;
      end
    endcase
  end

  assign FpuPlugin_wantKill = 1'b0;
  assign when_FpuPlugin_l350 = (! (FpuPlugin_stateReg == FpuPlugin_enumDef_IDLE));
  always @(*) begin
    fpuAccess_done = 1'b0;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
        fpuAccess_done = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fpuAccess_readDataValid = 1'b0;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
        fpuAccess_readDataValid = 1'b1;
      end
      FpuPlugin_enumDef_RSP_1 : begin
        fpuAccess_readDataValid = 1'b1;
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fpuAccess_readDataChunk = 1'bx;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
        fpuAccess_readDataChunk = 1'b0;
      end
      FpuPlugin_enumDef_RSP_1 : begin
        fpuAccess_readDataChunk = 1'b1;
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fpuAccess_readData = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
        fpuAccess_readData = FpuPlugin_port_rsp_payload_value[31 : 0];
      end
      FpuPlugin_enumDef_RSP_1 : begin
        fpuAccess_readData = FpuPlugin_port_rsp_payload_value[63 : 32];
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign when_CfuPlugin_l192 = (! execute_LEGAL_INSTRUCTION);
  assign execute_CfuPlugin_hazard = (|{(writeBack_arbitration_isValid && writeBack_HAS_SIDE_EFFECT),(memory_arbitration_isValid && memory_HAS_SIDE_EFFECT)});
  assign execute_CfuPlugin_scheduleWish = (execute_arbitration_isValid && execute_CfuPlugin_CFU_ENABLE);
  assign execute_CfuPlugin_schedule = (execute_CfuPlugin_scheduleWish && (! execute_CfuPlugin_hazard));
  assign when_CfuPlugin_l196 = (execute_CfuPlugin_scheduleWish && execute_CfuPlugin_hazard);
  assign CfuPlugin_bus_cmd_fire = (CfuPlugin_bus_cmd_valid && CfuPlugin_bus_cmd_ready);
  assign when_CfuPlugin_l199 = (! execute_arbitration_isStuck);
  assign CfuPlugin_bus_cmd_valid = ((execute_CfuPlugin_schedule || execute_CfuPlugin_hold) && (! execute_CfuPlugin_fired));
  assign when_CfuPlugin_l203 = (CfuPlugin_bus_cmd_valid && (! CfuPlugin_bus_cmd_ready));
  assign execute_CfuPlugin_functionsIds_0 = {execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[14 : 12]};
  assign CfuPlugin_bus_cmd_payload_function_id = execute_CfuPlugin_functionsIds_0;
  assign CfuPlugin_bus_cmd_payload_inputs_0 = execute_RS1;
  assign _zz_CfuPlugin_bus_cmd_payload_inputs_1 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[23] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[22] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[21] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[20] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[19] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[18] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[17] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[16] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[15] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[14] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[13] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[12] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[11] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[10] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[9] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[8] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[7] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[6] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[5] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[4] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[3] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[2] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[1] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[0] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
  end

  always @(*) begin
    case(execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : begin
        _zz_CfuPlugin_bus_cmd_payload_inputs_1_2 = execute_RS2;
      end
      default : begin
        _zz_CfuPlugin_bus_cmd_payload_inputs_1_2 = {_zz_CfuPlugin_bus_cmd_payload_inputs_1_1,execute_INSTRUCTION[31 : 24]};
      end
    endcase
  end

  assign CfuPlugin_bus_cmd_payload_inputs_1 = _zz_CfuPlugin_bus_cmd_payload_inputs_1_2;
  assign CfuPlugin_bus_rsp_ready = CfuPlugin_bus_rsp_rValidN;
  assign writeBack_CfuPlugin_rsp_valid = (CfuPlugin_bus_rsp_valid || (! CfuPlugin_bus_rsp_rValidN));
  assign writeBack_CfuPlugin_rsp_payload_outputs_0 = (CfuPlugin_bus_rsp_rValidN ? CfuPlugin_bus_rsp_payload_outputs_0 : CfuPlugin_bus_rsp_rData_outputs_0);
  always @(*) begin
    writeBack_CfuPlugin_rsp_ready = 1'b0;
    if(writeBack_CfuPlugin_CFU_IN_FLIGHT) begin
      writeBack_CfuPlugin_rsp_ready = (! writeBack_arbitration_isStuckByOthers);
    end
  end

  assign when_CfuPlugin_l239 = (! writeBack_CfuPlugin_rsp_valid);
  always @(*) begin
    _zz_decode_RS2_3[0] = memory_SHIFT_RIGHT[31];
    _zz_decode_RS2_3[1] = memory_SHIFT_RIGHT[30];
    _zz_decode_RS2_3[2] = memory_SHIFT_RIGHT[29];
    _zz_decode_RS2_3[3] = memory_SHIFT_RIGHT[28];
    _zz_decode_RS2_3[4] = memory_SHIFT_RIGHT[27];
    _zz_decode_RS2_3[5] = memory_SHIFT_RIGHT[26];
    _zz_decode_RS2_3[6] = memory_SHIFT_RIGHT[25];
    _zz_decode_RS2_3[7] = memory_SHIFT_RIGHT[24];
    _zz_decode_RS2_3[8] = memory_SHIFT_RIGHT[23];
    _zz_decode_RS2_3[9] = memory_SHIFT_RIGHT[22];
    _zz_decode_RS2_3[10] = memory_SHIFT_RIGHT[21];
    _zz_decode_RS2_3[11] = memory_SHIFT_RIGHT[20];
    _zz_decode_RS2_3[12] = memory_SHIFT_RIGHT[19];
    _zz_decode_RS2_3[13] = memory_SHIFT_RIGHT[18];
    _zz_decode_RS2_3[14] = memory_SHIFT_RIGHT[17];
    _zz_decode_RS2_3[15] = memory_SHIFT_RIGHT[16];
    _zz_decode_RS2_3[16] = memory_SHIFT_RIGHT[15];
    _zz_decode_RS2_3[17] = memory_SHIFT_RIGHT[14];
    _zz_decode_RS2_3[18] = memory_SHIFT_RIGHT[13];
    _zz_decode_RS2_3[19] = memory_SHIFT_RIGHT[12];
    _zz_decode_RS2_3[20] = memory_SHIFT_RIGHT[11];
    _zz_decode_RS2_3[21] = memory_SHIFT_RIGHT[10];
    _zz_decode_RS2_3[22] = memory_SHIFT_RIGHT[9];
    _zz_decode_RS2_3[23] = memory_SHIFT_RIGHT[8];
    _zz_decode_RS2_3[24] = memory_SHIFT_RIGHT[7];
    _zz_decode_RS2_3[25] = memory_SHIFT_RIGHT[6];
    _zz_decode_RS2_3[26] = memory_SHIFT_RIGHT[5];
    _zz_decode_RS2_3[27] = memory_SHIFT_RIGHT[4];
    _zz_decode_RS2_3[28] = memory_SHIFT_RIGHT[3];
    _zz_decode_RS2_3[29] = memory_SHIFT_RIGHT[2];
    _zz_decode_RS2_3[30] = memory_SHIFT_RIGHT[1];
    _zz_decode_RS2_3[31] = memory_SHIFT_RIGHT[0];
  end

  assign when_Pipeline_l124 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_1 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_2 = ((! writeBack_arbitration_isStuck) && (! CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack));
  assign when_Pipeline_l124_3 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_4 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_5 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_6 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_7 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_8 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_9 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_10 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_11 = (! execute_arbitration_isStuck);
  assign _zz_decode_SRC1_CTRL = _zz_decode_SRC1_CTRL_1;
  assign when_Pipeline_l124_12 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_13 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_14 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_15 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_CTRL_1 = decode_ALU_CTRL;
  assign _zz_decode_ALU_CTRL = _zz_decode_ALU_CTRL_1;
  assign when_Pipeline_l124_16 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_CTRL = decode_to_execute_ALU_CTRL;
  assign _zz_decode_SRC2_CTRL = _zz_decode_SRC2_CTRL_1;
  assign when_Pipeline_l124_17 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_18 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_19 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_20 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_21 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_22 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_23 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_24 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_25 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_26 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_27 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_28 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_29 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_30 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_31 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_32 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_33 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_34 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_35 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_36 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_37 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_38 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_39 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ENV_CTRL_1 = decode_ENV_CTRL;
  assign _zz_execute_to_memory_ENV_CTRL_1 = execute_ENV_CTRL;
  assign _zz_memory_to_writeBack_ENV_CTRL_1 = memory_ENV_CTRL;
  assign _zz_decode_ENV_CTRL = _zz_decode_ENV_CTRL_1;
  assign when_Pipeline_l124_40 = (! execute_arbitration_isStuck);
  assign _zz_execute_ENV_CTRL = decode_to_execute_ENV_CTRL;
  assign when_Pipeline_l124_41 = (! memory_arbitration_isStuck);
  assign _zz_memory_ENV_CTRL = execute_to_memory_ENV_CTRL;
  assign when_Pipeline_l124_42 = (! writeBack_arbitration_isStuck);
  assign _zz_writeBack_ENV_CTRL = memory_to_writeBack_ENV_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL_1 = decode_BRANCH_CTRL;
  assign _zz_decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL_1;
  assign when_Pipeline_l124_43 = (! execute_arbitration_isStuck);
  assign _zz_execute_BRANCH_CTRL = decode_to_execute_BRANCH_CTRL;
  assign when_Pipeline_l124_44 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_45 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_46 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_47 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_48 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_49 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_50 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_51 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_52 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_53 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_54 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_55 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_56 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_57 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_FPU_OPCODE_1 = decode_FPU_OPCODE;
  assign _zz_execute_to_memory_FPU_OPCODE_1 = execute_FPU_OPCODE;
  assign _zz_memory_to_writeBack_FPU_OPCODE_1 = memory_FPU_OPCODE;
  assign _zz_decode_FPU_OPCODE = _zz_decode_FPU_OPCODE_1;
  assign when_Pipeline_l124_58 = (! execute_arbitration_isStuck);
  assign _zz_execute_FPU_OPCODE = decode_to_execute_FPU_OPCODE;
  assign when_Pipeline_l124_59 = (! memory_arbitration_isStuck);
  assign _zz_memory_FPU_OPCODE = execute_to_memory_FPU_OPCODE;
  assign when_Pipeline_l124_60 = (! writeBack_arbitration_isStuck);
  assign _zz_writeBack_FPU_OPCODE = memory_to_writeBack_FPU_OPCODE;
  assign _zz_decode_FPU_FORMAT = _zz_decode_FPU_FORMAT_1;
  assign when_Pipeline_l124_61 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1 = decode_CfuPlugin_CFU_INPUT_2_KIND;
  assign _zz_decode_CfuPlugin_CFU_INPUT_2_KIND = _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1;
  assign when_Pipeline_l124_62 = (! execute_arbitration_isStuck);
  assign _zz_execute_CfuPlugin_CFU_INPUT_2_KIND = decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL_1 = decode_ALU_BITWISE_CTRL;
  assign _zz_decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL_1;
  assign when_Pipeline_l124_63 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_BITWISE_CTRL = decode_to_execute_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL_1 = decode_SHIFT_CTRL;
  assign _zz_execute_to_memory_SHIFT_CTRL_1 = execute_SHIFT_CTRL;
  assign _zz_decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL_1;
  assign when_Pipeline_l124_64 = (! execute_arbitration_isStuck);
  assign _zz_execute_SHIFT_CTRL = decode_to_execute_SHIFT_CTRL;
  assign when_Pipeline_l124_65 = (! memory_arbitration_isStuck);
  assign _zz_memory_SHIFT_CTRL = execute_to_memory_SHIFT_CTRL;
  assign when_Pipeline_l124_66 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_67 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_68 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_69 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_70 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_71 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_72 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_73 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_74 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_75 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_76 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_77 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_78 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_79 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_80 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_81 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_82 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_83 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_84 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_85 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_86 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_87 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_88 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_89 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_90 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_91 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_92 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_93 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_94 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_95 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_96 = (! writeBack_arbitration_isStuck);
  assign decode_arbitration_isFlushed = ((|{writeBack_arbitration_flushNext,{memory_arbitration_flushNext,execute_arbitration_flushNext}}) || (|{writeBack_arbitration_flushIt,{memory_arbitration_flushIt,{execute_arbitration_flushIt,decode_arbitration_flushIt}}}));
  assign execute_arbitration_isFlushed = ((|{writeBack_arbitration_flushNext,memory_arbitration_flushNext}) || (|{writeBack_arbitration_flushIt,{memory_arbitration_flushIt,execute_arbitration_flushIt}}));
  assign memory_arbitration_isFlushed = ((|writeBack_arbitration_flushNext) || (|{writeBack_arbitration_flushIt,memory_arbitration_flushIt}));
  assign writeBack_arbitration_isFlushed = (1'b0 || (|writeBack_arbitration_flushIt));
  assign decode_arbitration_isStuckByOthers = (decode_arbitration_haltByOther || (((1'b0 || execute_arbitration_isStuck) || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign decode_arbitration_isStuck = (decode_arbitration_haltItself || decode_arbitration_isStuckByOthers);
  assign decode_arbitration_isMoving = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign decode_arbitration_isFiring = ((decode_arbitration_isValid && (! decode_arbitration_isStuck)) && (! decode_arbitration_removeIt));
  assign execute_arbitration_isStuckByOthers = (execute_arbitration_haltByOther || ((1'b0 || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign execute_arbitration_isStuck = (execute_arbitration_haltItself || execute_arbitration_isStuckByOthers);
  assign execute_arbitration_isMoving = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign execute_arbitration_isFiring = ((execute_arbitration_isValid && (! execute_arbitration_isStuck)) && (! execute_arbitration_removeIt));
  assign memory_arbitration_isStuckByOthers = (memory_arbitration_haltByOther || (1'b0 || writeBack_arbitration_isStuck));
  assign memory_arbitration_isStuck = (memory_arbitration_haltItself || memory_arbitration_isStuckByOthers);
  assign memory_arbitration_isMoving = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  assign memory_arbitration_isFiring = ((memory_arbitration_isValid && (! memory_arbitration_isStuck)) && (! memory_arbitration_removeIt));
  assign writeBack_arbitration_isStuckByOthers = (writeBack_arbitration_haltByOther || 1'b0);
  assign writeBack_arbitration_isStuck = (writeBack_arbitration_haltItself || writeBack_arbitration_isStuckByOthers);
  assign writeBack_arbitration_isMoving = ((! writeBack_arbitration_isStuck) && (! writeBack_arbitration_removeIt));
  assign writeBack_arbitration_isFiring = ((writeBack_arbitration_isValid && (! writeBack_arbitration_isStuck)) && (! writeBack_arbitration_removeIt));
  assign when_Pipeline_l151 = ((! execute_arbitration_isStuck) || execute_arbitration_removeIt);
  assign when_Pipeline_l154 = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign when_Pipeline_l151_1 = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  assign when_Pipeline_l154_1 = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign when_Pipeline_l151_2 = ((! writeBack_arbitration_isStuck) || writeBack_arbitration_removeIt);
  assign when_Pipeline_l154_2 = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  always @(*) begin
    CsrPlugin_injectionPort_ready = 1'b0;
    case(IBusCachedPlugin_injector_port_state)
      3'b100 : begin
        CsrPlugin_injectionPort_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign when_Fetcher_l373 = (IBusCachedPlugin_injector_port_state != 3'b000);
  assign when_Fetcher_l391 = (! decode_arbitration_isStuck);
  assign when_Fetcher_l411 = (IBusCachedPlugin_injector_port_state != 3'b000);
  assign when_CsrPlugin_l1813 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_2 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_3 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_4 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_5 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_6 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_7 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_8 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_9 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_10 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_11 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_12 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_13 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_14 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_15 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_16 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_17 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_18 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_19 = (! execute_arbitration_isStuck);
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit = 32'h0;
    if(execute_CsrPlugin_csr_1972) begin
      _zz_CsrPlugin_csrMapping_readDataInit[31 : 0] = CsrPlugin_dataCsrw_value_0;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_1 = 32'h0;
    if(execute_CsrPlugin_csr_1969) begin
      _zz_CsrPlugin_csrMapping_readDataInit_1[31 : 0] = CsrPlugin_dpc;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_2 = 32'h0;
    if(execute_CsrPlugin_csr_1968) begin
      _zz_CsrPlugin_csrMapping_readDataInit_2[3 : 3] = CsrPlugin_dcsr_nmip;
      _zz_CsrPlugin_csrMapping_readDataInit_2[8 : 6] = CsrPlugin_dcsr_cause;
      _zz_CsrPlugin_csrMapping_readDataInit_2[31 : 28] = CsrPlugin_dcsr_xdebugver;
      _zz_CsrPlugin_csrMapping_readDataInit_2[4 : 4] = CsrPlugin_dcsr_mprven;
      _zz_CsrPlugin_csrMapping_readDataInit_2[1 : 0] = CsrPlugin_dcsr_prv;
      _zz_CsrPlugin_csrMapping_readDataInit_2[2 : 2] = CsrPlugin_dcsr_step;
      _zz_CsrPlugin_csrMapping_readDataInit_2[9 : 9] = CsrPlugin_dcsr_stoptime;
      _zz_CsrPlugin_csrMapping_readDataInit_2[10 : 10] = CsrPlugin_dcsr_stopcount;
      _zz_CsrPlugin_csrMapping_readDataInit_2[11 : 11] = CsrPlugin_dcsr_stepie;
      _zz_CsrPlugin_csrMapping_readDataInit_2[15 : 15] = CsrPlugin_dcsr_ebreakm;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_3 = 32'h0;
    if(execute_CsrPlugin_csr_3860) begin
      _zz_CsrPlugin_csrMapping_readDataInit_3[0 : 0] = 1'b1;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_4 = 32'h0;
    if(execute_CsrPlugin_csr_769) begin
      _zz_CsrPlugin_csrMapping_readDataInit_4[31 : 30] = CsrPlugin_misa_base;
      _zz_CsrPlugin_csrMapping_readDataInit_4[25 : 0] = CsrPlugin_misa_extensions;
    end
  end

  assign switch_CsrPlugin_l1167 = CsrPlugin_csrMapping_writeDataSignal[12 : 11];
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_5 = 32'h0;
    if(execute_CsrPlugin_csr_768) begin
      _zz_CsrPlugin_csrMapping_readDataInit_5[7 : 7] = CsrPlugin_mstatus_MPIE;
      _zz_CsrPlugin_csrMapping_readDataInit_5[3 : 3] = CsrPlugin_mstatus_MIE;
      _zz_CsrPlugin_csrMapping_readDataInit_5[12 : 11] = CsrPlugin_mstatus_MPP;
      _zz_CsrPlugin_csrMapping_readDataInit_5[14 : 13] = FpuPlugin_fs;
      _zz_CsrPlugin_csrMapping_readDataInit_5[31 : 31] = FpuPlugin_sd;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_6 = 32'h0;
    if(execute_CsrPlugin_csr_836) begin
      _zz_CsrPlugin_csrMapping_readDataInit_6[11 : 11] = CsrPlugin_mip_MEIP;
      _zz_CsrPlugin_csrMapping_readDataInit_6[7 : 7] = CsrPlugin_mip_MTIP;
      _zz_CsrPlugin_csrMapping_readDataInit_6[3 : 3] = CsrPlugin_mip_MSIP;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_7 = 32'h0;
    if(execute_CsrPlugin_csr_772) begin
      _zz_CsrPlugin_csrMapping_readDataInit_7[11 : 11] = CsrPlugin_mie_MEIE;
      _zz_CsrPlugin_csrMapping_readDataInit_7[7 : 7] = CsrPlugin_mie_MTIE;
      _zz_CsrPlugin_csrMapping_readDataInit_7[3 : 3] = CsrPlugin_mie_MSIE;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_8 = 32'h0;
    if(execute_CsrPlugin_csr_773) begin
      _zz_CsrPlugin_csrMapping_readDataInit_8[31 : 2] = CsrPlugin_mtvec_base;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_9 = 32'h0;
    if(execute_CsrPlugin_csr_833) begin
      _zz_CsrPlugin_csrMapping_readDataInit_9[31 : 0] = CsrPlugin_mepc;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_10 = 32'h0;
    if(execute_CsrPlugin_csr_832) begin
      _zz_CsrPlugin_csrMapping_readDataInit_10[31 : 0] = CsrPlugin_mscratch;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_11 = 32'h0;
    if(execute_CsrPlugin_csr_834) begin
      _zz_CsrPlugin_csrMapping_readDataInit_11[31 : 31] = CsrPlugin_mcause_interrupt;
      _zz_CsrPlugin_csrMapping_readDataInit_11[3 : 0] = CsrPlugin_mcause_exceptionCode;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_12 = 32'h0;
    if(execute_CsrPlugin_csr_835) begin
      _zz_CsrPlugin_csrMapping_readDataInit_12[31 : 0] = CsrPlugin_mtval;
    end
  end

  assign _zz_FpuPlugin_flags_NX = CsrPlugin_csrMapping_writeDataSignal[4 : 0];
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_13 = 32'h0;
    if(execute_CsrPlugin_csr_3) begin
      _zz_CsrPlugin_csrMapping_readDataInit_13[7 : 5] = FpuPlugin_rm;
      _zz_CsrPlugin_csrMapping_readDataInit_13[4 : 0] = {FpuPlugin_flags_NV,{FpuPlugin_flags_DZ,{FpuPlugin_flags_OF,{FpuPlugin_flags_UF,FpuPlugin_flags_NX}}}};
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_14 = 32'h0;
    if(execute_CsrPlugin_csr_2) begin
      _zz_CsrPlugin_csrMapping_readDataInit_14[2 : 0] = FpuPlugin_rm;
    end
  end

  assign _zz_FpuPlugin_flags_NX_1 = CsrPlugin_csrMapping_writeDataSignal[4 : 0];
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_15 = 32'h0;
    if(execute_CsrPlugin_csr_1) begin
      _zz_CsrPlugin_csrMapping_readDataInit_15[4 : 0] = {FpuPlugin_flags_NV,{FpuPlugin_flags_DZ,{FpuPlugin_flags_OF,{FpuPlugin_flags_UF,FpuPlugin_flags_NX}}}};
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_16 = 32'h0;
    if(execute_CsrPlugin_csr_256) begin
      _zz_CsrPlugin_csrMapping_readDataInit_16[14 : 13] = FpuPlugin_fs;
      _zz_CsrPlugin_csrMapping_readDataInit_16[31 : 31] = FpuPlugin_sd;
    end
  end

  assign CsrPlugin_csrMapping_readDataInit = (((((_zz_CsrPlugin_csrMapping_readDataInit | _zz_CsrPlugin_csrMapping_readDataInit_1) | (_zz_CsrPlugin_csrMapping_readDataInit_2 | _zz_CsrPlugin_csrMapping_readDataInit_17)) | ((_zz_CsrPlugin_csrMapping_readDataInit_18 | _zz_CsrPlugin_csrMapping_readDataInit_19) | (_zz_CsrPlugin_csrMapping_readDataInit_3 | _zz_CsrPlugin_csrMapping_readDataInit_4))) | (((_zz_CsrPlugin_csrMapping_readDataInit_5 | _zz_CsrPlugin_csrMapping_readDataInit_6) | (_zz_CsrPlugin_csrMapping_readDataInit_7 | _zz_CsrPlugin_csrMapping_readDataInit_8)) | ((_zz_CsrPlugin_csrMapping_readDataInit_9 | _zz_CsrPlugin_csrMapping_readDataInit_10) | (_zz_CsrPlugin_csrMapping_readDataInit_11 | _zz_CsrPlugin_csrMapping_readDataInit_12)))) | ((_zz_CsrPlugin_csrMapping_readDataInit_13 | _zz_CsrPlugin_csrMapping_readDataInit_14) | (_zz_CsrPlugin_csrMapping_readDataInit_15 | _zz_CsrPlugin_csrMapping_readDataInit_16)));
  assign when_CsrPlugin_l1846 = ((execute_arbitration_isValid && execute_IS_CSR) && (({execute_CsrPlugin_csrAddress[11 : 2],2'b00} == 12'h3a0) || ({execute_CsrPlugin_csrAddress[11 : 4],4'b0000} == 12'h3b0)));
  assign _zz_when_CsrPlugin_l1853 = (execute_CsrPlugin_csrAddress & 12'hf60);
  assign when_CsrPlugin_l1853 = (((execute_arbitration_isValid && execute_IS_CSR) && (5'h03 <= execute_CsrPlugin_csrAddress[4 : 0])) && (((_zz_when_CsrPlugin_l1853 == 12'hb00) || (((_zz_when_CsrPlugin_l1853 == 12'hc00) && (! execute_CsrPlugin_writeInstruction)) && (CsrPlugin_privilege == 2'b11))) || ((execute_CsrPlugin_csrAddress & 12'hfe0) == 12'h320)));
  always @(*) begin
    when_CsrPlugin_l1863 = CsrPlugin_csrMapping_doForceFailCsr;
    if(when_CsrPlugin_l1861) begin
      when_CsrPlugin_l1863 = 1'b1;
    end
    if(when_CsrPlugin_l1862) begin
      when_CsrPlugin_l1863 = 1'b1;
    end
  end

  assign when_CsrPlugin_l1861 = (CsrPlugin_privilege < execute_CsrPlugin_csrAddress[9 : 8]);
  assign when_CsrPlugin_l1862 = ((! debugMode) && (_zz_when_CsrPlugin_l1862 == 8'h7b));
  assign when_CsrPlugin_l1869 = ((! execute_arbitration_isValid) || (! execute_IS_CSR));
  always @(*) begin
    FpuPlugin_stateNext = FpuPlugin_stateReg;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
        if(fpuAccess_start) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_CMD;
        end
      end
      FpuPlugin_enumDef_CMD : begin
        if(fpuAccess_write) begin
          if(FpuPlugin_port_cmd_ready) begin
            FpuPlugin_stateNext = FpuPlugin_enumDef_COMMIT;
          end
        end else begin
          if(FpuPlugin_port_cmd_ready) begin
            FpuPlugin_stateNext = FpuPlugin_enumDef_RSP;
          end
        end
      end
      FpuPlugin_enumDef_RSP : begin
        if(FpuPlugin_port_rsp_valid) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_RSP_0;
        end
      end
      FpuPlugin_enumDef_RSP_0 : begin
        if(when_FpuPlugin_l402) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_RSP_1;
        end else begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_DONE;
        end
      end
      FpuPlugin_enumDef_RSP_1 : begin
        FpuPlugin_stateNext = FpuPlugin_enumDef_DONE;
      end
      FpuPlugin_enumDef_COMMIT : begin
        if(FpuPlugin_port_commit_ready) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_DONE;
        end
      end
      FpuPlugin_enumDef_DONE : begin
        FpuPlugin_stateNext = FpuPlugin_enumDef_IDLE;
      end
      default : begin
      end
    endcase
    if(FpuPlugin_wantStart) begin
      FpuPlugin_stateNext = FpuPlugin_enumDef_IDLE;
    end
    if(FpuPlugin_wantKill) begin
      FpuPlugin_stateNext = FpuPlugin_enumDef_BOOT;
    end
  end

  always @(*) begin
    _zz_FpuPlugin_port_cmd_payload_format = (1'bx);
    case(fpuAccess_size)
      3'b010 : begin
        _zz_FpuPlugin_port_cmd_payload_format = FpuFormat_FLOAT;
      end
      3'b011 : begin
        _zz_FpuPlugin_port_cmd_payload_format = FpuFormat_DOUBLE;
      end
      default : begin
      end
    endcase
  end

  assign when_FpuPlugin_l402 = (3'b010 < fpuAccess_size);
  assign DBusCachedPlugin_trigger_hitBefore = 1'b0;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      IBusCachedPlugin_fetchPc_pcReg <= 32'hf9000000;
      IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      IBusCachedPlugin_fetchPc_booted <= 1'b0;
      IBusCachedPlugin_fetchPc_inc <= 1'b0;
      IBusCachedPlugin_decodePc_pcReg <= 32'hf9000000;
      _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1 <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      IBusCachedPlugin_decompressor_bufferValid <= 1'b0;
      IBusCachedPlugin_decompressor_throw2BytesReg <= 1'b0;
      _zz_IBusCachedPlugin_injector_decodeInput_valid <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      IBusCachedPlugin_rspCounter <= 32'h0;
      dataCache_2_io_mem_cmd_rValidN <= 1'b1;
      dataCache_2_io_mem_cmd_s2mPipe_rValid <= 1'b0;
      dBus_rsp_valid_regNext <= 1'b0;
      DBusCachedPlugin_rspCounter <= 32'h0;
      _zz_5 <= 1'b1;
      HazardSimplePlugin_writeBackBuffer_valid <= 1'b0;
      _zz_CsrPlugin_privilege <= 2'b11;
      CsrPlugin_running <= 1'b1;
      CsrPlugin_reseting <= 1'b1;
      _zz_debugBus_haveReset <= 1'b0;
      CsrPlugin_running_aheadValue_regNext <= 1'b0;
      CsrPlugin_doHalt <= 1'b0;
      _zz_CsrPlugin_doResume <= 1'b0;
      CsrPlugin_timeout_state <= 1'b0;
      CsrPlugin_timeout_counter_value <= 3'b000;
      CsrPlugin_inject_cmd_toStream_rValid <= 1'b0;
      CsrPlugin_inject_pending <= 1'b0;
      CsrPlugin_dcsr_prv <= 2'b11;
      CsrPlugin_dcsr_step <= 1'b0;
      CsrPlugin_dcsr_cause <= 3'b000;
      CsrPlugin_dcsr_stoptime <= 1'b1;
      CsrPlugin_dcsr_stopcount <= 1'b0;
      CsrPlugin_dcsr_stepie <= 1'b0;
      CsrPlugin_dcsr_ebreakm <= 1'b0;
      CsrPlugin_dcsr_stepLogic_stateReg <= CsrPlugin_dcsr_stepLogic_enumDef_BOOT;
      stoptime <= 1'b0;
      CsrPlugin_mstatus_MIE <= 1'b0;
      CsrPlugin_mstatus_MPIE <= 1'b0;
      CsrPlugin_mstatus_MPP <= 2'b11;
      CsrPlugin_mie_MEIE <= 1'b0;
      CsrPlugin_mie_MTIE <= 1'b0;
      CsrPlugin_mie_MSIE <= 1'b0;
      CsrPlugin_counters_mcycle <= 64'h0;
      CsrPlugin_counters_minstret <= 64'h0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      CsrPlugin_interrupt_valid <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      CsrPlugin_hadException <= 1'b0;
      execute_CsrPlugin_wfiWake <= 1'b0;
      memory_MulDivIterativePlugin_div_counter_value <= 6'h0;
      FpuPlugin_pendings <= 6'h0;
      FpuPlugin_flags_NV <= 1'b0;
      FpuPlugin_flags_DZ <= 1'b0;
      FpuPlugin_flags_OF <= 1'b0;
      FpuPlugin_flags_UF <= 1'b0;
      FpuPlugin_flags_NX <= 1'b0;
      FpuPlugin_rm <= 3'b000;
      FpuPlugin_fs <= 2'b01;
      decode_FpuPlugin_forked <= 1'b0;
      writeBack_FpuPlugin_commit_rValidN <= 1'b1;
      execute_CfuPlugin_hold <= 1'b0;
      execute_CfuPlugin_fired <= 1'b0;
      CfuPlugin_bus_rsp_rValidN <= 1'b1;
      execute_arbitration_isValid <= 1'b0;
      memory_arbitration_isValid <= 1'b0;
      writeBack_arbitration_isValid <= 1'b0;
      IBusCachedPlugin_injector_port_state <= 3'b000;
      FpuPlugin_stateReg <= FpuPlugin_enumDef_BOOT;
      decode_to_execute_FPU_FORKED <= 1'b0;
      execute_to_memory_FPU_FORKED <= 1'b0;
      memory_to_writeBack_FPU_FORKED <= 1'b0;
      memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT <= 1'b0;
      execute_to_memory_CfuPlugin_CFU_IN_FLIGHT <= 1'b0;
    end else begin
      if(IBusCachedPlugin_fetchPc_correction) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_output_fire) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      end
      IBusCachedPlugin_fetchPc_booted <= 1'b1;
      if(when_Fetcher_l133) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_output_fire) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b1;
      end
      if(when_Fetcher_l133_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(when_Fetcher_l160) begin
        IBusCachedPlugin_fetchPc_pcReg <= IBusCachedPlugin_fetchPc_pc;
      end
      if(when_Fetcher_l182) begin
        IBusCachedPlugin_decodePc_pcReg <= IBusCachedPlugin_decodePc_pcPlus;
      end
      if(when_Fetcher_l194) begin
        IBusCachedPlugin_decodePc_pcReg <= IBusCachedPlugin_jump_pcLoad_payload;
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1 <= 1'b0;
      end
      if(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1 <= (IBusCachedPlugin_iBusRsp_stages_0_output_valid && (! 1'b0));
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      end
      if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= (IBusCachedPlugin_iBusRsp_stages_1_output_valid && (! IBusCachedPlugin_iBusRsp_flush));
      end
      if(IBusCachedPlugin_decompressor_output_fire) begin
        IBusCachedPlugin_decompressor_throw2BytesReg <= ((((! IBusCachedPlugin_decompressor_unaligned) && IBusCachedPlugin_decompressor_isInputLowRvc) && IBusCachedPlugin_decompressor_isInputHighRvc) || (IBusCachedPlugin_decompressor_bufferValid && IBusCachedPlugin_decompressor_isInputHighRvc));
      end
      if(when_Fetcher_l285) begin
        IBusCachedPlugin_decompressor_bufferValid <= 1'b0;
      end
      if(when_Fetcher_l288) begin
        if(IBusCachedPlugin_decompressor_bufferFill) begin
          IBusCachedPlugin_decompressor_bufferValid <= 1'b1;
        end
      end
      if(when_Fetcher_l293) begin
        IBusCachedPlugin_decompressor_throw2BytesReg <= 1'b0;
        IBusCachedPlugin_decompressor_bufferValid <= 1'b0;
      end
      if(decode_arbitration_removeIt) begin
        _zz_IBusCachedPlugin_injector_decodeInput_valid <= 1'b0;
      end
      if(IBusCachedPlugin_decompressor_output_ready) begin
        _zz_IBusCachedPlugin_injector_decodeInput_valid <= (IBusCachedPlugin_decompressor_output_valid && (! IBusCachedPlugin_externalFlush));
      end
      if(when_Fetcher_l331) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b1;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      end
      if(when_Fetcher_l331_1) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= IBusCachedPlugin_injector_nextPcCalc_valids_0;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(when_Fetcher_l331_2) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= IBusCachedPlugin_injector_nextPcCalc_valids_1;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(when_Fetcher_l331_3) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= IBusCachedPlugin_injector_nextPcCalc_valids_2;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(iBus_rsp_valid) begin
        IBusCachedPlugin_rspCounter <= (IBusCachedPlugin_rspCounter + 32'h00000001);
      end
      if(dataCache_2_io_mem_cmd_valid) begin
        dataCache_2_io_mem_cmd_rValidN <= 1'b0;
      end
      if(dataCache_2_io_mem_cmd_s2mPipe_ready) begin
        dataCache_2_io_mem_cmd_rValidN <= 1'b1;
      end
      if(dataCache_2_io_mem_cmd_s2mPipe_ready) begin
        dataCache_2_io_mem_cmd_s2mPipe_rValid <= dataCache_2_io_mem_cmd_s2mPipe_valid;
      end
      dBus_rsp_valid_regNext <= dBus_rsp_valid;
      if(dBus_rsp_valid) begin
        DBusCachedPlugin_rspCounter <= (DBusCachedPlugin_rspCounter + 32'h00000001);
      end
      _zz_5 <= 1'b0;
      HazardSimplePlugin_writeBackBuffer_valid <= HazardSimplePlugin_writeBackWrites_valid;
      CsrPlugin_reseting <= 1'b0;
      if(CsrPlugin_reseting) begin
        _zz_debugBus_haveReset <= 1'b1;
      end
      if(debugBus_ackReset) begin
        _zz_debugBus_haveReset <= 1'b0;
      end
      CsrPlugin_running_aheadValue_regNext <= CsrPlugin_running_aheadValue;
      if(when_CsrPlugin_l747) begin
        CsrPlugin_doHalt <= 1'b1;
      end
      if(CsrPlugin_enterHalt) begin
        CsrPlugin_doHalt <= 1'b0;
      end
      if(debugBus_resume_cmd_valid) begin
        _zz_CsrPlugin_doResume <= 1'b1;
      end
      if(debugBus_resume_rsp_valid) begin
        _zz_CsrPlugin_doResume <= 1'b0;
      end
      CsrPlugin_timeout_counter_value <= CsrPlugin_timeout_counter_valueNext;
      if(CsrPlugin_timeout_counter_willOverflow) begin
        CsrPlugin_timeout_state <= 1'b1;
      end
      if(when_CsrPlugin_l753) begin
        CsrPlugin_timeout_state <= 1'b0;
      end
      if(CsrPlugin_inject_cmd_toStream_ready) begin
        CsrPlugin_inject_cmd_toStream_rValid <= CsrPlugin_inject_cmd_toStream_valid;
      end
      if(when_CsrPlugin_l804) begin
        CsrPlugin_inject_pending <= 1'b1;
      end
      if(when_CsrPlugin_l804_1) begin
        CsrPlugin_inject_pending <= 1'b0;
      end
      if(CsrPlugin_inject_cmd_valid) begin
        CsrPlugin_timeout_state <= 1'b0;
      end
      CsrPlugin_dcsr_stepLogic_stateReg <= CsrPlugin_dcsr_stepLogic_stateNext;
      case(CsrPlugin_dcsr_stepLogic_stateReg)
        CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
        end
        CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
          CsrPlugin_timeout_state <= 1'b0;
          if(when_CsrPlugin_l836) begin
            CsrPlugin_doHalt <= 1'b1;
          end
        end
        CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
          if(!when_CsrPlugin_l848) begin
            if(writeBack_arbitration_isFiring) begin
              CsrPlugin_doHalt <= 1'b1;
            end
          end
        end
        default : begin
        end
      endcase
      stoptime <= (debugMode && CsrPlugin_dcsr_stoptime);
      CsrPlugin_counters_mcycle <= (CsrPlugin_counters_mcycle + _zz_CsrPlugin_counters_mcycle);
      if(writeBack_arbitration_isFiring) begin
        CsrPlugin_counters_minstret <= (CsrPlugin_counters_minstret + _zz_CsrPlugin_counters_minstret);
      end
      if(when_CsrPlugin_l1403) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
      end
      if(when_CsrPlugin_l1403_1) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= (CsrPlugin_exceptionPortCtrl_exceptionValids_decode && (! decode_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
      end
      if(when_CsrPlugin_l1403_2) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= (CsrPlugin_exceptionPortCtrl_exceptionValids_execute && (! execute_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
      end
      if(when_CsrPlugin_l1403_3) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= (CsrPlugin_exceptionPortCtrl_exceptionValids_memory && (! memory_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      end
      CsrPlugin_interrupt_valid <= 1'b0;
      if(when_CsrPlugin_l1440) begin
        if(when_CsrPlugin_l1446) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l1446_1) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l1446_2) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
      end
      if(when_CsrPlugin_l1459) begin
        CsrPlugin_interrupt_valid <= 1'b0;
      end
      if(CsrPlugin_doHalt) begin
        CsrPlugin_interrupt_valid <= 1'b1;
      end
      if(CsrPlugin_pipelineLiberator_active) begin
        if(when_CsrPlugin_l1479) begin
          CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b1;
        end
        if(when_CsrPlugin_l1479_1) begin
          CsrPlugin_pipelineLiberator_pcValids_1 <= CsrPlugin_pipelineLiberator_pcValids_0;
        end
        if(when_CsrPlugin_l1479_2) begin
          CsrPlugin_pipelineLiberator_pcValids_2 <= CsrPlugin_pipelineLiberator_pcValids_1;
        end
      end
      if(when_CsrPlugin_l1484) begin
        CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      end
      if(CsrPlugin_interruptJump) begin
        CsrPlugin_interrupt_valid <= 1'b0;
      end
      CsrPlugin_hadException <= CsrPlugin_exception;
      if(when_CsrPlugin_l1534) begin
        if(when_CsrPlugin_l1542) begin
          _zz_CsrPlugin_privilege <= CsrPlugin_targetPrivilege;
          case(CsrPlugin_targetPrivilege)
            2'b11 : begin
              CsrPlugin_mstatus_MIE <= 1'b0;
              CsrPlugin_mstatus_MPIE <= CsrPlugin_mstatus_MIE;
              CsrPlugin_mstatus_MPP <= CsrPlugin_privilege;
            end
            default : begin
            end
          endcase
        end else begin
          if(when_CsrPlugin_l1572) begin
            CsrPlugin_dcsr_cause <= 3'b011;
            if(CsrPlugin_dcsr_step) begin
              CsrPlugin_dcsr_cause <= 3'b100;
            end
            if(CsrPlugin_trapCauseEbreakDebug) begin
              CsrPlugin_dcsr_cause <= 3'b001;
            end
            CsrPlugin_dcsr_prv <= CsrPlugin_privilege;
          end
          _zz_CsrPlugin_privilege <= 2'b11;
        end
      end
      if(when_CsrPlugin_l1600) begin
        case(switch_CsrPlugin_l1604)
          2'b11 : begin
            CsrPlugin_mstatus_MPP <= 2'b00;
            CsrPlugin_mstatus_MIE <= CsrPlugin_mstatus_MPIE;
            CsrPlugin_mstatus_MPIE <= 1'b1;
            _zz_CsrPlugin_privilege <= CsrPlugin_mstatus_MPP;
          end
          default : begin
          end
        endcase
      end
      if(CsrPlugin_doResume) begin
        _zz_CsrPlugin_privilege <= CsrPlugin_dcsr_prv;
      end
      execute_CsrPlugin_wfiWake <= ((|{_zz_when_CsrPlugin_l1446_2,{_zz_when_CsrPlugin_l1446_1,_zz_when_CsrPlugin_l1446}}) || CsrPlugin_thirdPartyWake);
      memory_MulDivIterativePlugin_div_counter_value <= memory_MulDivIterativePlugin_div_counter_valueNext;
      FpuPlugin_pendings <= (_zz_FpuPlugin_pendings - _zz_FpuPlugin_pendings_6);
      if(when_FpuPlugin_l215) begin
        FpuPlugin_flags_NV <= 1'b1;
      end
      if(when_FpuPlugin_l216) begin
        FpuPlugin_flags_DZ <= 1'b1;
      end
      if(when_FpuPlugin_l217) begin
        FpuPlugin_flags_OF <= 1'b1;
      end
      if(when_FpuPlugin_l218) begin
        FpuPlugin_flags_UF <= 1'b1;
      end
      if(when_FpuPlugin_l219) begin
        FpuPlugin_flags_NX <= 1'b1;
      end
      if(when_FpuPlugin_l234) begin
        FpuPlugin_fs <= 2'b11;
      end
      if(when_FpuPlugin_l237) begin
        FpuPlugin_fs <= 2'b11;
      end
      if(when_FpuPlugin_l268) begin
        decode_FpuPlugin_forked <= 1'b1;
      end
      if(when_FpuPlugin_l268_1) begin
        decode_FpuPlugin_forked <= 1'b0;
      end
      if(writeBack_FpuPlugin_isRsp) begin
        if(writeBack_arbitration_isValid) begin
          if(when_FpuPlugin_l315) begin
            if(FpuPlugin_port_rsp_payload_NV) begin
              FpuPlugin_flags_NV <= 1'b1;
            end
            if(FpuPlugin_port_rsp_payload_NX) begin
              FpuPlugin_flags_NX <= 1'b1;
            end
            if(when_FpuPlugin_l318) begin
              FpuPlugin_fs <= 2'b11;
            end
          end
        end
      end
      if(writeBack_FpuPlugin_commit_valid) begin
        writeBack_FpuPlugin_commit_rValidN <= 1'b0;
      end
      if(writeBack_FpuPlugin_commit_s2mPipe_ready) begin
        writeBack_FpuPlugin_commit_rValidN <= 1'b1;
      end
      if(execute_CfuPlugin_schedule) begin
        execute_CfuPlugin_hold <= 1'b1;
      end
      if(CfuPlugin_bus_cmd_ready) begin
        execute_CfuPlugin_hold <= 1'b0;
      end
      if(CfuPlugin_bus_cmd_fire) begin
        execute_CfuPlugin_fired <= 1'b1;
      end
      if(when_CfuPlugin_l199) begin
        execute_CfuPlugin_fired <= 1'b0;
      end
      if(CfuPlugin_bus_rsp_valid) begin
        CfuPlugin_bus_rsp_rValidN <= 1'b0;
      end
      if(writeBack_CfuPlugin_rsp_ready) begin
        CfuPlugin_bus_rsp_rValidN <= 1'b1;
      end
      if(when_Pipeline_l124_75) begin
        decode_to_execute_FPU_FORKED <= _zz_decode_to_execute_FPU_FORKED;
      end
      if(when_Pipeline_l124_76) begin
        execute_to_memory_FPU_FORKED <= _zz_execute_to_memory_FPU_FORKED;
      end
      if(when_Pipeline_l124_77) begin
        memory_to_writeBack_FPU_FORKED <= _zz_memory_to_writeBack_FPU_FORKED;
      end
      if(when_Pipeline_l124_91) begin
        execute_to_memory_CfuPlugin_CFU_IN_FLIGHT <= _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
      end
      if(when_Pipeline_l124_92) begin
        memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT <= _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
      end
      if(when_Pipeline_l151) begin
        execute_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154) begin
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end
      if(when_Pipeline_l151_1) begin
        memory_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_1) begin
        memory_arbitration_isValid <= execute_arbitration_isValid;
      end
      if(when_Pipeline_l151_2) begin
        writeBack_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_2) begin
        writeBack_arbitration_isValid <= memory_arbitration_isValid;
      end
      case(IBusCachedPlugin_injector_port_state)
        3'b000 : begin
          if(CsrPlugin_injectionPort_valid) begin
            IBusCachedPlugin_injector_port_state <= 3'b001;
          end
        end
        3'b001 : begin
          IBusCachedPlugin_injector_port_state <= 3'b010;
        end
        3'b010 : begin
          IBusCachedPlugin_injector_port_state <= 3'b011;
        end
        3'b011 : begin
          if(when_Fetcher_l391) begin
            IBusCachedPlugin_injector_port_state <= 3'b100;
          end
        end
        3'b100 : begin
          IBusCachedPlugin_injector_port_state <= 3'b000;
        end
        default : begin
        end
      endcase
      if(execute_CsrPlugin_csr_1968) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_dcsr_prv <= CsrPlugin_csrMapping_writeDataSignal[1 : 0];
          CsrPlugin_dcsr_step <= CsrPlugin_csrMapping_writeDataSignal[2];
          CsrPlugin_dcsr_stoptime <= CsrPlugin_csrMapping_writeDataSignal[9];
          CsrPlugin_dcsr_stopcount <= CsrPlugin_csrMapping_writeDataSignal[10];
          CsrPlugin_dcsr_stepie <= CsrPlugin_csrMapping_writeDataSignal[11];
          CsrPlugin_dcsr_ebreakm <= CsrPlugin_csrMapping_writeDataSignal[15];
        end
      end
      if(execute_CsrPlugin_csr_768) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mstatus_MPIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mstatus_MIE <= CsrPlugin_csrMapping_writeDataSignal[3];
          case(switch_CsrPlugin_l1167)
            2'b11 : begin
              CsrPlugin_mstatus_MPP <= 2'b11;
            end
            default : begin
            end
          endcase
          FpuPlugin_fs <= CsrPlugin_csrMapping_writeDataSignal[14 : 13];
        end
      end
      if(execute_CsrPlugin_csr_772) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mie_MEIE <= CsrPlugin_csrMapping_writeDataSignal[11];
          CsrPlugin_mie_MTIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mie_MSIE <= CsrPlugin_csrMapping_writeDataSignal[3];
        end
      end
      if(execute_CsrPlugin_csr_3) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_rm <= CsrPlugin_csrMapping_writeDataSignal[7 : 5];
          FpuPlugin_flags_NX <= _zz_FpuPlugin_flags_NX[0];
          FpuPlugin_flags_UF <= _zz_FpuPlugin_flags_NX[1];
          FpuPlugin_flags_OF <= _zz_FpuPlugin_flags_NX[2];
          FpuPlugin_flags_DZ <= _zz_FpuPlugin_flags_NX[3];
          FpuPlugin_flags_NV <= _zz_FpuPlugin_flags_NX[4];
        end
      end
      if(execute_CsrPlugin_csr_2) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_rm <= CsrPlugin_csrMapping_writeDataSignal[2 : 0];
        end
      end
      if(execute_CsrPlugin_csr_1) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_flags_NX <= _zz_FpuPlugin_flags_NX_1[0];
          FpuPlugin_flags_UF <= _zz_FpuPlugin_flags_NX_1[1];
          FpuPlugin_flags_OF <= _zz_FpuPlugin_flags_NX_1[2];
          FpuPlugin_flags_DZ <= _zz_FpuPlugin_flags_NX_1[3];
          FpuPlugin_flags_NV <= _zz_FpuPlugin_flags_NX_1[4];
        end
      end
      if(execute_CsrPlugin_csr_256) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_fs <= CsrPlugin_csrMapping_writeDataSignal[14 : 13];
        end
      end
      FpuPlugin_stateReg <= FpuPlugin_stateNext;
      CsrPlugin_running <= CsrPlugin_running_aheadValue;
    end
  end

  always @(posedge io_systemClk) begin
    if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload <= IBusCachedPlugin_iBusRsp_stages_1_output_payload;
    end
    if(IBusCachedPlugin_decompressor_input_valid) begin
      IBusCachedPlugin_decompressor_bufferValidLatch <= IBusCachedPlugin_decompressor_bufferValid;
    end
    if(IBusCachedPlugin_decompressor_input_valid) begin
      IBusCachedPlugin_decompressor_throw2BytesLatch <= IBusCachedPlugin_decompressor_throw2Bytes;
    end
    if(when_Fetcher_l288) begin
      IBusCachedPlugin_decompressor_bufferData <= IBusCachedPlugin_decompressor_input_payload_rsp_inst[31 : 16];
    end
    if(IBusCachedPlugin_decompressor_output_ready) begin
      _zz_IBusCachedPlugin_injector_decodeInput_payload_pc <= IBusCachedPlugin_decompressor_output_payload_pc;
      _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_error <= IBusCachedPlugin_decompressor_output_payload_rsp_error;
      _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst <= IBusCachedPlugin_decompressor_output_payload_rsp_inst;
      _zz_IBusCachedPlugin_injector_decodeInput_payload_isRvc <= IBusCachedPlugin_decompressor_output_payload_isRvc;
    end
    if(IBusCachedPlugin_injector_decodeInput_ready) begin
      IBusCachedPlugin_injector_formal_rawInDecode <= IBusCachedPlugin_decompressor_raw;
    end
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_s1_tightlyCoupledHit <= IBusCachedPlugin_s0_tightlyCoupledHit;
    end
    if(IBusCachedPlugin_iBusRsp_stages_2_input_ready) begin
      IBusCachedPlugin_s2_tightlyCoupledHit <= IBusCachedPlugin_s1_tightlyCoupledHit;
    end
    if(dataCache_2_io_mem_cmd_rValidN) begin
      dataCache_2_io_mem_cmd_rData_wr <= dataCache_2_io_mem_cmd_payload_wr;
      dataCache_2_io_mem_cmd_rData_uncached <= dataCache_2_io_mem_cmd_payload_uncached;
      dataCache_2_io_mem_cmd_rData_address <= dataCache_2_io_mem_cmd_payload_address;
      dataCache_2_io_mem_cmd_rData_data <= dataCache_2_io_mem_cmd_payload_data;
      dataCache_2_io_mem_cmd_rData_mask <= dataCache_2_io_mem_cmd_payload_mask;
      dataCache_2_io_mem_cmd_rData_size <= dataCache_2_io_mem_cmd_payload_size;
      dataCache_2_io_mem_cmd_rData_exclusive <= dataCache_2_io_mem_cmd_payload_exclusive;
      dataCache_2_io_mem_cmd_rData_last <= dataCache_2_io_mem_cmd_payload_last;
    end
    if(dataCache_2_io_mem_cmd_s2mPipe_ready) begin
      dataCache_2_io_mem_cmd_s2mPipe_rData_wr <= dataCache_2_io_mem_cmd_s2mPipe_payload_wr;
      dataCache_2_io_mem_cmd_s2mPipe_rData_uncached <= dataCache_2_io_mem_cmd_s2mPipe_payload_uncached;
      dataCache_2_io_mem_cmd_s2mPipe_rData_address <= dataCache_2_io_mem_cmd_s2mPipe_payload_address;
      dataCache_2_io_mem_cmd_s2mPipe_rData_data <= dataCache_2_io_mem_cmd_s2mPipe_payload_data;
      dataCache_2_io_mem_cmd_s2mPipe_rData_mask <= dataCache_2_io_mem_cmd_s2mPipe_payload_mask;
      dataCache_2_io_mem_cmd_s2mPipe_rData_size <= dataCache_2_io_mem_cmd_s2mPipe_payload_size;
      dataCache_2_io_mem_cmd_s2mPipe_rData_exclusive <= dataCache_2_io_mem_cmd_s2mPipe_payload_exclusive;
      dataCache_2_io_mem_cmd_s2mPipe_rData_last <= dataCache_2_io_mem_cmd_s2mPipe_payload_last;
    end
    dBus_rsp_payload_exclusive_regNext <= dBus_rsp_payload_exclusive;
    dBus_rsp_payload_error_regNext <= dBus_rsp_payload_error;
    dBus_rsp_payload_last_regNext <= dBus_rsp_payload_last;
    dBus_rsp_payload_aggregated_regNext <= dBus_rsp_payload_aggregated;
    if(when_DBusCachedPlugin_l334) begin
      dBus_rsp_payload_data_regNextWhen <= dBus_rsp_payload_data;
    end
    HazardSimplePlugin_writeBackBuffer_payload_address <= HazardSimplePlugin_writeBackWrites_payload_address;
    HazardSimplePlugin_writeBackBuffer_payload_data <= HazardSimplePlugin_writeBackWrites_payload_data;
    if(when_CsrPlugin_l768) begin
      if(_zz_6[0]) begin
        CsrPlugin_dataCsrw_value_0 <= debugBus_dmToHart_payload_data;
      end
      if(_zz_6[1]) begin
        CsrPlugin_dataCsrw_value_1 <= debugBus_dmToHart_payload_data;
      end
    end
    if(CsrPlugin_inject_cmd_toStream_ready) begin
      CsrPlugin_inject_cmd_toStream_rData_op <= CsrPlugin_inject_cmd_toStream_payload_op;
      CsrPlugin_inject_cmd_toStream_rData_address <= CsrPlugin_inject_cmd_toStream_payload_address;
      CsrPlugin_inject_cmd_toStream_rData_data <= CsrPlugin_inject_cmd_toStream_payload_data;
      CsrPlugin_inject_cmd_toStream_rData_size <= CsrPlugin_inject_cmd_toStream_payload_size;
    end
    CsrPlugin_mip_MEIP <= externalInterrupt;
    CsrPlugin_mip_MTIP <= timerInterrupt;
    CsrPlugin_mip_MSIP <= softwareInterrupt;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_code : decodeExceptionPort_payload_code);
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_badAddr : decodeExceptionPort_payload_badAddr);
    end
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= CsrPlugin_selfException_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= CsrPlugin_selfException_payload_badAddr;
    end
    if(DBusCachedPlugin_exceptionBus_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= DBusCachedPlugin_exceptionBus_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= DBusCachedPlugin_exceptionBus_payload_badAddr;
    end
    if(when_CsrPlugin_l1440) begin
      if(when_CsrPlugin_l1446) begin
        CsrPlugin_interrupt_code <= 4'b0111;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l1446_1) begin
        CsrPlugin_interrupt_code <= 4'b0011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l1446_2) begin
        CsrPlugin_interrupt_code <= 4'b1011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
    end
    if(when_CsrPlugin_l1534) begin
      if(when_CsrPlugin_l1542) begin
        case(CsrPlugin_targetPrivilege)
          2'b11 : begin
            CsrPlugin_mcause_interrupt <= (! CsrPlugin_hadException);
            CsrPlugin_mcause_exceptionCode <= CsrPlugin_trapCause;
            CsrPlugin_mepc <= writeBack_PC;
            if(CsrPlugin_hadException) begin
              CsrPlugin_mtval <= CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
            end
          end
          default : begin
          end
        endcase
      end else begin
        if(when_CsrPlugin_l1572) begin
          CsrPlugin_dpc <= writeBack_PC;
        end
      end
    end
    execute_MulPlugin_delayLogic_counter <= (execute_MulPlugin_delayLogic_counter + 1'b1);
    if(when_MulPlugin_l70) begin
      execute_MulPlugin_delayLogic_counter <= 1'b0;
    end
    execute_MulPlugin_withOuputBuffer_mul_ll <= (execute_MulPlugin_aULow * execute_MulPlugin_bULow);
    execute_MulPlugin_withOuputBuffer_mul_lh <= ($signed(execute_MulPlugin_aSLow) * $signed(execute_MulPlugin_bHigh));
    execute_MulPlugin_withOuputBuffer_mul_hl <= ($signed(execute_MulPlugin_aHigh) * $signed(execute_MulPlugin_bSLow));
    execute_MulPlugin_withOuputBuffer_mul_hh <= ($signed(execute_MulPlugin_aHigh) * $signed(execute_MulPlugin_bHigh));
    if(when_MulDivIterativePlugin_l126) begin
      memory_MulDivIterativePlugin_div_done <= 1'b1;
    end
    if(when_MulDivIterativePlugin_l126_1) begin
      memory_MulDivIterativePlugin_div_done <= 1'b0;
    end
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l132) begin
        memory_MulDivIterativePlugin_rs1[31 : 0] <= memory_MulDivIterativePlugin_div_stage_0_outNumerator;
        memory_MulDivIterativePlugin_accumulator[31 : 0] <= memory_MulDivIterativePlugin_div_stage_0_outRemainder;
        if(when_MulDivIterativePlugin_l151) begin
          memory_MulDivIterativePlugin_div_result <= _zz_memory_MulDivIterativePlugin_div_result_1[31:0];
        end
      end
    end
    if(when_MulDivIterativePlugin_l162) begin
      memory_MulDivIterativePlugin_accumulator <= 65'h0;
      memory_MulDivIterativePlugin_rs1 <= ((_zz_memory_MulDivIterativePlugin_rs1 ? (~ _zz_memory_MulDivIterativePlugin_rs1_1) : _zz_memory_MulDivIterativePlugin_rs1_1) + _zz_memory_MulDivIterativePlugin_rs1_2);
      memory_MulDivIterativePlugin_rs2 <= ((_zz_memory_MulDivIterativePlugin_rs2 ? (~ execute_RS2) : execute_RS2) + _zz_memory_MulDivIterativePlugin_rs2_1);
      memory_MulDivIterativePlugin_div_needRevert <= ((_zz_memory_MulDivIterativePlugin_rs1 ^ (_zz_memory_MulDivIterativePlugin_rs2 && (! execute_INSTRUCTION[13]))) && (! (((execute_RS2 == 32'h0) && execute_IS_RS2_SIGNED) && (! execute_INSTRUCTION[13]))));
    end
    if(writeBack_FpuPlugin_commit_ready) begin
      writeBack_FpuPlugin_commit_rData_opcode <= writeBack_FpuPlugin_commit_payload_opcode;
      writeBack_FpuPlugin_commit_rData_rd <= writeBack_FpuPlugin_commit_payload_rd;
      writeBack_FpuPlugin_commit_rData_write <= writeBack_FpuPlugin_commit_payload_write;
      writeBack_FpuPlugin_commit_rData_value <= writeBack_FpuPlugin_commit_payload_value;
    end
    if(CfuPlugin_bus_rsp_ready) begin
      CfuPlugin_bus_rsp_rData_outputs_0 <= CfuPlugin_bus_rsp_payload_outputs_0;
    end
    if(when_Pipeline_l124) begin
      decode_to_execute_PC <= _zz_decode_to_execute_PC;
    end
    if(when_Pipeline_l124_1) begin
      execute_to_memory_PC <= execute_PC;
    end
    if(when_Pipeline_l124_2) begin
      memory_to_writeBack_PC <= memory_PC;
    end
    if(when_Pipeline_l124_3) begin
      decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
    end
    if(when_Pipeline_l124_4) begin
      execute_to_memory_INSTRUCTION <= execute_INSTRUCTION;
    end
    if(when_Pipeline_l124_5) begin
      memory_to_writeBack_INSTRUCTION <= memory_INSTRUCTION;
    end
    if(when_Pipeline_l124_6) begin
      decode_to_execute_FORMAL_PC_NEXT <= decode_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_7) begin
      execute_to_memory_FORMAL_PC_NEXT <= execute_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_8) begin
      memory_to_writeBack_FORMAL_PC_NEXT <= _zz_memory_to_writeBack_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_9) begin
      decode_to_execute_MEMORY_FORCE_CONSTISTENCY <= decode_MEMORY_FORCE_CONSTISTENCY;
    end
    if(when_Pipeline_l124_10) begin
      decode_to_execute_LEGAL_INSTRUCTION <= decode_LEGAL_INSTRUCTION;
    end
    if(when_Pipeline_l124_11) begin
      decode_to_execute_MEMORY_FENCE_WR <= decode_MEMORY_FENCE_WR;
    end
    if(when_Pipeline_l124_12) begin
      decode_to_execute_SRC_USE_SUB_LESS <= decode_SRC_USE_SUB_LESS;
    end
    if(when_Pipeline_l124_13) begin
      decode_to_execute_MEMORY_ENABLE <= decode_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_14) begin
      execute_to_memory_MEMORY_ENABLE <= execute_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_15) begin
      memory_to_writeBack_MEMORY_ENABLE <= memory_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_16) begin
      decode_to_execute_ALU_CTRL <= _zz_decode_to_execute_ALU_CTRL;
    end
    if(when_Pipeline_l124_17) begin
      decode_to_execute_REGFILE_WRITE_VALID <= decode_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_18) begin
      execute_to_memory_REGFILE_WRITE_VALID <= execute_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_19) begin
      memory_to_writeBack_REGFILE_WRITE_VALID <= memory_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_20) begin
      decode_to_execute_BYPASSABLE_EXECUTE_STAGE <= decode_BYPASSABLE_EXECUTE_STAGE;
    end
    if(when_Pipeline_l124_21) begin
      decode_to_execute_BYPASSABLE_MEMORY_STAGE <= decode_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_22) begin
      execute_to_memory_BYPASSABLE_MEMORY_STAGE <= execute_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_23) begin
      decode_to_execute_MEMORY_WR <= decode_MEMORY_WR;
    end
    if(when_Pipeline_l124_24) begin
      execute_to_memory_MEMORY_WR <= execute_MEMORY_WR;
    end
    if(when_Pipeline_l124_25) begin
      memory_to_writeBack_MEMORY_WR <= memory_MEMORY_WR;
    end
    if(when_Pipeline_l124_26) begin
      decode_to_execute_HAS_SIDE_EFFECT <= decode_HAS_SIDE_EFFECT;
    end
    if(when_Pipeline_l124_27) begin
      execute_to_memory_HAS_SIDE_EFFECT <= execute_HAS_SIDE_EFFECT;
    end
    if(when_Pipeline_l124_28) begin
      memory_to_writeBack_HAS_SIDE_EFFECT <= memory_HAS_SIDE_EFFECT;
    end
    if(when_Pipeline_l124_29) begin
      decode_to_execute_MEMORY_LRSC <= decode_MEMORY_LRSC;
    end
    if(when_Pipeline_l124_30) begin
      execute_to_memory_MEMORY_LRSC <= execute_MEMORY_LRSC;
    end
    if(when_Pipeline_l124_31) begin
      memory_to_writeBack_MEMORY_LRSC <= memory_MEMORY_LRSC;
    end
    if(when_Pipeline_l124_32) begin
      decode_to_execute_MEMORY_AMO <= decode_MEMORY_AMO;
    end
    if(when_Pipeline_l124_33) begin
      execute_to_memory_MEMORY_AMO <= execute_MEMORY_AMO;
    end
    if(when_Pipeline_l124_34) begin
      memory_to_writeBack_MEMORY_AMO <= memory_MEMORY_AMO;
    end
    if(when_Pipeline_l124_35) begin
      decode_to_execute_MEMORY_MANAGMENT <= decode_MEMORY_MANAGMENT;
    end
    if(when_Pipeline_l124_36) begin
      decode_to_execute_MEMORY_FENCE <= decode_MEMORY_FENCE;
    end
    if(when_Pipeline_l124_37) begin
      execute_to_memory_MEMORY_FENCE <= execute_MEMORY_FENCE;
    end
    if(when_Pipeline_l124_38) begin
      memory_to_writeBack_MEMORY_FENCE <= memory_MEMORY_FENCE;
    end
    if(when_Pipeline_l124_39) begin
      decode_to_execute_IS_CSR <= decode_IS_CSR;
    end
    if(when_Pipeline_l124_40) begin
      decode_to_execute_ENV_CTRL <= _zz_decode_to_execute_ENV_CTRL;
    end
    if(when_Pipeline_l124_41) begin
      execute_to_memory_ENV_CTRL <= _zz_execute_to_memory_ENV_CTRL;
    end
    if(when_Pipeline_l124_42) begin
      memory_to_writeBack_ENV_CTRL <= _zz_memory_to_writeBack_ENV_CTRL;
    end
    if(when_Pipeline_l124_43) begin
      decode_to_execute_BRANCH_CTRL <= _zz_decode_to_execute_BRANCH_CTRL;
    end
    if(when_Pipeline_l124_44) begin
      decode_to_execute_SRC_LESS_UNSIGNED <= decode_SRC_LESS_UNSIGNED;
    end
    if(when_Pipeline_l124_45) begin
      decode_to_execute_IS_MUL <= decode_IS_MUL;
    end
    if(when_Pipeline_l124_46) begin
      execute_to_memory_IS_MUL <= execute_IS_MUL;
    end
    if(when_Pipeline_l124_47) begin
      memory_to_writeBack_IS_MUL <= memory_IS_MUL;
    end
    if(when_Pipeline_l124_48) begin
      decode_to_execute_IS_DIV <= decode_IS_DIV;
    end
    if(when_Pipeline_l124_49) begin
      execute_to_memory_IS_DIV <= execute_IS_DIV;
    end
    if(when_Pipeline_l124_50) begin
      decode_to_execute_IS_RS1_SIGNED <= decode_IS_RS1_SIGNED;
    end
    if(when_Pipeline_l124_51) begin
      decode_to_execute_IS_RS2_SIGNED <= decode_IS_RS2_SIGNED;
    end
    if(when_Pipeline_l124_52) begin
      decode_to_execute_FPU_COMMIT <= decode_FPU_COMMIT;
    end
    if(when_Pipeline_l124_53) begin
      execute_to_memory_FPU_COMMIT <= execute_FPU_COMMIT;
    end
    if(when_Pipeline_l124_54) begin
      memory_to_writeBack_FPU_COMMIT <= memory_FPU_COMMIT;
    end
    if(when_Pipeline_l124_55) begin
      decode_to_execute_FPU_RSP <= decode_FPU_RSP;
    end
    if(when_Pipeline_l124_56) begin
      execute_to_memory_FPU_RSP <= execute_FPU_RSP;
    end
    if(when_Pipeline_l124_57) begin
      memory_to_writeBack_FPU_RSP <= memory_FPU_RSP;
    end
    if(when_Pipeline_l124_58) begin
      decode_to_execute_FPU_OPCODE <= _zz_decode_to_execute_FPU_OPCODE;
    end
    if(when_Pipeline_l124_59) begin
      execute_to_memory_FPU_OPCODE <= _zz_execute_to_memory_FPU_OPCODE;
    end
    if(when_Pipeline_l124_60) begin
      memory_to_writeBack_FPU_OPCODE <= _zz_memory_to_writeBack_FPU_OPCODE;
    end
    if(when_Pipeline_l124_61) begin
      decode_to_execute_CfuPlugin_CFU_ENABLE <= decode_CfuPlugin_CFU_ENABLE;
    end
    if(when_Pipeline_l124_62) begin
      decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND <= _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
    end
    if(when_Pipeline_l124_63) begin
      decode_to_execute_ALU_BITWISE_CTRL <= _zz_decode_to_execute_ALU_BITWISE_CTRL;
    end
    if(when_Pipeline_l124_64) begin
      decode_to_execute_SHIFT_CTRL <= _zz_decode_to_execute_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_65) begin
      execute_to_memory_SHIFT_CTRL <= _zz_execute_to_memory_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_66) begin
      decode_to_execute_RS1 <= _zz_decode_to_execute_RS1;
    end
    if(when_Pipeline_l124_67) begin
      execute_to_memory_RS1 <= execute_RS1;
    end
    if(when_Pipeline_l124_68) begin
      memory_to_writeBack_RS1 <= memory_RS1;
    end
    if(when_Pipeline_l124_69) begin
      decode_to_execute_RS2 <= _zz_decode_to_execute_RS2;
    end
    if(when_Pipeline_l124_70) begin
      decode_to_execute_SRC2_FORCE_ZERO <= decode_SRC2_FORCE_ZERO;
    end
    if(when_Pipeline_l124_71) begin
      decode_to_execute_SRC1 <= decode_SRC1;
    end
    if(when_Pipeline_l124_72) begin
      decode_to_execute_SRC2 <= decode_SRC2;
    end
    if(when_Pipeline_l124_73) begin
      decode_to_execute_CSR_WRITE_OPCODE <= decode_CSR_WRITE_OPCODE;
    end
    if(when_Pipeline_l124_74) begin
      decode_to_execute_CSR_READ_OPCODE <= decode_CSR_READ_OPCODE;
    end
    if(when_Pipeline_l124_78) begin
      decode_to_execute_FPU_COMMIT_LOAD <= decode_FPU_COMMIT_LOAD;
    end
    if(when_Pipeline_l124_79) begin
      execute_to_memory_FPU_COMMIT_LOAD <= execute_FPU_COMMIT_LOAD;
    end
    if(when_Pipeline_l124_80) begin
      memory_to_writeBack_FPU_COMMIT_LOAD <= memory_FPU_COMMIT_LOAD;
    end
    if(when_Pipeline_l124_81) begin
      execute_to_memory_MEMORY_STORE_DATA_RF <= execute_MEMORY_STORE_DATA_RF;
    end
    if(when_Pipeline_l124_82) begin
      memory_to_writeBack_MEMORY_STORE_DATA_RF <= memory_MEMORY_STORE_DATA_RF;
    end
    if(when_Pipeline_l124_83) begin
      execute_to_memory_MEMORY_VIRTUAL_ADDRESS <= execute_MEMORY_VIRTUAL_ADDRESS;
    end
    if(when_Pipeline_l124_84) begin
      execute_to_memory_BRANCH_DO <= execute_BRANCH_DO;
    end
    if(when_Pipeline_l124_85) begin
      execute_to_memory_BRANCH_CALC <= execute_BRANCH_CALC;
    end
    if(when_Pipeline_l124_86) begin
      execute_to_memory_MUL_LL <= execute_MUL_LL;
    end
    if(when_Pipeline_l124_87) begin
      execute_to_memory_MUL_LH <= execute_MUL_LH;
    end
    if(when_Pipeline_l124_88) begin
      execute_to_memory_MUL_HL <= execute_MUL_HL;
    end
    if(when_Pipeline_l124_89) begin
      execute_to_memory_MUL_HH <= execute_MUL_HH;
    end
    if(when_Pipeline_l124_90) begin
      memory_to_writeBack_MUL_HH <= memory_MUL_HH;
    end
    if(when_Pipeline_l124_93) begin
      execute_to_memory_REGFILE_WRITE_DATA <= _zz_decode_RS2;
    end
    if(when_Pipeline_l124_94) begin
      memory_to_writeBack_REGFILE_WRITE_DATA <= _zz_decode_RS2_1;
    end
    if(when_Pipeline_l124_95) begin
      execute_to_memory_SHIFT_RIGHT <= execute_SHIFT_RIGHT;
    end
    if(when_Pipeline_l124_96) begin
      memory_to_writeBack_MUL_LOW <= memory_MUL_LOW;
    end
    if(when_Fetcher_l411) begin
      _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst <= CsrPlugin_injectionPort_payload;
    end
    if(when_CsrPlugin_l1813) begin
      execute_CsrPlugin_csr_1972 <= (decode_INSTRUCTION[31 : 20] == 12'h7b4);
    end
    if(when_CsrPlugin_l1813_1) begin
      execute_CsrPlugin_csr_1969 <= (decode_INSTRUCTION[31 : 20] == 12'h7b1);
    end
    if(when_CsrPlugin_l1813_2) begin
      execute_CsrPlugin_csr_1968 <= (decode_INSTRUCTION[31 : 20] == 12'h7b0);
    end
    if(when_CsrPlugin_l1813_3) begin
      execute_CsrPlugin_csr_3857 <= (decode_INSTRUCTION[31 : 20] == 12'hf11);
    end
    if(when_CsrPlugin_l1813_4) begin
      execute_CsrPlugin_csr_3858 <= (decode_INSTRUCTION[31 : 20] == 12'hf12);
    end
    if(when_CsrPlugin_l1813_5) begin
      execute_CsrPlugin_csr_3859 <= (decode_INSTRUCTION[31 : 20] == 12'hf13);
    end
    if(when_CsrPlugin_l1813_6) begin
      execute_CsrPlugin_csr_3860 <= (decode_INSTRUCTION[31 : 20] == 12'hf14);
    end
    if(when_CsrPlugin_l1813_7) begin
      execute_CsrPlugin_csr_769 <= (decode_INSTRUCTION[31 : 20] == 12'h301);
    end
    if(when_CsrPlugin_l1813_8) begin
      execute_CsrPlugin_csr_768 <= (decode_INSTRUCTION[31 : 20] == 12'h300);
    end
    if(when_CsrPlugin_l1813_9) begin
      execute_CsrPlugin_csr_836 <= (decode_INSTRUCTION[31 : 20] == 12'h344);
    end
    if(when_CsrPlugin_l1813_10) begin
      execute_CsrPlugin_csr_772 <= (decode_INSTRUCTION[31 : 20] == 12'h304);
    end
    if(when_CsrPlugin_l1813_11) begin
      execute_CsrPlugin_csr_773 <= (decode_INSTRUCTION[31 : 20] == 12'h305);
    end
    if(when_CsrPlugin_l1813_12) begin
      execute_CsrPlugin_csr_833 <= (decode_INSTRUCTION[31 : 20] == 12'h341);
    end
    if(when_CsrPlugin_l1813_13) begin
      execute_CsrPlugin_csr_832 <= (decode_INSTRUCTION[31 : 20] == 12'h340);
    end
    if(when_CsrPlugin_l1813_14) begin
      execute_CsrPlugin_csr_834 <= (decode_INSTRUCTION[31 : 20] == 12'h342);
    end
    if(when_CsrPlugin_l1813_15) begin
      execute_CsrPlugin_csr_835 <= (decode_INSTRUCTION[31 : 20] == 12'h343);
    end
    if(when_CsrPlugin_l1813_16) begin
      execute_CsrPlugin_csr_3 <= (decode_INSTRUCTION[31 : 20] == 12'h003);
    end
    if(when_CsrPlugin_l1813_17) begin
      execute_CsrPlugin_csr_2 <= (decode_INSTRUCTION[31 : 20] == 12'h002);
    end
    if(when_CsrPlugin_l1813_18) begin
      execute_CsrPlugin_csr_1 <= (decode_INSTRUCTION[31 : 20] == 12'h001);
    end
    if(when_CsrPlugin_l1813_19) begin
      execute_CsrPlugin_csr_256 <= (decode_INSTRUCTION[31 : 20] == 12'h100);
    end
    if(execute_CsrPlugin_csr_1969) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_dpc <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    if(execute_CsrPlugin_csr_836) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mip_MSIP <= CsrPlugin_csrMapping_writeDataSignal[3];
      end
    end
    if(execute_CsrPlugin_csr_773) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mtvec_base <= CsrPlugin_csrMapping_writeDataSignal[31 : 2];
      end
    end
    if(execute_CsrPlugin_csr_833) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mepc <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    if(execute_CsrPlugin_csr_832) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mscratch <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
  end


endmodule

module VexRiscv (
  output wire          dBus_cmd_valid,
  input  wire          dBus_cmd_ready,
  output wire          dBus_cmd_payload_wr,
  output wire          dBus_cmd_payload_uncached,
  output wire [31:0]   dBus_cmd_payload_address,
  output wire [63:0]   dBus_cmd_payload_data,
  output wire [7:0]    dBus_cmd_payload_mask,
  output wire [2:0]    dBus_cmd_payload_size,
  output wire          dBus_cmd_payload_exclusive,
  output wire          dBus_cmd_payload_last,
  input  wire          dBus_rsp_valid,
  input  wire [3:0]    dBus_rsp_payload_aggregated,
  input  wire          dBus_rsp_payload_last,
  input  wire [63:0]   dBus_rsp_payload_data,
  input  wire          dBus_rsp_payload_error,
  input  wire          dBus_rsp_payload_exclusive,
  input  wire          dBus_inv_valid,
  output wire          dBus_inv_ready,
  input  wire          dBus_inv_payload_last,
  input  wire          dBus_inv_payload_fragment_enable,
  input  wire [31:0]   dBus_inv_payload_fragment_address,
  output wire          dBus_ack_valid,
  input  wire          dBus_ack_ready,
  output wire          dBus_ack_payload_last,
  output wire          dBus_ack_payload_fragment_hit,
  input  wire          dBus_sync_valid,
  output wire          dBus_sync_ready,
  input  wire [3:0]    dBus_sync_payload_aggregated,
  input  wire          timerInterrupt,
  input  wire          externalInterrupt,
  input  wire          softwareInterrupt,
  output wire          debugBus_halted,
  output wire          debugBus_running,
  output wire          debugBus_unavailable,
  output reg           debugBus_exception,
  output wire          debugBus_commit,
  output reg           debugBus_ebreak,
  output wire          debugBus_redo,
  output wire          debugBus_regSuccess,
  input  wire          debugBus_ackReset,
  output wire          debugBus_haveReset,
  input  wire          debugBus_resume_cmd_valid,
  output reg           debugBus_resume_rsp_valid,
  input  wire          debugBus_haltReq,
  input  wire          debugBus_dmToHart_valid,
  input  wire [1:0]    debugBus_dmToHart_payload_op,
  input  wire [4:0]    debugBus_dmToHart_payload_address,
  input  wire [31:0]   debugBus_dmToHart_payload_data,
  input  wire [2:0]    debugBus_dmToHart_payload_size,
  output reg           debugBus_hartToDm_valid,
  output reg  [3:0]    debugBus_hartToDm_payload_address,
  output reg  [31:0]   debugBus_hartToDm_payload_data,
  output reg           FpuPlugin_port_cmd_valid /* verilator public */ ,
  input  wire          FpuPlugin_port_cmd_ready /* verilator public */ ,
  output reg  [3:0]    FpuPlugin_port_cmd_payload_opcode /* verilator public */ ,
  output wire [1:0]    FpuPlugin_port_cmd_payload_arg /* verilator public */ ,
  output wire [4:0]    FpuPlugin_port_cmd_payload_rs1 /* verilator public */ ,
  output reg  [4:0]    FpuPlugin_port_cmd_payload_rs2 /* verilator public */ ,
  output wire [4:0]    FpuPlugin_port_cmd_payload_rs3 /* verilator public */ ,
  output reg  [4:0]    FpuPlugin_port_cmd_payload_rd /* verilator public */ ,
  output reg  [0:0]    FpuPlugin_port_cmd_payload_format /* verilator public */ ,
  output wire [2:0]    FpuPlugin_port_cmd_payload_roundMode /* verilator public */ ,
  output reg           FpuPlugin_port_commit_valid /* verilator public */ ,
  input  wire          FpuPlugin_port_commit_ready /* verilator public */ ,
  output reg  [3:0]    FpuPlugin_port_commit_payload_opcode /* verilator public */ ,
  output reg  [4:0]    FpuPlugin_port_commit_payload_rd /* verilator public */ ,
  output reg           FpuPlugin_port_commit_payload_write /* verilator public */ ,
  output reg  [63:0]   FpuPlugin_port_commit_payload_value /* verilator public */ ,
  input  wire          FpuPlugin_port_rsp_valid /* verilator public */ ,
  output reg           FpuPlugin_port_rsp_ready /* verilator public */ ,
  input  wire [63:0]   FpuPlugin_port_rsp_payload_value /* verilator public */ ,
  input  wire          FpuPlugin_port_rsp_payload_NV /* verilator public */ ,
  input  wire          FpuPlugin_port_rsp_payload_NX /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_valid /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_NX /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_UF /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_OF /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_DZ /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_flags_NV /* verilator public */ ,
  input  wire          FpuPlugin_port_completion_payload_written /* verilator public */ ,
  output wire          CfuPlugin_bus_cmd_valid,
  input  wire          CfuPlugin_bus_cmd_ready,
  output wire [9:0]    CfuPlugin_bus_cmd_payload_function_id,
  output wire [31:0]   CfuPlugin_bus_cmd_payload_inputs_0,
  output wire [31:0]   CfuPlugin_bus_cmd_payload_inputs_1,
  input  wire          CfuPlugin_bus_rsp_valid,
  output wire          CfuPlugin_bus_rsp_ready,
  input  wire [31:0]   CfuPlugin_bus_rsp_payload_outputs_0,
  output wire          iBus_cmd_valid,
  input  wire          iBus_cmd_ready,
  output reg  [31:0]   iBus_cmd_payload_address,
  output wire [2:0]    iBus_cmd_payload_size,
  input  wire          iBus_rsp_valid,
  input  wire [63:0]   iBus_rsp_payload_data,
  input  wire          iBus_rsp_payload_error,
  input  wire          systemCd_logic_outputReset,
  output reg           stoptime,
  input  wire          io_systemClk
);
  localparam FpuOpcode_LOAD = 4'd0;
  localparam FpuOpcode_STORE = 4'd1;
  localparam FpuOpcode_MUL = 4'd2;
  localparam FpuOpcode_ADD = 4'd3;
  localparam FpuOpcode_FMA = 4'd4;
  localparam FpuOpcode_I2F = 4'd5;
  localparam FpuOpcode_F2I = 4'd6;
  localparam FpuOpcode_CMP = 4'd7;
  localparam FpuOpcode_DIV = 4'd8;
  localparam FpuOpcode_SQRT = 4'd9;
  localparam FpuOpcode_MIN_MAX = 4'd10;
  localparam FpuOpcode_SGNJ = 4'd11;
  localparam FpuOpcode_FMV_X_W = 4'd12;
  localparam FpuOpcode_FMV_W_X = 4'd13;
  localparam FpuOpcode_FCLASS = 4'd14;
  localparam FpuOpcode_FCVT_X_X = 4'd15;
  localparam ShiftCtrlEnum_DISABLE_1 = 2'd0;
  localparam ShiftCtrlEnum_SLL_1 = 2'd1;
  localparam ShiftCtrlEnum_SRL_1 = 2'd2;
  localparam ShiftCtrlEnum_SRA_1 = 2'd3;
  localparam AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam Input2Kind_RS = 1'd0;
  localparam Input2Kind_IMM_I = 1'd1;
  localparam BranchCtrlEnum_INC = 2'd0;
  localparam BranchCtrlEnum_B = 2'd1;
  localparam BranchCtrlEnum_JAL = 2'd2;
  localparam BranchCtrlEnum_JALR = 2'd3;
  localparam EnvCtrlEnum_NONE = 2'd0;
  localparam EnvCtrlEnum_XRET = 2'd1;
  localparam EnvCtrlEnum_ECALL = 2'd2;
  localparam EnvCtrlEnum_EBREAK = 2'd3;
  localparam AluCtrlEnum_ADD_SUB = 2'd0;
  localparam AluCtrlEnum_SLT_SLTU = 2'd1;
  localparam AluCtrlEnum_BITWISE = 2'd2;
  localparam FpuFormat_FLOAT = 1'd0;
  localparam FpuFormat_DOUBLE = 1'd1;
  localparam Src2CtrlEnum_RS = 2'd0;
  localparam Src2CtrlEnum_IMI = 2'd1;
  localparam Src2CtrlEnum_IMS = 2'd2;
  localparam Src2CtrlEnum_PC = 2'd3;
  localparam Src1CtrlEnum_RS = 2'd0;
  localparam Src1CtrlEnum_IMU = 2'd1;
  localparam Src1CtrlEnum_PC_INCREMENT = 2'd2;
  localparam Src1CtrlEnum_URS1 = 2'd3;
  localparam DebugDmToHartOp_DATA = 2'd0;
  localparam DebugDmToHartOp_EXECUTE = 2'd1;
  localparam DebugDmToHartOp_REG_WRITE = 2'd2;
  localparam DebugDmToHartOp_REG_READ = 2'd3;
  localparam FpuRoundMode_RNE = 3'd0;
  localparam FpuRoundMode_RTZ = 3'd1;
  localparam FpuRoundMode_RDN = 3'd2;
  localparam FpuRoundMode_RUP = 3'd3;
  localparam FpuRoundMode_RMM = 3'd4;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_BOOT = 2'd0;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_IDLE = 2'd1;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_SINGLE = 2'd2;
  localparam CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 = 2'd3;
  localparam FpuPlugin_enumDef_BOOT = 3'd0;
  localparam FpuPlugin_enumDef_IDLE = 3'd1;
  localparam FpuPlugin_enumDef_CMD = 3'd2;
  localparam FpuPlugin_enumDef_RSP = 3'd3;
  localparam FpuPlugin_enumDef_RSP_0 = 3'd4;
  localparam FpuPlugin_enumDef_RSP_1 = 3'd5;
  localparam FpuPlugin_enumDef_COMMIT = 3'd6;
  localparam FpuPlugin_enumDef_DONE = 3'd7;

  wire                IBusCachedPlugin_cache_io_flush;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isRemoved;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isUser;
  reg                 IBusCachedPlugin_cache_io_cpu_fill_valid;
  wire                dataCache_2_io_cpu_execute_isValid;
  wire       [31:0]   dataCache_2_io_cpu_execute_address;
  reg                 dataCache_2_io_cpu_execute_args_isLrsc;
  wire                dataCache_2_io_cpu_execute_args_amoCtrl_swap;
  wire       [2:0]    dataCache_2_io_cpu_execute_args_amoCtrl_alu;
  wire                dataCache_2_io_cpu_memory_isValid;
  reg                 dataCache_2_io_cpu_memory_mmuRsp_isIoAccess;
  reg                 dataCache_2_io_cpu_writeBack_isValid;
  wire                dataCache_2_io_cpu_writeBack_isUser;
  reg        [63:0]   dataCache_2_io_cpu_writeBack_storeData;
  wire       [31:0]   dataCache_2_io_cpu_writeBack_address;
  reg                 dataCache_2_io_cpu_writeBack_fence_SW;
  reg                 dataCache_2_io_cpu_writeBack_fence_SR;
  reg                 dataCache_2_io_cpu_writeBack_fence_SO;
  reg                 dataCache_2_io_cpu_writeBack_fence_SI;
  reg                 dataCache_2_io_cpu_writeBack_fence_PW;
  reg                 dataCache_2_io_cpu_writeBack_fence_PR;
  reg                 dataCache_2_io_cpu_writeBack_fence_PO;
  reg                 dataCache_2_io_cpu_writeBack_fence_PI;
  wire       [3:0]    dataCache_2_io_cpu_writeBack_fence_FM;
  wire                dataCache_2_io_cpu_flush_valid;
  wire                dataCache_2_io_cpu_flush_payload_singleLine;
  wire       [5:0]    dataCache_2_io_cpu_flush_payload_lineId;
  reg        [31:0]   RegFilePlugin_regFile_spinal_port0;
  reg        [31:0]   RegFilePlugin_regFile_spinal_port1;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_haltIt;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_data;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress;
  wire                IBusCachedPlugin_cache_io_cpu_decode_error;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuException;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_data;
  wire                IBusCachedPlugin_cache_io_cpu_decode_cacheMiss;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_physicalAddress;
  wire                IBusCachedPlugin_cache_io_mem_cmd_valid;
  wire       [31:0]   IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  wire       [2:0]    IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  wire                dataCache_2_io_cpu_execute_haltIt;
  wire                dataCache_2_io_cpu_execute_refilling;
  wire                dataCache_2_io_cpu_memory_isWrite;
  wire                dataCache_2_io_cpu_writeBack_haltIt;
  wire       [63:0]   dataCache_2_io_cpu_writeBack_data;
  wire                dataCache_2_io_cpu_writeBack_mmuException;
  wire                dataCache_2_io_cpu_writeBack_unalignedAccess;
  wire                dataCache_2_io_cpu_writeBack_accessError;
  wire                dataCache_2_io_cpu_writeBack_isWrite;
  wire                dataCache_2_io_cpu_writeBack_keepMemRspData;
  wire                dataCache_2_io_cpu_writeBack_exclusiveOk;
  wire                dataCache_2_io_cpu_flush_ready;
  wire                dataCache_2_io_cpu_redo;
  wire                dataCache_2_io_cpu_writesPending;
  wire                dataCache_2_io_mem_cmd_valid;
  wire                dataCache_2_io_mem_cmd_payload_wr;
  wire                dataCache_2_io_mem_cmd_payload_uncached;
  wire       [31:0]   dataCache_2_io_mem_cmd_payload_address;
  wire       [63:0]   dataCache_2_io_mem_cmd_payload_data;
  wire       [7:0]    dataCache_2_io_mem_cmd_payload_mask;
  wire       [2:0]    dataCache_2_io_mem_cmd_payload_size;
  wire                dataCache_2_io_mem_cmd_payload_exclusive;
  wire                dataCache_2_io_mem_cmd_payload_last;
  wire                dataCache_2_io_mem_inv_ready;
  wire                dataCache_2_io_mem_ack_valid;
  wire                dataCache_2_io_mem_ack_payload_last;
  wire                dataCache_2_io_mem_ack_payload_fragment_hit;
  wire                dataCache_2_io_mem_sync_ready;
  wire                systemCd_logic_outputReset_buffercc_io_dataOut;
  wire       [31:0]   EfxCPUSp1_inst_result;
  wire       [31:0]   EfxCPUSp2_inst_result;
  wire       [51:0]   _zz_memory_MUL_LOW;
  wire       [51:0]   _zz_memory_MUL_LOW_1;
  wire       [51:0]   _zz_memory_MUL_LOW_2;
  wire       [32:0]   _zz_memory_MUL_LOW_3;
  wire       [51:0]   _zz_memory_MUL_LOW_4;
  wire       [49:0]   _zz_memory_MUL_LOW_5;
  wire       [51:0]   _zz_memory_MUL_LOW_6;
  wire       [49:0]   _zz_memory_MUL_LOW_7;
  wire       [31:0]   _zz_decode_FORMAL_PC_NEXT;
  wire       [2:0]    _zz_decode_FORMAL_PC_NEXT_1;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_1;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_2;
  wire                _zz_decode_LEGAL_INSTRUCTION_3;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_4;
  wire       [29:0]   _zz_decode_LEGAL_INSTRUCTION_5;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_6;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_7;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_8;
  wire                _zz_decode_LEGAL_INSTRUCTION_9;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_10;
  wire       [23:0]   _zz_decode_LEGAL_INSTRUCTION_11;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_12;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_13;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_14;
  wire                _zz_decode_LEGAL_INSTRUCTION_15;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_16;
  wire       [17:0]   _zz_decode_LEGAL_INSTRUCTION_17;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_18;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_19;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_20;
  wire                _zz_decode_LEGAL_INSTRUCTION_21;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_22;
  wire       [11:0]   _zz_decode_LEGAL_INSTRUCTION_23;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_24;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_25;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_26;
  wire                _zz_decode_LEGAL_INSTRUCTION_27;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_28;
  wire       [5:0]    _zz_decode_LEGAL_INSTRUCTION_29;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_30;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_31;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_32;
  wire                _zz_decode_LEGAL_INSTRUCTION_33;
  wire                _zz_decode_LEGAL_INSTRUCTION_34;
  wire       [2:0]    _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  reg        [31:0]   _zz_IBusCachedPlugin_jump_pcLoad_payload_4;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_5;
  wire       [31:0]   _zz_IBusCachedPlugin_fetchPc_pc;
  wire       [2:0]    _zz_IBusCachedPlugin_fetchPc_pc_1;
  wire       [31:0]   _zz_IBusCachedPlugin_decodePc_pcPlus;
  wire       [2:0]    _zz_IBusCachedPlugin_decodePc_pcPlus_1;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_28;
  wire       [0:0]    _zz_IBusCachedPlugin_decompressor_decompressed_29;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_30;
  wire       [31:0]   _zz_IBusCachedPlugin_decompressor_decompressed_31;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_32;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_33;
  wire       [6:0]    _zz_IBusCachedPlugin_decompressor_decompressed_34;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_35;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_36;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_37;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_38;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_39;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_40;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_41;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_42;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_43;
  wire       [25:0]   _zz_io_cpu_flush_payload_lineId;
  wire       [25:0]   _zz_io_cpu_flush_payload_lineId_1;
  wire       [2:0]    _zz_DBusCachedPlugin_exceptionBus_payload_code;
  wire       [2:0]    _zz_DBusCachedPlugin_exceptionBus_payload_code_1;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted;
  wire       [2:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_1;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_2;
  wire       [1:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_3;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_4;
  wire       [0:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_5;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_6;
  wire       [0:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_7;
  wire       [0:0]    _zz_writeBack_DBusCachedPlugin_rspRf;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_1;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_2;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_3;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_4;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_5;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_6;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_7;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_8;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_9;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_10;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_11;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_12;
  wire       [40:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_13;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_14;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_15;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_16;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_17;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_18;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_19;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_20;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_21;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_22;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_23;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_24;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_25;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_26;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_27;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_28;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_29;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_30;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_31;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_32;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_33;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_34;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_35;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_36;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_37;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_38;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_39;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_40;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_41;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_42;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_43;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_44;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_45;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_46;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_47;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_48;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_49;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_50;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_51;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_52;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_53;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_54;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_55;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_56;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_57;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_58;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_59;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_60;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_61;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_62;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_63;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_64;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_65;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_66;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_67;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_68;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_69;
  wire       [35:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_70;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_71;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_72;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_73;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_74;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_75;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_76;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_77;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_78;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_79;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_80;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_81;
  wire       [33:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_82;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_83;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_84;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_85;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_86;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_87;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_88;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_89;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_90;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_91;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_92;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_93;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_94;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_95;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_96;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_97;
  wire       [29:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_98;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_99;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_100;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_101;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_102;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_103;
  wire       [27:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_104;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_105;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_106;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_107;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_108;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_109;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_110;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_111;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_112;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_113;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_114;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_115;
  wire       [24:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_116;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_117;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_118;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_119;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_120;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_121;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_122;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_123;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_124;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_125;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_126;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_127;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_128;
  wire       [20:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_129;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_130;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_131;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_132;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_133;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_134;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_135;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_136;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_137;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_138;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_139;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_140;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_141;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_142;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_143;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_144;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_145;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_146;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_147;
  wire       [16:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_148;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_149;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_150;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_151;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_152;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_153;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_154;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_155;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_156;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_157;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_158;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_159;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_160;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_161;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_162;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_163;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_164;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_165;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_166;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_167;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_168;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_169;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_170;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_171;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_172;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_173;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_174;
  wire       [13:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_175;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_176;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_177;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_178;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_179;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_180;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_181;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_182;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_183;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_184;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_185;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_186;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_187;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_188;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_189;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_190;
  wire       [3:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_191;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_192;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_193;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_194;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_195;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_196;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_197;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_198;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_199;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_200;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_201;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_202;
  wire       [6:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_203;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_204;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_205;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_206;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_207;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_208;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_209;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_210;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_211;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_212;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_213;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_214;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_215;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_216;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_217;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_218;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_219;
  wire       [10:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_220;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_221;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_222;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_223;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_224;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_225;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_226;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_227;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_228;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_229;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_230;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_231;
  wire       [8:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_232;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_233;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_234;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_235;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_236;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_237;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_238;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_239;
  wire       [6:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_240;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_241;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_242;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_243;
  wire       [5:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_244;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_245;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_246;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_247;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_248;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_249;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_250;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_251;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_252;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_253;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_254;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_255;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_256;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_257;
  wire       [4:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_258;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_259;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_260;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_261;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_262;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_263;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_264;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_265;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_266;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_267;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_268;
  wire       [0:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_269;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_270;
  wire       [31:0]   _zz__zz_decode_CfuPlugin_CFU_ENABLE_271;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_272;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_273;
  wire       [2:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_274;
  wire       [1:0]    _zz__zz_decode_CfuPlugin_CFU_ENABLE_275;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_276;
  wire                _zz__zz_decode_CfuPlugin_CFU_ENABLE_277;
  wire                _zz_RegFilePlugin_regFile_port;
  wire                _zz_decode_RegFilePlugin_rs1Data;
  wire                _zz_RegFilePlugin_regFile_port_1;
  wire                _zz_decode_RegFilePlugin_rs2Data;
  wire       [2:0]    _zz__zz_decode_SRC1;
  wire       [4:0]    _zz__zz_decode_SRC1_1;
  wire       [11:0]   _zz__zz_decode_SRC2_2;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_1;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_2;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_4;
  wire       [2:0]    _zz_CsrPlugin_timeout_counter_valueNext;
  wire       [0:0]    _zz_CsrPlugin_timeout_counter_valueNext_1;
  wire       [0:0]    _zz__zz_6;
  wire       [63:0]   _zz_CsrPlugin_counters_mcycle;
  wire       [0:0]    _zz_CsrPlugin_counters_mcycle_1;
  wire       [63:0]   _zz_CsrPlugin_counters_minstret;
  wire       [0:0]    _zz_CsrPlugin_counters_minstret_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1;
  wire                _zz_when;
  wire       [19:0]   _zz__zz_execute_BranchPlugin_branch_src2;
  wire       [11:0]   _zz__zz_execute_BranchPlugin_branch_src2_4;
  wire       [65:0]   _zz_writeBack_MulPlugin_result;
  wire       [65:0]   _zz_writeBack_MulPlugin_result_1;
  wire       [31:0]   _zz__zz_decode_RS2_2;
  wire       [31:0]   _zz__zz_decode_RS2_2_1;
  wire       [5:0]    _zz_memory_MulDivIterativePlugin_div_counter_valueNext;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_div_counter_valueNext_1;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder_1;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_outNumerator;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_1;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_2;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_3;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_div_result_4;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_div_result_5;
  wire       [32:0]   _zz_memory_MulDivIterativePlugin_rs1_2;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_rs1_3;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_rs2_1;
  wire       [0:0]    _zz_memory_MulDivIterativePlugin_rs2_2;
  wire       [5:0]    _zz_FpuPlugin_pendings;
  wire       [5:0]    _zz_FpuPlugin_pendings_1;
  wire       [5:0]    _zz_FpuPlugin_pendings_2;
  wire       [0:0]    _zz_FpuPlugin_pendings_3;
  wire       [5:0]    _zz_FpuPlugin_pendings_4;
  wire       [0:0]    _zz_FpuPlugin_pendings_5;
  wire       [5:0]    _zz_FpuPlugin_pendings_6;
  wire       [0:0]    _zz_FpuPlugin_pendings_7;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_16;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_17;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_18;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_19;
  wire       [7:0]    _zz_when_CsrPlugin_l1862;
  wire       [63:0]   writeBack_MEMORY_LOAD_DATA;
  wire       [51:0]   memory_MUL_LOW;
  wire       [31:0]   execute_SHIFT_RIGHT;
  wire       [31:0]   execute_REGFILE_WRITE_DATA;
  wire                memory_CfuPlugin_CFU_IN_FLIGHT;
  wire                execute_CfuPlugin_CFU_IN_FLIGHT;
  wire       [33:0]   memory_MUL_HH;
  wire       [33:0]   execute_MUL_HH;
  wire       [33:0]   execute_MUL_HL;
  wire       [33:0]   execute_MUL_LH;
  wire       [31:0]   execute_MUL_LL;
  wire       [31:0]   execute_BRANCH_CALC;
  wire                execute_BRANCH_DO;
  wire       [31:0]   execute_MEMORY_VIRTUAL_ADDRESS;
  wire       [31:0]   execute_MEMORY_STORE_DATA_RF;
  wire                memory_FPU_COMMIT_LOAD;
  wire                execute_FPU_COMMIT_LOAD;
  wire                decode_FPU_COMMIT_LOAD;
  wire                memory_FPU_FORKED;
  wire                execute_FPU_FORKED;
  wire                decode_FPU_FORKED;
  wire                decode_CSR_READ_OPCODE;
  wire                decode_CSR_WRITE_OPCODE;
  wire       [31:0]   decode_SRC2;
  wire       [31:0]   decode_SRC1;
  wire                decode_SRC2_FORCE_ZERO;
  wire       [31:0]   memory_RS1;
  wire       [1:0]    _zz_execute_to_memory_SHIFT_CTRL;
  wire       [1:0]    _zz_execute_to_memory_SHIFT_CTRL_1;
  wire       [1:0]    decode_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SHIFT_CTRL_1;
  wire       [1:0]    decode_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  wire       [0:0]    decode_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_decode_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1;
  wire                decode_CfuPlugin_CFU_ENABLE;
  wire       [3:0]    memory_FPU_OPCODE;
  wire       [3:0]    _zz_memory_FPU_OPCODE;
  wire       [3:0]    _zz_memory_to_writeBack_FPU_OPCODE;
  wire       [3:0]    _zz_memory_to_writeBack_FPU_OPCODE_1;
  wire       [3:0]    execute_FPU_OPCODE;
  wire       [3:0]    _zz_execute_FPU_OPCODE;
  wire       [3:0]    _zz_execute_to_memory_FPU_OPCODE;
  wire       [3:0]    _zz_execute_to_memory_FPU_OPCODE_1;
  wire       [3:0]    _zz_decode_to_execute_FPU_OPCODE;
  wire       [3:0]    _zz_decode_to_execute_FPU_OPCODE_1;
  wire                memory_FPU_RSP;
  wire                execute_FPU_RSP;
  wire                decode_FPU_RSP;
  wire                memory_FPU_COMMIT;
  wire                execute_FPU_COMMIT;
  wire                decode_FPU_COMMIT;
  wire                decode_IS_RS2_SIGNED;
  wire                decode_IS_RS1_SIGNED;
  wire                decode_IS_DIV;
  wire                memory_IS_MUL;
  wire                decode_IS_MUL;
  wire                decode_SRC_LESS_UNSIGNED;
  wire       [1:0]    decode_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_to_execute_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_to_execute_BRANCH_CTRL_1;
  wire       [1:0]    _zz_memory_to_writeBack_ENV_CTRL;
  wire       [1:0]    _zz_memory_to_writeBack_ENV_CTRL_1;
  wire       [1:0]    _zz_execute_to_memory_ENV_CTRL;
  wire       [1:0]    _zz_execute_to_memory_ENV_CTRL_1;
  wire       [1:0]    decode_ENV_CTRL;
  wire       [1:0]    _zz_decode_ENV_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ENV_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ENV_CTRL_1;
  wire                decode_IS_CSR;
  wire                memory_MEMORY_FENCE;
  wire                execute_MEMORY_FENCE;
  wire                decode_MEMORY_FENCE;
  wire                decode_MEMORY_MANAGMENT;
  wire                memory_MEMORY_AMO;
  wire                memory_MEMORY_LRSC;
  wire                execute_HAS_SIDE_EFFECT;
  wire                decode_HAS_SIDE_EFFECT;
  wire                decode_MEMORY_WR;
  wire                execute_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_EXECUTE_STAGE;
  wire       [1:0]    decode_ALU_CTRL;
  wire       [1:0]    _zz_decode_ALU_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_CTRL_1;
  wire                decode_MEMORY_FENCE_WR;
  wire                decode_MEMORY_FORCE_CONSTISTENCY;
  wire       [31:0]   writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   memory_FORMAL_PC_NEXT;
  wire       [31:0]   execute_FORMAL_PC_NEXT;
  wire       [31:0]   decode_FORMAL_PC_NEXT;
  wire       [31:0]   memory_SHIFT_RIGHT;
  wire       [1:0]    memory_SHIFT_CTRL;
  wire       [1:0]    _zz_memory_SHIFT_CTRL;
  wire       [1:0]    execute_SHIFT_CTRL;
  wire       [1:0]    _zz_execute_SHIFT_CTRL;
  wire       [31:0]   execute_SRC_ADD_SUB;
  wire       [1:0]    execute_ALU_CTRL;
  wire       [1:0]    _zz_execute_ALU_CTRL;
  wire       [1:0]    execute_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_execute_ALU_BITWISE_CTRL;
  reg                 _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
  reg                 _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
  wire                writeBack_CfuPlugin_CFU_IN_FLIGHT;
  wire       [0:0]    execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire       [0:0]    _zz_execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire                writeBack_HAS_SIDE_EFFECT;
  wire                memory_HAS_SIDE_EFFECT;
  wire                execute_LEGAL_INSTRUCTION;
  reg                 execute_CfuPlugin_CFU_ENABLE;
  reg                 _zz_memory_to_writeBack_FPU_FORKED;
  reg                 _zz_execute_to_memory_FPU_FORKED;
  reg                 _zz_decode_to_execute_FPU_FORKED;
  wire       [3:0]    writeBack_FPU_OPCODE;
  wire       [3:0]    _zz_writeBack_FPU_OPCODE;
  wire       [31:0]   writeBack_RS1;
  wire       [63:0]   _zz_writeBack_FpuPlugin_commit_payload_value;
  wire                writeBack_FPU_COMMIT_LOAD;
  reg                 DBusBypass0_cond;
  wire                writeBack_FPU_COMMIT;
  wire                writeBack_FPU_RSP;
  wire                writeBack_FPU_FORKED;
  wire       [0:0]    decode_FPU_FORMAT;
  wire       [0:0]    _zz_decode_FPU_FORMAT;
  wire       [1:0]    decode_FPU_ARG;
  wire       [3:0]    decode_FPU_OPCODE;
  wire       [3:0]    _zz_decode_FPU_OPCODE;
  reg                 decode_FPU_ENABLE;
  wire                execute_IS_RS1_SIGNED;
  wire                execute_IS_DIV;
  wire                execute_IS_RS2_SIGNED;
  wire                memory_IS_DIV;
  wire                writeBack_IS_MUL;
  wire       [33:0]   writeBack_MUL_HH;
  wire       [51:0]   writeBack_MUL_LOW;
  wire       [33:0]   memory_MUL_HL;
  wire       [33:0]   memory_MUL_LH;
  wire       [31:0]   memory_MUL_LL;
  wire                execute_IS_MUL;
  wire       [31:0]   memory_BRANCH_CALC;
  wire                memory_BRANCH_DO;
  wire       [31:0]   execute_PC;
  wire       [1:0]    execute_BRANCH_CTRL;
  wire       [1:0]    _zz_execute_BRANCH_CTRL;
  wire                execute_SRC_LESS;
  wire                execute_CSR_READ_OPCODE;
  wire                execute_CSR_WRITE_OPCODE;
  wire                execute_IS_CSR;
  wire       [1:0]    memory_ENV_CTRL;
  wire       [1:0]    _zz_memory_ENV_CTRL;
  wire       [1:0]    execute_ENV_CTRL;
  wire       [1:0]    _zz_execute_ENV_CTRL;
  wire       [1:0]    writeBack_ENV_CTRL;
  wire       [1:0]    _zz_writeBack_ENV_CTRL;
  reg                 CsrPlugin_running_aheadValue;
  wire                decode_RS2_USE;
  wire                decode_RS1_USE;
  reg        [31:0]   _zz_decode_RS2;
  wire                execute_REGFILE_WRITE_VALID;
  wire                execute_BYPASSABLE_EXECUTE_STAGE;
  reg        [31:0]   _zz_decode_RS2_1;
  wire                memory_REGFILE_WRITE_VALID;
  wire                memory_BYPASSABLE_MEMORY_STAGE;
  wire                writeBack_REGFILE_WRITE_VALID;
  reg        [31:0]   decode_RS2;
  reg        [31:0]   decode_RS1;
  wire                execute_SRC_LESS_UNSIGNED;
  wire                execute_SRC2_FORCE_ZERO;
  wire       [31:0]   execute_SRC2;
  wire                execute_SRC_USE_SUB_LESS;
  wire       [31:0]   execute_SRC1;
  wire       [31:0]   _zz_decode_to_execute_PC;
  wire       [31:0]   _zz_decode_to_execute_RS2;
  wire       [1:0]    decode_SRC2_CTRL;
  wire       [1:0]    _zz_decode_SRC2_CTRL;
  wire       [31:0]   _zz_decode_to_execute_RS1;
  wire       [1:0]    decode_SRC1_CTRL;
  wire       [1:0]    _zz_decode_SRC1_CTRL;
  wire                decode_SRC_USE_SUB_LESS;
  wire                decode_SRC_ADD_ZERO;
  wire       [31:0]   _zz_lastStageRegFileWrite_payload_address;
  wire                _zz_lastStageRegFileWrite_valid;
  reg                 _zz_1;
  wire       [31:0]   decode_INSTRUCTION_ANTICIPATED;
  reg                 decode_REGFILE_WRITE_VALID;
  reg                 decode_LEGAL_INSTRUCTION;
  wire       [1:0]    _zz_decode_SHIFT_CTRL_1;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL_1;
  wire       [0:0]    _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1;
  wire       [0:0]    _zz_decode_FPU_FORMAT_1;
  wire       [3:0]    _zz_decode_FPU_OPCODE_1;
  wire                _zz_decode_FPU_ENABLE;
  wire       [1:0]    _zz_decode_BRANCH_CTRL_1;
  wire       [1:0]    _zz_decode_ENV_CTRL_1;
  wire       [1:0]    _zz_decode_SRC2_CTRL_1;
  wire       [1:0]    _zz_decode_ALU_CTRL_1;
  wire       [1:0]    _zz_decode_SRC1_CTRL_1;
  reg        [31:0]   _zz_decode_RS2_2;
  wire                writeBack_MEMORY_WR;
  wire                writeBack_MEMORY_FENCE;
  wire                writeBack_MEMORY_AMO;
  wire                writeBack_MEMORY_LRSC;
  wire       [31:0]   writeBack_MEMORY_STORE_DATA_RF;
  wire       [31:0]   writeBack_REGFILE_WRITE_DATA;
  wire                writeBack_MEMORY_ENABLE;
  wire       [31:0]   memory_PC;
  wire       [31:0]   memory_MEMORY_STORE_DATA_RF;
  wire       [31:0]   memory_REGFILE_WRITE_DATA;
  wire       [31:0]   memory_INSTRUCTION;
  wire                memory_MEMORY_WR;
  wire                memory_MEMORY_ENABLE;
  wire                execute_MEMORY_FENCE_WR;
  wire       [31:0]   memory_MEMORY_VIRTUAL_ADDRESS;
  wire                execute_MEMORY_AMO;
  wire                execute_MEMORY_LRSC;
  wire                execute_MEMORY_FORCE_CONSTISTENCY;
  (* keep , syn_keep *) wire       [31:0]   execute_RS1 /* synthesis syn_keep = 1 */ ;
  wire                execute_MEMORY_MANAGMENT;
  (* keep , syn_keep *) wire       [31:0]   execute_RS2 /* synthesis syn_keep = 1 */ ;
  wire                execute_MEMORY_WR;
  wire       [31:0]   execute_SRC_ADD;
  wire                execute_MEMORY_ENABLE;
  wire       [31:0]   execute_INSTRUCTION;
  wire                decode_MEMORY_AMO;
  wire                decode_MEMORY_LRSC;
  reg                 _zz_decode_MEMORY_FORCE_CONSTISTENCY;
  wire                decode_MEMORY_ENABLE;
  wire                decode_FLUSH_ALL;
  reg                 IBusCachedPlugin_rsp_issueDetected_4;
  reg                 IBusCachedPlugin_rsp_issueDetected_3;
  reg                 IBusCachedPlugin_rsp_issueDetected_2;
  reg                 IBusCachedPlugin_rsp_issueDetected_1;
  reg        [31:0]   _zz_memory_to_writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   decode_PC;
  wire       [31:0]   decode_INSTRUCTION;
  wire                decode_IS_RVC;
  wire       [31:0]   writeBack_PC;
  wire       [31:0]   writeBack_INSTRUCTION;
  reg                 decode_arbitration_haltItself;
  reg                 decode_arbitration_haltByOther;
  reg                 decode_arbitration_removeIt;
  wire                decode_arbitration_flushIt;
  reg                 decode_arbitration_flushNext;
  reg                 decode_arbitration_isValid;
  wire                decode_arbitration_isStuck;
  wire                decode_arbitration_isStuckByOthers;
  wire                decode_arbitration_isFlushed;
  wire                decode_arbitration_isMoving;
  wire                decode_arbitration_isFiring;
  reg                 execute_arbitration_haltItself;
  reg                 execute_arbitration_haltByOther;
  reg                 execute_arbitration_removeIt;
  wire                execute_arbitration_flushIt;
  reg                 execute_arbitration_flushNext;
  reg                 execute_arbitration_isValid;
  wire                execute_arbitration_isStuck;
  wire                execute_arbitration_isStuckByOthers;
  wire                execute_arbitration_isFlushed;
  wire                execute_arbitration_isMoving;
  wire                execute_arbitration_isFiring;
  reg                 memory_arbitration_haltItself;
  reg                 memory_arbitration_haltByOther;
  reg                 memory_arbitration_removeIt;
  wire                memory_arbitration_flushIt;
  reg                 memory_arbitration_flushNext;
  reg                 memory_arbitration_isValid;
  wire                memory_arbitration_isStuck;
  wire                memory_arbitration_isStuckByOthers;
  wire                memory_arbitration_isFlushed;
  wire                memory_arbitration_isMoving;
  wire                memory_arbitration_isFiring;
  reg                 writeBack_arbitration_haltItself;
  reg                 writeBack_arbitration_haltByOther;
  reg                 writeBack_arbitration_removeIt;
  reg                 writeBack_arbitration_flushIt;
  reg                 writeBack_arbitration_flushNext;
  reg                 writeBack_arbitration_isValid;
  wire                writeBack_arbitration_isStuck;
  wire                writeBack_arbitration_isStuckByOthers;
  wire                writeBack_arbitration_isFlushed;
  wire                writeBack_arbitration_isMoving;
  wire                writeBack_arbitration_isFiring;
  wire       [31:0]   lastStageInstruction /* verilator public */ ;
  wire       [31:0]   lastStagePc /* verilator public */ ;
  wire                lastStageIsValid /* verilator public */ ;
  wire                lastStageIsFiring /* verilator public */ ;
  reg                 IBusCachedPlugin_fetcherHalt;
  wire                IBusCachedPlugin_forceNoDecodeCond;
  reg                 IBusCachedPlugin_incomingInstruction;
  wire                IBusCachedPlugin_pcValids_0;
  wire                IBusCachedPlugin_pcValids_1;
  wire                IBusCachedPlugin_pcValids_2;
  wire                IBusCachedPlugin_pcValids_3;
  reg                 IBusCachedPlugin_decodeExceptionPort_valid;
  reg        [3:0]    IBusCachedPlugin_decodeExceptionPort_payload_code;
  wire       [31:0]   IBusCachedPlugin_decodeExceptionPort_payload_badAddr;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   IBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                IBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                IBusCachedPlugin_mmuBus_rsp_isPaging;
  wire                IBusCachedPlugin_mmuBus_rsp_allowRead;
  wire                IBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire                IBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                IBusCachedPlugin_mmuBus_rsp_exception;
  wire                IBusCachedPlugin_mmuBus_rsp_refilling;
  wire                IBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                IBusCachedPlugin_mmuBus_end;
  wire                IBusCachedPlugin_mmuBus_busy;
  wire                DBusCachedPlugin_trigger_valid;
  wire                DBusCachedPlugin_trigger_load;
  wire                DBusCachedPlugin_trigger_store;
  wire       [31:0]   DBusCachedPlugin_trigger_virtual;
  wire       [31:0]   DBusCachedPlugin_trigger_writeData;
  wire       [31:0]   DBusCachedPlugin_trigger_readData;
  wire                DBusCachedPlugin_trigger_readDataValid;
  wire       [1:0]    DBusCachedPlugin_trigger_size;
  wire       [31:0]   DBusCachedPlugin_trigger_dpc;
  wire                DBusCachedPlugin_trigger_hit;
  wire                DBusCachedPlugin_trigger_hitBefore;
  wire                DBusCachedPlugin_writesPending;
  wire                DBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                DBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   DBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   DBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                DBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                DBusCachedPlugin_mmuBus_rsp_isPaging;
  wire                DBusCachedPlugin_mmuBus_rsp_allowRead;
  wire                DBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire                DBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                DBusCachedPlugin_mmuBus_rsp_exception;
  wire                DBusCachedPlugin_mmuBus_rsp_refilling;
  wire                DBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                DBusCachedPlugin_mmuBus_end;
  wire                DBusCachedPlugin_mmuBus_busy;
  reg                 DBusCachedPlugin_redoBranch_valid;
  wire       [31:0]   DBusCachedPlugin_redoBranch_payload;
  reg                 DBusCachedPlugin_exceptionBus_valid;
  reg        [3:0]    DBusCachedPlugin_exceptionBus_payload_code;
  wire       [31:0]   DBusCachedPlugin_exceptionBus_payload_badAddr;
  wire                decodeExceptionPort_valid;
  wire       [3:0]    decodeExceptionPort_payload_code;
  wire       [31:0]   decodeExceptionPort_payload_badAddr;
  wire       [31:0]   CsrPlugin_csrMapping_readDataSignal;
  wire       [31:0]   CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   CsrPlugin_csrMapping_writeDataSignal;
  reg                 CsrPlugin_csrMapping_allowCsrSignal;
  wire                CsrPlugin_csrMapping_hazardFree;
  reg                 CsrPlugin_csrMapping_doForceFailCsr;
  wire                CsrPlugin_inWfi /* verilator public */ ;
  reg                 CsrPlugin_thirdPartyWake;
  reg                 CsrPlugin_jumpInterface_valid;
  reg        [31:0]   CsrPlugin_jumpInterface_payload;
  wire                CsrPlugin_exceptionPendings_0;
  wire                CsrPlugin_exceptionPendings_1;
  wire                CsrPlugin_exceptionPendings_2;
  wire                CsrPlugin_exceptionPendings_3;
  wire                contextSwitching;
  reg        [1:0]    CsrPlugin_privilege;
  wire                CsrPlugin_forceMachineWire;
  reg                 CsrPlugin_selfException_valid;
  reg        [3:0]    CsrPlugin_selfException_payload_code;
  wire       [31:0]   CsrPlugin_selfException_payload_badAddr;
  reg                 CsrPlugin_allowInterrupts;
  wire                CsrPlugin_allowException;
  wire                CsrPlugin_allowEbreakException;
  reg                 CsrPlugin_xretAwayFromMachine;
  wire                fpuAccess_start;
  wire       [4:0]    fpuAccess_regId;
  wire       [2:0]    fpuAccess_size;
  wire                fpuAccess_write;
  wire       [63:0]   fpuAccess_writeData;
  reg        [31:0]   fpuAccess_readData;
  reg                 fpuAccess_readDataValid;
  reg        [0:0]    fpuAccess_readDataChunk;
  reg                 fpuAccess_done;
  wire                CsrPlugin_injectionPort_valid;
  reg                 CsrPlugin_injectionPort_ready;
  wire       [31:0]   CsrPlugin_injectionPort_payload;
  wire                debugMode;
  wire                BranchPlugin_jumpInterface_valid;
  wire       [31:0]   BranchPlugin_jumpInterface_payload;
  reg                 BranchPlugin_inDebugNoFetchFlag;
  wire                IBusCachedPlugin_externalFlush;
  wire                IBusCachedPlugin_jump_pcLoad_valid;
  wire       [31:0]   IBusCachedPlugin_jump_pcLoad_payload;
  wire       [2:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload;
  wire       [2:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  wire                _zz_IBusCachedPlugin_jump_pcLoad_payload_2;
  wire                _zz_IBusCachedPlugin_jump_pcLoad_payload_3;
  wire                IBusCachedPlugin_fetchPc_output_valid;
  wire                IBusCachedPlugin_fetchPc_output_ready;
  wire       [31:0]   IBusCachedPlugin_fetchPc_output_payload;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pcReg /* verilator public */ ;
  reg                 IBusCachedPlugin_fetchPc_correction;
  reg                 IBusCachedPlugin_fetchPc_correctionReg;
  wire                IBusCachedPlugin_fetchPc_output_fire;
  wire                IBusCachedPlugin_fetchPc_corrected;
  reg                 IBusCachedPlugin_fetchPc_pcRegPropagate;
  reg                 IBusCachedPlugin_fetchPc_booted;
  reg                 IBusCachedPlugin_fetchPc_inc;
  wire                when_Fetcher_l133;
  wire                when_Fetcher_l133_1;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pc;
  wire                IBusCachedPlugin_fetchPc_redo_valid;
  reg        [31:0]   IBusCachedPlugin_fetchPc_redo_payload;
  reg                 IBusCachedPlugin_fetchPc_flushed;
  wire                when_Fetcher_l160;
  reg                 IBusCachedPlugin_decodePc_flushed;
  reg        [31:0]   IBusCachedPlugin_decodePc_pcReg /* verilator public */ ;
  wire       [31:0]   IBusCachedPlugin_decodePc_pcPlus;
  reg                 IBusCachedPlugin_decodePc_injectedDecode;
  wire                when_Fetcher_l182;
  wire                when_Fetcher_l194;
  reg                 IBusCachedPlugin_iBusRsp_redoFetch;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_0_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_1_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_2_halt;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire                IBusCachedPlugin_iBusRsp_flush;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  reg        [31:0]   _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 IBusCachedPlugin_iBusRsp_readyForError;
  wire                IBusCachedPlugin_iBusRsp_output_valid;
  wire                IBusCachedPlugin_iBusRsp_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_pc;
  wire                IBusCachedPlugin_iBusRsp_output_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  wire                IBusCachedPlugin_iBusRsp_output_payload_isRvc;
  wire                when_Fetcher_l242;
  wire                IBusCachedPlugin_decompressor_input_valid;
  wire                IBusCachedPlugin_decompressor_input_ready;
  wire       [31:0]   IBusCachedPlugin_decompressor_input_payload_pc;
  wire                IBusCachedPlugin_decompressor_input_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_decompressor_input_payload_rsp_inst;
  wire                IBusCachedPlugin_decompressor_input_payload_isRvc;
  wire                IBusCachedPlugin_decompressor_output_valid;
  wire                IBusCachedPlugin_decompressor_output_ready;
  wire       [31:0]   IBusCachedPlugin_decompressor_output_payload_pc;
  wire                IBusCachedPlugin_decompressor_output_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_decompressor_output_payload_rsp_inst;
  wire                IBusCachedPlugin_decompressor_output_payload_isRvc;
  wire                IBusCachedPlugin_decompressor_flushNext;
  wire                IBusCachedPlugin_decompressor_consumeCurrent;
  reg                 IBusCachedPlugin_decompressor_bufferValid;
  reg        [15:0]   IBusCachedPlugin_decompressor_bufferData;
  wire                IBusCachedPlugin_decompressor_isInputLowRvc;
  wire                IBusCachedPlugin_decompressor_isInputHighRvc;
  reg                 IBusCachedPlugin_decompressor_throw2BytesReg;
  wire                IBusCachedPlugin_decompressor_throw2Bytes;
  wire                IBusCachedPlugin_decompressor_unaligned;
  reg                 IBusCachedPlugin_decompressor_bufferValidLatch;
  reg                 IBusCachedPlugin_decompressor_throw2BytesLatch;
  wire                IBusCachedPlugin_decompressor_bufferValidPatched;
  wire                IBusCachedPlugin_decompressor_throw2BytesPatched;
  wire       [31:0]   IBusCachedPlugin_decompressor_raw;
  wire                IBusCachedPlugin_decompressor_isRvc;
  wire       [15:0]   _zz_IBusCachedPlugin_decompressor_decompressed;
  reg        [31:0]   IBusCachedPlugin_decompressor_decompressed;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_1;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_2;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_3;
  wire       [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_4;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_5;
  reg        [11:0]   _zz_IBusCachedPlugin_decompressor_decompressed_6;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_7;
  reg        [9:0]    _zz_IBusCachedPlugin_decompressor_decompressed_8;
  wire       [20:0]   _zz_IBusCachedPlugin_decompressor_decompressed_9;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_10;
  reg        [14:0]   _zz_IBusCachedPlugin_decompressor_decompressed_11;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_12;
  reg        [2:0]    _zz_IBusCachedPlugin_decompressor_decompressed_13;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_14;
  reg        [9:0]    _zz_IBusCachedPlugin_decompressor_decompressed_15;
  wire       [20:0]   _zz_IBusCachedPlugin_decompressor_decompressed_16;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_17;
  reg        [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_18;
  wire       [12:0]   _zz_IBusCachedPlugin_decompressor_decompressed_19;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_20;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_21;
  wire       [4:0]    _zz_IBusCachedPlugin_decompressor_decompressed_22;
  wire       [4:0]    switch_Misc_l44;
  wire                when_Misc_l47;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_23;
  wire       [1:0]    switch_Misc_l241;
  wire       [1:0]    switch_Misc_l241_1;
  reg        [2:0]    _zz_IBusCachedPlugin_decompressor_decompressed_24;
  reg        [2:0]    _zz_IBusCachedPlugin_decompressor_decompressed_25;
  wire                _zz_IBusCachedPlugin_decompressor_decompressed_26;
  reg        [6:0]    _zz_IBusCachedPlugin_decompressor_decompressed_27;
  wire                IBusCachedPlugin_decompressor_output_fire;
  wire                IBusCachedPlugin_decompressor_bufferFill;
  wire                when_Fetcher_l285;
  wire                when_Fetcher_l288;
  wire                when_Fetcher_l293;
  wire                IBusCachedPlugin_injector_decodeInput_valid;
  wire                IBusCachedPlugin_injector_decodeInput_ready;
  wire       [31:0]   IBusCachedPlugin_injector_decodeInput_payload_pc;
  wire                IBusCachedPlugin_injector_decodeInput_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  wire                IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  reg                 _zz_IBusCachedPlugin_injector_decodeInput_valid;
  reg        [31:0]   _zz_IBusCachedPlugin_injector_decodeInput_payload_pc;
  reg                 _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_error;
  reg        [31:0]   _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  reg                 _zz_IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_0;
  wire                when_Fetcher_l331;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_1;
  wire                when_Fetcher_l331_1;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_2;
  wire                when_Fetcher_l331_2;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_3;
  wire                when_Fetcher_l331_3;
  reg        [31:0]   IBusCachedPlugin_injector_formal_rawInDecode;
  reg        [31:0]   IBusCachedPlugin_rspCounter;
  wire                IBusCachedPlugin_s0_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s1_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s2_tightlyCoupledHit;
  wire                IBusCachedPlugin_rsp_iBusRspOutputHalt;
  wire                IBusCachedPlugin_rsp_issueDetected;
  reg                 IBusCachedPlugin_rsp_redoFetch;
  wire                when_IBusCachedPlugin_l245;
  wire                when_IBusCachedPlugin_l250;
  wire                when_IBusCachedPlugin_l256;
  wire                when_IBusCachedPlugin_l262;
  wire                when_IBusCachedPlugin_l273;
  wire                dataCache_2_io_mem_cmd_s2mPipe_valid;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_ready;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_wr;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_uncached;
  wire       [31:0]   dataCache_2_io_mem_cmd_s2mPipe_payload_address;
  wire       [63:0]   dataCache_2_io_mem_cmd_s2mPipe_payload_data;
  wire       [7:0]    dataCache_2_io_mem_cmd_s2mPipe_payload_mask;
  wire       [2:0]    dataCache_2_io_mem_cmd_s2mPipe_payload_size;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_exclusive;
  wire                dataCache_2_io_mem_cmd_s2mPipe_payload_last;
  reg                 dataCache_2_io_mem_cmd_rValidN;
  reg                 dataCache_2_io_mem_cmd_rData_wr;
  reg                 dataCache_2_io_mem_cmd_rData_uncached;
  reg        [31:0]   dataCache_2_io_mem_cmd_rData_address;
  reg        [63:0]   dataCache_2_io_mem_cmd_rData_data;
  reg        [7:0]    dataCache_2_io_mem_cmd_rData_mask;
  reg        [2:0]    dataCache_2_io_mem_cmd_rData_size;
  reg                 dataCache_2_io_mem_cmd_rData_exclusive;
  reg                 dataCache_2_io_mem_cmd_rData_last;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_ready;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_wr;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached;
  wire       [31:0]   dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_address;
  wire       [63:0]   dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_data;
  wire       [7:0]    dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_mask;
  wire       [2:0]    dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_size;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_exclusive;
  wire                dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_last;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rValid;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_wr;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_uncached;
  reg        [31:0]   dataCache_2_io_mem_cmd_s2mPipe_rData_address;
  reg        [63:0]   dataCache_2_io_mem_cmd_s2mPipe_rData_data;
  reg        [7:0]    dataCache_2_io_mem_cmd_s2mPipe_rData_mask;
  reg        [2:0]    dataCache_2_io_mem_cmd_s2mPipe_rData_size;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_exclusive;
  reg                 dataCache_2_io_mem_cmd_s2mPipe_rData_last;
  wire                when_Stream_l375;
  reg                 dBus_rsp_valid_regNext;
  reg                 dBus_rsp_payload_exclusive_regNext;
  reg                 dBus_rsp_payload_error_regNext;
  reg                 dBus_rsp_payload_last_regNext;
  reg        [3:0]    dBus_rsp_payload_aggregated_regNext;
  wire                when_DBusCachedPlugin_l334;
  reg        [63:0]   dBus_rsp_payload_data_regNextWhen;
  reg        [31:0]   DBusCachedPlugin_rspCounter;
  wire                when_DBusCachedPlugin_l356;
  wire                when_DBusCachedPlugin_l364;
  wire       [1:0]    execute_DBusCachedPlugin_size;
  reg        [31:0]   _zz_execute_MEMORY_STORE_DATA_RF;
  wire                dataCache_2_io_cpu_flush_isStall;
  wire                when_DBusCachedPlugin_l398;
  wire                when_DBusCachedPlugin_l414;
  wire                when_DBusCachedPlugin_l427;
  wire                when_DBusCachedPlugin_l476;
  wire       [11:0]   _zz_io_cpu_writeBack_fence_SW;
  reg                 writeBack_DBusCachedPlugin_fence_aquire;
  wire                when_DBusCachedPlugin_l518;
  wire                when_DBusCachedPlugin_l531;
  wire                when_DBusCachedPlugin_l535;
  wire                when_DBusCachedPlugin_l552;
  wire                when_DBusCachedPlugin_l572;
  wire       [63:0]   writeBack_DBusCachedPlugin_rspData;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_0;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_1;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_2;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_3;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_4;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_5;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_6;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_7;
  reg        [63:0]   writeBack_DBusCachedPlugin_rspShifted;
  reg        [31:0]   writeBack_DBusCachedPlugin_rspRf;
  wire                when_DBusCachedPlugin_l589;
  wire       [1:0]    switch_Misc_l241_2;
  wire                _zz_writeBack_DBusCachedPlugin_rspFormated;
  reg        [31:0]   _zz_writeBack_DBusCachedPlugin_rspFormated_1;
  wire                _zz_writeBack_DBusCachedPlugin_rspFormated_2;
  reg        [31:0]   _zz_writeBack_DBusCachedPlugin_rspFormated_3;
  reg        [31:0]   writeBack_DBusCachedPlugin_rspFormated;
  wire                when_DBusCachedPlugin_l599;
  wire       [47:0]   _zz_decode_CfuPlugin_CFU_ENABLE;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_1;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_2;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_3;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_4;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_5;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_6;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_7;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_8;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_9;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_10;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_11;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_12;
  wire                _zz_decode_CfuPlugin_CFU_ENABLE_13;
  wire       [1:0]    _zz_decode_SRC1_CTRL_2;
  wire       [1:0]    _zz_decode_ALU_CTRL_2;
  wire       [1:0]    _zz_decode_SRC2_CTRL_2;
  wire       [1:0]    _zz_decode_ENV_CTRL_2;
  wire       [1:0]    _zz_decode_BRANCH_CTRL_2;
  wire       [3:0]    _zz_decode_FPU_OPCODE_2;
  wire       [0:0]    _zz_decode_FPU_FORMAT_2;
  wire       [0:0]    _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL_2;
  wire       [1:0]    _zz_decode_SHIFT_CTRL_2;
  wire                when_RegFilePlugin_l63;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress1;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress2;
  wire       [31:0]   decode_RegFilePlugin_rs1Data;
  wire       [31:0]   decode_RegFilePlugin_rs2Data;
  reg                 lastStageRegFileWrite_valid /* verilator public */ ;
  reg        [4:0]    lastStageRegFileWrite_payload_address /* verilator public */ ;
  reg        [31:0]   lastStageRegFileWrite_payload_data /* verilator public */ ;
  reg                 _zz_5;
  reg        [31:0]   _zz_decode_SRC1;
  wire                _zz_decode_SRC2;
  reg        [19:0]   _zz_decode_SRC2_1;
  wire                _zz_decode_SRC2_2;
  reg        [19:0]   _zz_decode_SRC2_3;
  reg        [31:0]   _zz_decode_SRC2_4;
  reg        [31:0]   execute_SrcPlugin_addSub;
  wire                execute_SrcPlugin_less;
  reg                 HazardSimplePlugin_src0Hazard;
  reg                 HazardSimplePlugin_src1Hazard;
  wire                HazardSimplePlugin_writeBackWrites_valid;
  wire       [4:0]    HazardSimplePlugin_writeBackWrites_payload_address;
  wire       [31:0]   HazardSimplePlugin_writeBackWrites_payload_data;
  reg                 HazardSimplePlugin_writeBackBuffer_valid;
  reg        [4:0]    HazardSimplePlugin_writeBackBuffer_payload_address;
  reg        [31:0]   HazardSimplePlugin_writeBackBuffer_payload_data;
  wire                HazardSimplePlugin_addr0Match;
  wire                HazardSimplePlugin_addr1Match;
  wire                when_HazardSimplePlugin_l47;
  wire                when_HazardSimplePlugin_l48;
  wire                when_HazardSimplePlugin_l51;
  wire                when_HazardSimplePlugin_l45;
  wire                when_HazardSimplePlugin_l57;
  wire                when_HazardSimplePlugin_l58;
  wire                when_HazardSimplePlugin_l48_1;
  wire                when_HazardSimplePlugin_l51_1;
  wire                when_HazardSimplePlugin_l45_1;
  wire                when_HazardSimplePlugin_l57_1;
  wire                when_HazardSimplePlugin_l58_1;
  wire                when_HazardSimplePlugin_l48_2;
  wire                when_HazardSimplePlugin_l51_2;
  wire                when_HazardSimplePlugin_l45_2;
  wire                when_HazardSimplePlugin_l57_2;
  wire                when_HazardSimplePlugin_l58_2;
  wire                when_HazardSimplePlugin_l105;
  wire                when_HazardSimplePlugin_l108;
  wire                when_HazardSimplePlugin_l113;
  reg                 when_CsrPlugin_l836;
  reg        [1:0]    _zz_CsrPlugin_privilege;
  reg                 CsrPlugin_running;
  wire                when_CsrPlugin_l729;
  reg                 CsrPlugin_reseting;
  reg                 _zz_debugBus_haveReset;
  reg                 CsrPlugin_running_aheadValue_regNext;
  wire                CsrPlugin_enterHalt;
  reg                 CsrPlugin_doHalt;
  wire                when_CsrPlugin_l747;
  wire                CsrPlugin_forceResume;
  reg                 _zz_CsrPlugin_doResume;
  wire                CsrPlugin_doResume;
  reg                 CsrPlugin_timeout_state;
  reg                 CsrPlugin_timeout_stateRise;
  wire                CsrPlugin_timeout_counter_willIncrement;
  reg                 CsrPlugin_timeout_counter_willClear;
  reg        [2:0]    CsrPlugin_timeout_counter_valueNext;
  reg        [2:0]    CsrPlugin_timeout_counter_value;
  wire                CsrPlugin_timeout_counter_willOverflowIfInc;
  wire                CsrPlugin_timeout_counter_willOverflow;
  wire                when_CsrPlugin_l753;
  reg                 _zz_debugBus_hartToDm_valid;
  reg        [31:0]   CsrPlugin_dataCsrw_value_0;
  reg        [31:0]   CsrPlugin_dataCsrw_value_1;
  wire                when_CsrPlugin_l768;
  wire       [1:0]    _zz_6;
  wire                CsrPlugin_inject_cmd_valid;
  wire       [1:0]    CsrPlugin_inject_cmd_payload_op;
  wire       [4:0]    CsrPlugin_inject_cmd_payload_address;
  wire       [31:0]   CsrPlugin_inject_cmd_payload_data;
  wire       [2:0]    CsrPlugin_inject_cmd_payload_size;
  wire                CsrPlugin_inject_cmd_toStream_valid;
  reg                 CsrPlugin_inject_cmd_toStream_ready;
  wire       [1:0]    CsrPlugin_inject_cmd_toStream_payload_op;
  wire       [4:0]    CsrPlugin_inject_cmd_toStream_payload_address;
  wire       [31:0]   CsrPlugin_inject_cmd_toStream_payload_data;
  wire       [2:0]    CsrPlugin_inject_cmd_toStream_payload_size;
  wire                CsrPlugin_inject_buffer_valid;
  reg                 CsrPlugin_inject_buffer_ready;
  wire       [1:0]    CsrPlugin_inject_buffer_payload_op;
  wire       [4:0]    CsrPlugin_inject_buffer_payload_address;
  wire       [31:0]   CsrPlugin_inject_buffer_payload_data;
  wire       [2:0]    CsrPlugin_inject_buffer_payload_size;
  reg                 CsrPlugin_inject_cmd_toStream_rValid;
  reg        [1:0]    CsrPlugin_inject_cmd_toStream_rData_op;
  reg        [4:0]    CsrPlugin_inject_cmd_toStream_rData_address;
  reg        [31:0]   CsrPlugin_inject_cmd_toStream_rData_data;
  reg        [2:0]    CsrPlugin_inject_cmd_toStream_rData_size;
  wire                when_Stream_l375_1;
  wire                CsrPlugin_injectionPort_fire;
  reg                 CsrPlugin_inject_pending;
  wire                when_CsrPlugin_l804;
  wire                when_CsrPlugin_l804_1;
  reg        [31:0]   CsrPlugin_dpc;
  reg        [1:0]    CsrPlugin_dcsr_prv;
  reg                 CsrPlugin_dcsr_step;
  wire                CsrPlugin_dcsr_nmip;
  wire                CsrPlugin_dcsr_mprven;
  reg        [2:0]    CsrPlugin_dcsr_cause;
  reg                 CsrPlugin_dcsr_stoptime;
  reg                 CsrPlugin_dcsr_stopcount;
  reg                 CsrPlugin_dcsr_stepie;
  reg                 CsrPlugin_dcsr_ebreakm;
  wire       [3:0]    CsrPlugin_dcsr_xdebugver;
  wire                CsrPlugin_dcsr_stepLogic_wantExit;
  reg                 CsrPlugin_dcsr_stepLogic_wantStart;
  wire                CsrPlugin_dcsr_stepLogic_wantKill;
  reg        [1:0]    CsrPlugin_dcsr_stepLogic_stateReg;
  reg        [1:0]    CsrPlugin_dcsr_stepLogic_stateNext;
  wire                when_CsrPlugin_l830;
  wire                when_CsrPlugin_l848;
  wire                when_CsrPlugin_l880;
  wire       [1:0]    CsrPlugin_misa_base;
  wire       [25:0]   CsrPlugin_misa_extensions;
  reg        [1:0]    CsrPlugin_mtvec_mode;
  reg        [29:0]   CsrPlugin_mtvec_base;
  reg        [31:0]   CsrPlugin_mepc;
  reg                 CsrPlugin_mstatus_MIE;
  reg                 CsrPlugin_mstatus_MPIE;
  reg        [1:0]    CsrPlugin_mstatus_MPP;
  reg                 CsrPlugin_mip_MEIP;
  reg                 CsrPlugin_mip_MTIP;
  reg                 CsrPlugin_mip_MSIP;
  reg                 CsrPlugin_mie_MEIE;
  reg                 CsrPlugin_mie_MTIE;
  reg                 CsrPlugin_mie_MSIE;
  reg        [31:0]   CsrPlugin_mscratch;
  reg                 CsrPlugin_mcause_interrupt;
  reg        [3:0]    CsrPlugin_mcause_exceptionCode;
  reg        [31:0]   CsrPlugin_mtval;
  reg        [63:0]   CsrPlugin_counters_mcycle;
  reg        [63:0]   CsrPlugin_counters_minstret;
  wire                _zz_when_CsrPlugin_l1446;
  wire                _zz_when_CsrPlugin_l1446_1;
  wire                _zz_when_CsrPlugin_l1446_2;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  reg        [3:0]    CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  reg        [31:0]   CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
  wire       [1:0]    _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  wire                _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire                when_CsrPlugin_l1403;
  wire                when_CsrPlugin_l1403_1;
  wire                when_CsrPlugin_l1403_2;
  wire                when_CsrPlugin_l1403_3;
  wire                when_CsrPlugin_l1416;
  reg                 CsrPlugin_interrupt_valid;
  reg        [3:0]    CsrPlugin_interrupt_code /* verilator public */ ;
  reg        [1:0]    CsrPlugin_interrupt_targetPrivilege;
  wire                when_CsrPlugin_l1440;
  wire                when_CsrPlugin_l1446;
  wire                when_CsrPlugin_l1446_1;
  wire                when_CsrPlugin_l1446_2;
  wire                when_CsrPlugin_l1459;
  wire                CsrPlugin_exception;
  wire                CsrPlugin_lastStageWasWfi;
  reg                 CsrPlugin_pipelineLiberator_pcValids_0;
  reg                 CsrPlugin_pipelineLiberator_pcValids_1;
  reg                 CsrPlugin_pipelineLiberator_pcValids_2;
  wire                CsrPlugin_pipelineLiberator_active;
  wire                when_CsrPlugin_l1479;
  wire                when_CsrPlugin_l1479_1;
  wire                when_CsrPlugin_l1479_2;
  wire                when_CsrPlugin_l1484;
  reg                 CsrPlugin_pipelineLiberator_done;
  wire                when_CsrPlugin_l1490;
  wire                CsrPlugin_interruptJump /* verilator public */ ;
  reg                 CsrPlugin_hadException /* verilator public */ ;
  reg        [1:0]    CsrPlugin_targetPrivilege;
  reg        [3:0]    CsrPlugin_trapCause;
  reg                 CsrPlugin_trapCauseEbreakDebug;
  wire                when_CsrPlugin_l1517;
  wire                when_CsrPlugin_l1519;
  reg        [1:0]    CsrPlugin_xtvec_mode;
  reg        [29:0]   CsrPlugin_xtvec_base;
  reg                 CsrPlugin_trapEnterDebug;
  wire                when_CsrPlugin_l1533;
  wire                when_CsrPlugin_l1534;
  wire                when_CsrPlugin_l1542;
  wire                when_CsrPlugin_l1572;
  wire                when_CsrPlugin_l1600;
  wire       [1:0]    switch_CsrPlugin_l1604;
  wire                when_CsrPlugin_l1612;
  reg                 execute_CsrPlugin_wfiWake;
  wire                when_CsrPlugin_l1671;
  wire                execute_CsrPlugin_blockedBySideEffects;
  reg                 execute_CsrPlugin_illegalAccess;
  reg                 execute_CsrPlugin_illegalInstruction;
  wire                when_CsrPlugin_l1684;
  wire                when_CsrPlugin_l1691;
  wire                when_CsrPlugin_l1692;
  wire                when_CsrPlugin_l1699;
  wire                when_CsrPlugin_l1709;
  reg                 execute_CsrPlugin_writeInstruction;
  reg                 execute_CsrPlugin_readInstruction;
  wire                execute_CsrPlugin_writeEnable;
  wire                execute_CsrPlugin_readEnable;
  wire       [31:0]   execute_CsrPlugin_readToWriteData;
  wire                switch_Misc_l241_3;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_writeDataSignal;
  wire                when_CsrPlugin_l1731;
  wire                when_CsrPlugin_l1735;
  wire       [11:0]   execute_CsrPlugin_csrAddress;
  wire                execute_BranchPlugin_eq;
  wire       [2:0]    switch_Misc_l241_4;
  reg                 _zz_execute_BRANCH_DO;
  reg                 _zz_execute_BRANCH_DO_1;
  wire       [31:0]   execute_BranchPlugin_branch_src1;
  wire                _zz_execute_BranchPlugin_branch_src2;
  reg        [10:0]   _zz_execute_BranchPlugin_branch_src2_1;
  wire                _zz_execute_BranchPlugin_branch_src2_2;
  reg        [19:0]   _zz_execute_BranchPlugin_branch_src2_3;
  wire                _zz_execute_BranchPlugin_branch_src2_4;
  reg        [18:0]   _zz_execute_BranchPlugin_branch_src2_5;
  reg        [31:0]   _zz_execute_BranchPlugin_branch_src2_6;
  wire       [31:0]   execute_BranchPlugin_branch_src2;
  wire       [31:0]   execute_BranchPlugin_branchAdder;
  reg                 execute_MulPlugin_aSigned;
  reg                 execute_MulPlugin_bSigned;
  wire       [31:0]   execute_MulPlugin_a;
  wire       [31:0]   execute_MulPlugin_b;
  reg        [0:0]    execute_MulPlugin_delayLogic_counter;
  wire                when_MulPlugin_l65;
  wire                when_MulPlugin_l70;
  wire       [1:0]    switch_MulPlugin_l87;
  wire       [15:0]   execute_MulPlugin_aULow;
  wire       [15:0]   execute_MulPlugin_bULow;
  wire       [16:0]   execute_MulPlugin_aSLow;
  wire       [16:0]   execute_MulPlugin_bSLow;
  wire       [16:0]   execute_MulPlugin_aHigh;
  wire       [16:0]   execute_MulPlugin_bHigh;
  reg        [31:0]   execute_MulPlugin_withOuputBuffer_mul_ll;
  reg        [33:0]   execute_MulPlugin_withOuputBuffer_mul_lh;
  reg        [33:0]   execute_MulPlugin_withOuputBuffer_mul_hl;
  reg        [33:0]   execute_MulPlugin_withOuputBuffer_mul_hh;
  wire       [65:0]   writeBack_MulPlugin_result;
  wire                when_MulPlugin_l147;
  wire       [1:0]    switch_MulPlugin_l148;
  reg        [32:0]   memory_MulDivIterativePlugin_rs1;
  reg        [31:0]   memory_MulDivIterativePlugin_rs2;
  reg        [64:0]   memory_MulDivIterativePlugin_accumulator;
  wire                memory_MulDivIterativePlugin_frontendOk;
  reg                 memory_MulDivIterativePlugin_div_needRevert;
  reg                 memory_MulDivIterativePlugin_div_counter_willIncrement;
  reg                 memory_MulDivIterativePlugin_div_counter_willClear;
  reg        [5:0]    memory_MulDivIterativePlugin_div_counter_valueNext;
  reg        [5:0]    memory_MulDivIterativePlugin_div_counter_value;
  wire                memory_MulDivIterativePlugin_div_counter_willOverflowIfInc;
  wire                memory_MulDivIterativePlugin_div_counter_willOverflow;
  reg                 memory_MulDivIterativePlugin_div_done;
  wire                when_MulDivIterativePlugin_l126;
  wire                when_MulDivIterativePlugin_l126_1;
  reg        [31:0]   memory_MulDivIterativePlugin_div_result;
  wire                when_MulDivIterativePlugin_l128;
  wire                when_MulDivIterativePlugin_l129;
  wire                when_MulDivIterativePlugin_l132;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted;
  wire       [32:0]   memory_MulDivIterativePlugin_div_stage_0_remainderShifted;
  wire       [32:0]   memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator;
  wire       [31:0]   memory_MulDivIterativePlugin_div_stage_0_outRemainder;
  wire       [31:0]   memory_MulDivIterativePlugin_div_stage_0_outNumerator;
  wire                when_MulDivIterativePlugin_l151;
  wire       [31:0]   _zz_memory_MulDivIterativePlugin_div_result;
  wire                when_MulDivIterativePlugin_l162;
  wire                _zz_memory_MulDivIterativePlugin_rs2;
  wire                _zz_memory_MulDivIterativePlugin_rs1;
  reg        [32:0]   _zz_memory_MulDivIterativePlugin_rs1_1;
  reg        [5:0]    FpuPlugin_pendings;
  wire                FpuPlugin_port_cmd_fire;
  wire                FpuPlugin_port_rsp_fire;
  wire                FpuPlugin_hasPending;
  reg                 FpuPlugin_flags_NX;
  reg                 FpuPlugin_flags_UF;
  reg                 FpuPlugin_flags_OF;
  reg                 FpuPlugin_flags_DZ;
  reg                 FpuPlugin_flags_NV;
  wire                when_FpuPlugin_l215;
  wire                when_FpuPlugin_l216;
  wire                when_FpuPlugin_l217;
  wire                when_FpuPlugin_l218;
  wire                when_FpuPlugin_l219;
  reg        [2:0]    FpuPlugin_rm;
  wire                FpuPlugin_csrActive;
  wire                when_FpuPlugin_l229;
  reg        [1:0]    FpuPlugin_fs;
  wire                FpuPlugin_sd;
  wire                when_FpuPlugin_l234;
  reg                 _zz_when_FpuPlugin_l237;
  reg                 _zz_when_FpuPlugin_l237_1;
  reg                 _zz_when_FpuPlugin_l237_2;
  wire                when_FpuPlugin_l237;
  reg                 FpuPlugin_accessFpuCsr;
  wire                when_FpuPlugin_l253;
  reg                 _zz_decode_FPU_FORKED;
  wire                decode_FpuPlugin_trap;
  reg                 decode_FpuPlugin_forked;
  wire                when_FpuPlugin_l268;
  wire                when_FpuPlugin_l268_1;
  wire                decode_FpuPlugin_hazard;
  wire                when_FpuPlugin_l272;
  wire                when_FpuPlugin_l273;
  wire                FpuPlugin_port_cmd_isStall;
  wire       [2:0]    decode_FpuPlugin_iRoundMode;
  wire       [2:0]    decode_FpuPlugin_roundMode;
  wire       [2:0]    _zz_FpuPlugin_port_cmd_payload_roundMode;
  wire       [2:0]    _zz_FpuPlugin_port_cmd_payload_roundMode_1;
  wire                writeBack_FpuPlugin_isRsp;
  wire                writeBack_FpuPlugin_isCommit;
  reg        [63:0]   writeBack_FpuPlugin_storeFormated;
  wire                when_FpuPlugin_l306;
  wire       [63:0]   DBusBypass0_value;
  wire                when_FpuPlugin_l315;
  wire                when_FpuPlugin_l318;
  wire                when_FpuPlugin_l323;
  wire                when_FpuPlugin_l325;
  wire                writeBack_FpuPlugin_commit_valid /* verilator public */ ;
  wire                writeBack_FpuPlugin_commit_ready /* verilator public */ ;
  wire       [3:0]    writeBack_FpuPlugin_commit_payload_opcode /* verilator public */ ;
  wire       [4:0]    writeBack_FpuPlugin_commit_payload_rd /* verilator public */ ;
  wire                writeBack_FpuPlugin_commit_payload_write /* verilator public */ ;
  reg        [63:0]   writeBack_FpuPlugin_commit_payload_value /* verilator public */ ;
  wire                when_FpuPlugin_l339;
  wire                writeBack_FpuPlugin_commit_s2mPipe_valid;
  wire                writeBack_FpuPlugin_commit_s2mPipe_ready;
  wire       [3:0]    writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
  wire       [4:0]    writeBack_FpuPlugin_commit_s2mPipe_payload_rd;
  wire                writeBack_FpuPlugin_commit_s2mPipe_payload_write;
  wire       [63:0]   writeBack_FpuPlugin_commit_s2mPipe_payload_value;
  reg                 writeBack_FpuPlugin_commit_rValidN;
  reg        [3:0]    writeBack_FpuPlugin_commit_rData_opcode;
  reg        [4:0]    writeBack_FpuPlugin_commit_rData_rd;
  reg                 writeBack_FpuPlugin_commit_rData_write;
  reg        [63:0]   writeBack_FpuPlugin_commit_rData_value;
  wire       [3:0]    _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
  wire                FpuPlugin_wantExit;
  reg                 FpuPlugin_wantStart;
  wire                FpuPlugin_wantKill;
  wire                when_FpuPlugin_l350;
  wire                when_CfuPlugin_l192;
  wire                execute_CfuPlugin_hazard;
  wire                execute_CfuPlugin_scheduleWish;
  wire                execute_CfuPlugin_schedule;
  wire                when_CfuPlugin_l196;
  reg                 execute_CfuPlugin_hold;
  reg                 execute_CfuPlugin_fired;
  wire                CfuPlugin_bus_cmd_fire;
  wire                when_CfuPlugin_l199;
  wire                when_CfuPlugin_l203;
  wire       [9:0]    execute_CfuPlugin_functionsIds_0;
  wire                _zz_CfuPlugin_bus_cmd_payload_inputs_1;
  reg        [23:0]   _zz_CfuPlugin_bus_cmd_payload_inputs_1_1;
  reg        [31:0]   _zz_CfuPlugin_bus_cmd_payload_inputs_1_2;
  wire                writeBack_CfuPlugin_rsp_valid;
  reg                 writeBack_CfuPlugin_rsp_ready;
  wire       [31:0]   writeBack_CfuPlugin_rsp_payload_outputs_0;
  reg                 CfuPlugin_bus_rsp_rValidN;
  reg        [31:0]   CfuPlugin_bus_rsp_rData_outputs_0;
  wire                when_CfuPlugin_l239;
  reg        [31:0]   _zz_decode_RS2_3;
  wire                when_Pipeline_l124;
  reg        [31:0]   decode_to_execute_PC;
  wire                when_Pipeline_l124_1;
  reg        [31:0]   execute_to_memory_PC;
  wire                when_Pipeline_l124_2;
  reg        [31:0]   memory_to_writeBack_PC;
  wire                when_Pipeline_l124_3;
  reg        [31:0]   decode_to_execute_INSTRUCTION;
  wire                when_Pipeline_l124_4;
  reg        [31:0]   execute_to_memory_INSTRUCTION;
  wire                when_Pipeline_l124_5;
  reg        [31:0]   memory_to_writeBack_INSTRUCTION;
  wire                when_Pipeline_l124_6;
  reg        [31:0]   decode_to_execute_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_7;
  reg        [31:0]   execute_to_memory_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_8;
  reg        [31:0]   memory_to_writeBack_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_9;
  reg                 decode_to_execute_MEMORY_FORCE_CONSTISTENCY;
  wire                when_Pipeline_l124_10;
  reg                 decode_to_execute_LEGAL_INSTRUCTION;
  wire                when_Pipeline_l124_11;
  reg                 decode_to_execute_MEMORY_FENCE_WR;
  wire                when_Pipeline_l124_12;
  reg                 decode_to_execute_SRC_USE_SUB_LESS;
  wire                when_Pipeline_l124_13;
  reg                 decode_to_execute_MEMORY_ENABLE;
  wire                when_Pipeline_l124_14;
  reg                 execute_to_memory_MEMORY_ENABLE;
  wire                when_Pipeline_l124_15;
  reg                 memory_to_writeBack_MEMORY_ENABLE;
  wire                when_Pipeline_l124_16;
  reg        [1:0]    decode_to_execute_ALU_CTRL;
  wire                when_Pipeline_l124_17;
  reg                 decode_to_execute_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_18;
  reg                 execute_to_memory_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_19;
  reg                 memory_to_writeBack_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_20;
  reg                 decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  wire                when_Pipeline_l124_21;
  reg                 decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_22;
  reg                 execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_23;
  reg                 decode_to_execute_MEMORY_WR;
  wire                when_Pipeline_l124_24;
  reg                 execute_to_memory_MEMORY_WR;
  wire                when_Pipeline_l124_25;
  reg                 memory_to_writeBack_MEMORY_WR;
  wire                when_Pipeline_l124_26;
  reg                 decode_to_execute_HAS_SIDE_EFFECT;
  wire                when_Pipeline_l124_27;
  reg                 execute_to_memory_HAS_SIDE_EFFECT;
  wire                when_Pipeline_l124_28;
  reg                 memory_to_writeBack_HAS_SIDE_EFFECT;
  wire                when_Pipeline_l124_29;
  reg                 decode_to_execute_MEMORY_LRSC;
  wire                when_Pipeline_l124_30;
  reg                 execute_to_memory_MEMORY_LRSC;
  wire                when_Pipeline_l124_31;
  reg                 memory_to_writeBack_MEMORY_LRSC;
  wire                when_Pipeline_l124_32;
  reg                 decode_to_execute_MEMORY_AMO;
  wire                when_Pipeline_l124_33;
  reg                 execute_to_memory_MEMORY_AMO;
  wire                when_Pipeline_l124_34;
  reg                 memory_to_writeBack_MEMORY_AMO;
  wire                when_Pipeline_l124_35;
  reg                 decode_to_execute_MEMORY_MANAGMENT;
  wire                when_Pipeline_l124_36;
  reg                 decode_to_execute_MEMORY_FENCE;
  wire                when_Pipeline_l124_37;
  reg                 execute_to_memory_MEMORY_FENCE;
  wire                when_Pipeline_l124_38;
  reg                 memory_to_writeBack_MEMORY_FENCE;
  wire                when_Pipeline_l124_39;
  reg                 decode_to_execute_IS_CSR;
  wire                when_Pipeline_l124_40;
  reg        [1:0]    decode_to_execute_ENV_CTRL;
  wire                when_Pipeline_l124_41;
  reg        [1:0]    execute_to_memory_ENV_CTRL;
  wire                when_Pipeline_l124_42;
  reg        [1:0]    memory_to_writeBack_ENV_CTRL;
  wire                when_Pipeline_l124_43;
  reg        [1:0]    decode_to_execute_BRANCH_CTRL;
  wire                when_Pipeline_l124_44;
  reg                 decode_to_execute_SRC_LESS_UNSIGNED;
  wire                when_Pipeline_l124_45;
  reg                 decode_to_execute_IS_MUL;
  wire                when_Pipeline_l124_46;
  reg                 execute_to_memory_IS_MUL;
  wire                when_Pipeline_l124_47;
  reg                 memory_to_writeBack_IS_MUL;
  wire                when_Pipeline_l124_48;
  reg                 decode_to_execute_IS_DIV;
  wire                when_Pipeline_l124_49;
  reg                 execute_to_memory_IS_DIV;
  wire                when_Pipeline_l124_50;
  reg                 decode_to_execute_IS_RS1_SIGNED;
  wire                when_Pipeline_l124_51;
  reg                 decode_to_execute_IS_RS2_SIGNED;
  wire                when_Pipeline_l124_52;
  reg                 decode_to_execute_FPU_COMMIT;
  wire                when_Pipeline_l124_53;
  reg                 execute_to_memory_FPU_COMMIT;
  wire                when_Pipeline_l124_54;
  reg                 memory_to_writeBack_FPU_COMMIT;
  wire                when_Pipeline_l124_55;
  reg                 decode_to_execute_FPU_RSP;
  wire                when_Pipeline_l124_56;
  reg                 execute_to_memory_FPU_RSP;
  wire                when_Pipeline_l124_57;
  reg                 memory_to_writeBack_FPU_RSP;
  wire                when_Pipeline_l124_58;
  reg        [3:0]    decode_to_execute_FPU_OPCODE;
  wire                when_Pipeline_l124_59;
  reg        [3:0]    execute_to_memory_FPU_OPCODE;
  wire                when_Pipeline_l124_60;
  reg        [3:0]    memory_to_writeBack_FPU_OPCODE;
  wire                when_Pipeline_l124_61;
  reg                 decode_to_execute_CfuPlugin_CFU_ENABLE;
  wire                when_Pipeline_l124_62;
  reg        [0:0]    decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
  wire                when_Pipeline_l124_63;
  reg        [1:0]    decode_to_execute_ALU_BITWISE_CTRL;
  wire                when_Pipeline_l124_64;
  reg        [1:0]    decode_to_execute_SHIFT_CTRL;
  wire                when_Pipeline_l124_65;
  reg        [1:0]    execute_to_memory_SHIFT_CTRL;
  wire                when_Pipeline_l124_66;
  reg        [31:0]   decode_to_execute_RS1;
  wire                when_Pipeline_l124_67;
  reg        [31:0]   execute_to_memory_RS1;
  wire                when_Pipeline_l124_68;
  reg        [31:0]   memory_to_writeBack_RS1;
  wire                when_Pipeline_l124_69;
  reg        [31:0]   decode_to_execute_RS2;
  wire                when_Pipeline_l124_70;
  reg                 decode_to_execute_SRC2_FORCE_ZERO;
  wire                when_Pipeline_l124_71;
  reg        [31:0]   decode_to_execute_SRC1;
  wire                when_Pipeline_l124_72;
  reg        [31:0]   decode_to_execute_SRC2;
  wire                when_Pipeline_l124_73;
  reg                 decode_to_execute_CSR_WRITE_OPCODE;
  wire                when_Pipeline_l124_74;
  reg                 decode_to_execute_CSR_READ_OPCODE;
  wire                when_Pipeline_l124_75;
  reg                 decode_to_execute_FPU_FORKED;
  wire                when_Pipeline_l124_76;
  reg                 execute_to_memory_FPU_FORKED;
  wire                when_Pipeline_l124_77;
  reg                 memory_to_writeBack_FPU_FORKED;
  wire                when_Pipeline_l124_78;
  reg                 decode_to_execute_FPU_COMMIT_LOAD;
  wire                when_Pipeline_l124_79;
  reg                 execute_to_memory_FPU_COMMIT_LOAD;
  wire                when_Pipeline_l124_80;
  reg                 memory_to_writeBack_FPU_COMMIT_LOAD;
  wire                when_Pipeline_l124_81;
  reg        [31:0]   execute_to_memory_MEMORY_STORE_DATA_RF;
  wire                when_Pipeline_l124_82;
  reg        [31:0]   memory_to_writeBack_MEMORY_STORE_DATA_RF;
  wire                when_Pipeline_l124_83;
  (* keep , syn_keep *) reg        [31:0]   execute_to_memory_MEMORY_VIRTUAL_ADDRESS /* synthesis syn_keep = 1 */ ;
  wire                when_Pipeline_l124_84;
  reg                 execute_to_memory_BRANCH_DO;
  wire                when_Pipeline_l124_85;
  reg        [31:0]   execute_to_memory_BRANCH_CALC;
  wire                when_Pipeline_l124_86;
  reg        [31:0]   execute_to_memory_MUL_LL;
  wire                when_Pipeline_l124_87;
  reg        [33:0]   execute_to_memory_MUL_LH;
  wire                when_Pipeline_l124_88;
  reg        [33:0]   execute_to_memory_MUL_HL;
  wire                when_Pipeline_l124_89;
  reg        [33:0]   execute_to_memory_MUL_HH;
  wire                when_Pipeline_l124_90;
  reg        [33:0]   memory_to_writeBack_MUL_HH;
  wire                when_Pipeline_l124_91;
  reg                 execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
  wire                when_Pipeline_l124_92;
  reg                 memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
  wire                when_Pipeline_l124_93;
  reg        [31:0]   execute_to_memory_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_94;
  reg        [31:0]   memory_to_writeBack_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_95;
  reg        [31:0]   execute_to_memory_SHIFT_RIGHT;
  wire                when_Pipeline_l124_96;
  reg        [51:0]   memory_to_writeBack_MUL_LOW;
  wire                when_Pipeline_l151;
  wire                when_Pipeline_l154;
  wire                when_Pipeline_l151_1;
  wire                when_Pipeline_l154_1;
  wire                when_Pipeline_l151_2;
  wire                when_Pipeline_l154_2;
  reg        [2:0]    IBusCachedPlugin_injector_port_state;
  wire                when_Fetcher_l373;
  wire                when_Fetcher_l391;
  wire                when_Fetcher_l411;
  wire                when_CsrPlugin_l1813;
  reg                 execute_CsrPlugin_csr_1972;
  wire                when_CsrPlugin_l1813_1;
  reg                 execute_CsrPlugin_csr_1969;
  wire                when_CsrPlugin_l1813_2;
  reg                 execute_CsrPlugin_csr_1968;
  wire                when_CsrPlugin_l1813_3;
  reg                 execute_CsrPlugin_csr_3857;
  wire                when_CsrPlugin_l1813_4;
  reg                 execute_CsrPlugin_csr_3858;
  wire                when_CsrPlugin_l1813_5;
  reg                 execute_CsrPlugin_csr_3859;
  wire                when_CsrPlugin_l1813_6;
  reg                 execute_CsrPlugin_csr_3860;
  wire                when_CsrPlugin_l1813_7;
  reg                 execute_CsrPlugin_csr_769;
  wire                when_CsrPlugin_l1813_8;
  reg                 execute_CsrPlugin_csr_768;
  wire                when_CsrPlugin_l1813_9;
  reg                 execute_CsrPlugin_csr_836;
  wire                when_CsrPlugin_l1813_10;
  reg                 execute_CsrPlugin_csr_772;
  wire                when_CsrPlugin_l1813_11;
  reg                 execute_CsrPlugin_csr_773;
  wire                when_CsrPlugin_l1813_12;
  reg                 execute_CsrPlugin_csr_833;
  wire                when_CsrPlugin_l1813_13;
  reg                 execute_CsrPlugin_csr_832;
  wire                when_CsrPlugin_l1813_14;
  reg                 execute_CsrPlugin_csr_834;
  wire                when_CsrPlugin_l1813_15;
  reg                 execute_CsrPlugin_csr_835;
  wire                when_CsrPlugin_l1813_16;
  reg                 execute_CsrPlugin_csr_3;
  wire                when_CsrPlugin_l1813_17;
  reg                 execute_CsrPlugin_csr_2;
  wire                when_CsrPlugin_l1813_18;
  reg                 execute_CsrPlugin_csr_1;
  wire                when_CsrPlugin_l1813_19;
  reg                 execute_CsrPlugin_csr_256;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_1;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_3;
  wire       [1:0]    switch_CsrPlugin_l1167;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_4;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_5;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_6;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_7;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_8;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_9;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_10;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_11;
  wire       [4:0]    _zz_FpuPlugin_flags_NX;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_12;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_13;
  wire       [4:0]    _zz_FpuPlugin_flags_NX_1;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_14;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_15;
  wire                when_CsrPlugin_l1846;
  wire       [11:0]   _zz_when_CsrPlugin_l1853;
  wire                when_CsrPlugin_l1853;
  reg                 when_CsrPlugin_l1863;
  wire                when_CsrPlugin_l1861;
  wire                when_CsrPlugin_l1862;
  wire                when_CsrPlugin_l1869;
  reg        [2:0]    FpuPlugin_stateReg;
  reg        [2:0]    FpuPlugin_stateNext;
  reg        [0:0]    _zz_FpuPlugin_port_cmd_payload_format;
  wire                when_FpuPlugin_l402;
  `ifndef SYNTHESIS
  reg [71:0] _zz_execute_to_memory_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_to_memory_SHIFT_CTRL_1_string;
  reg [71:0] decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_1_string;
  reg [39:0] decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string;
  reg [39:0] decode_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string;
  reg [63:0] memory_FPU_OPCODE_string;
  reg [63:0] _zz_memory_FPU_OPCODE_string;
  reg [63:0] _zz_memory_to_writeBack_FPU_OPCODE_string;
  reg [63:0] _zz_memory_to_writeBack_FPU_OPCODE_1_string;
  reg [63:0] execute_FPU_OPCODE_string;
  reg [63:0] _zz_execute_FPU_OPCODE_string;
  reg [63:0] _zz_execute_to_memory_FPU_OPCODE_string;
  reg [63:0] _zz_execute_to_memory_FPU_OPCODE_1_string;
  reg [63:0] _zz_decode_to_execute_FPU_OPCODE_string;
  reg [63:0] _zz_decode_to_execute_FPU_OPCODE_1_string;
  reg [31:0] decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_1_string;
  reg [47:0] _zz_memory_to_writeBack_ENV_CTRL_string;
  reg [47:0] _zz_memory_to_writeBack_ENV_CTRL_1_string;
  reg [47:0] _zz_execute_to_memory_ENV_CTRL_string;
  reg [47:0] _zz_execute_to_memory_ENV_CTRL_1_string;
  reg [47:0] decode_ENV_CTRL_string;
  reg [47:0] _zz_decode_ENV_CTRL_string;
  reg [47:0] _zz_decode_to_execute_ENV_CTRL_string;
  reg [47:0] _zz_decode_to_execute_ENV_CTRL_1_string;
  reg [63:0] decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_1_string;
  reg [71:0] memory_SHIFT_CTRL_string;
  reg [71:0] _zz_memory_SHIFT_CTRL_string;
  reg [71:0] execute_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_SHIFT_CTRL_string;
  reg [63:0] execute_ALU_CTRL_string;
  reg [63:0] _zz_execute_ALU_CTRL_string;
  reg [39:0] execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [63:0] writeBack_FPU_OPCODE_string;
  reg [63:0] _zz_writeBack_FPU_OPCODE_string;
  reg [47:0] decode_FPU_FORMAT_string;
  reg [47:0] _zz_decode_FPU_FORMAT_string;
  reg [63:0] decode_FPU_OPCODE_string;
  reg [63:0] _zz_decode_FPU_OPCODE_string;
  reg [31:0] execute_BRANCH_CTRL_string;
  reg [31:0] _zz_execute_BRANCH_CTRL_string;
  reg [47:0] memory_ENV_CTRL_string;
  reg [47:0] _zz_memory_ENV_CTRL_string;
  reg [47:0] execute_ENV_CTRL_string;
  reg [47:0] _zz_execute_ENV_CTRL_string;
  reg [47:0] writeBack_ENV_CTRL_string;
  reg [47:0] _zz_writeBack_ENV_CTRL_string;
  reg [23:0] decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_SRC2_CTRL_string;
  reg [95:0] decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_SRC1_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_1_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_1_string;
  reg [39:0] _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string;
  reg [47:0] _zz_decode_FPU_FORMAT_1_string;
  reg [63:0] _zz_decode_FPU_OPCODE_1_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_1_string;
  reg [47:0] _zz_decode_ENV_CTRL_1_string;
  reg [23:0] _zz_decode_SRC2_CTRL_1_string;
  reg [63:0] _zz_decode_ALU_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_1_string;
  reg [71:0] debugBus_dmToHart_payload_op_string;
  reg [63:0] FpuPlugin_port_cmd_payload_opcode_string;
  reg [47:0] FpuPlugin_port_cmd_payload_format_string;
  reg [23:0] FpuPlugin_port_cmd_payload_roundMode_string;
  reg [63:0] FpuPlugin_port_commit_payload_opcode_string;
  reg [95:0] _zz_decode_SRC1_CTRL_2_string;
  reg [63:0] _zz_decode_ALU_CTRL_2_string;
  reg [23:0] _zz_decode_SRC2_CTRL_2_string;
  reg [47:0] _zz_decode_ENV_CTRL_2_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_2_string;
  reg [63:0] _zz_decode_FPU_OPCODE_2_string;
  reg [47:0] _zz_decode_FPU_FORMAT_2_string;
  reg [39:0] _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_2_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_2_string;
  reg [71:0] CsrPlugin_inject_cmd_payload_op_string;
  reg [71:0] CsrPlugin_inject_cmd_toStream_payload_op_string;
  reg [71:0] CsrPlugin_inject_buffer_payload_op_string;
  reg [71:0] CsrPlugin_inject_cmd_toStream_rData_op_string;
  reg [47:0] CsrPlugin_dcsr_stepLogic_stateReg_string;
  reg [47:0] CsrPlugin_dcsr_stepLogic_stateNext_string;
  reg [23:0] _zz_FpuPlugin_port_cmd_payload_roundMode_string;
  reg [23:0] _zz_FpuPlugin_port_cmd_payload_roundMode_1_string;
  reg [63:0] writeBack_FpuPlugin_commit_payload_opcode_string;
  reg [63:0] writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string;
  reg [63:0] writeBack_FpuPlugin_commit_rData_opcode_string;
  reg [63:0] _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string;
  reg [63:0] decode_to_execute_ALU_CTRL_string;
  reg [47:0] decode_to_execute_ENV_CTRL_string;
  reg [47:0] execute_to_memory_ENV_CTRL_string;
  reg [47:0] memory_to_writeBack_ENV_CTRL_string;
  reg [31:0] decode_to_execute_BRANCH_CTRL_string;
  reg [63:0] decode_to_execute_FPU_OPCODE_string;
  reg [63:0] execute_to_memory_FPU_OPCODE_string;
  reg [63:0] memory_to_writeBack_FPU_OPCODE_string;
  reg [39:0] decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string;
  reg [39:0] decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [71:0] decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] execute_to_memory_SHIFT_CTRL_string;
  reg [47:0] FpuPlugin_stateReg_string;
  reg [47:0] FpuPlugin_stateNext_string;
  reg [47:0] _zz_FpuPlugin_port_cmd_payload_format_string;
  `endif

  reg [31:0] RegFilePlugin_regFile [0:31] /* verilator public */ ;

  assign _zz_when = (|{decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid});
  assign _zz_memory_MUL_LOW = ($signed(_zz_memory_MUL_LOW_1) + $signed(_zz_memory_MUL_LOW_4));
  assign _zz_memory_MUL_LOW_1 = ($signed(52'h0) + $signed(_zz_memory_MUL_LOW_2));
  assign _zz_memory_MUL_LOW_3 = {1'b0,memory_MUL_LL};
  assign _zz_memory_MUL_LOW_2 = {{19{_zz_memory_MUL_LOW_3[32]}}, _zz_memory_MUL_LOW_3};
  assign _zz_memory_MUL_LOW_5 = ({16'd0,memory_MUL_LH} <<< 5'd16);
  assign _zz_memory_MUL_LOW_4 = {{2{_zz_memory_MUL_LOW_5[49]}}, _zz_memory_MUL_LOW_5};
  assign _zz_memory_MUL_LOW_7 = ({16'd0,memory_MUL_HL} <<< 5'd16);
  assign _zz_memory_MUL_LOW_6 = {{2{_zz_memory_MUL_LOW_7[49]}}, _zz_memory_MUL_LOW_7};
  assign _zz_decode_FORMAL_PC_NEXT_1 = (decode_IS_RVC ? 3'b010 : 3'b100);
  assign _zz_decode_FORMAL_PC_NEXT = {29'd0, _zz_decode_FORMAL_PC_NEXT_1};
  assign _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload - 3'b001);
  assign _zz_IBusCachedPlugin_fetchPc_pc_1 = {IBusCachedPlugin_fetchPc_inc,2'b00};
  assign _zz_IBusCachedPlugin_fetchPc_pc = {29'd0, _zz_IBusCachedPlugin_fetchPc_pc_1};
  assign _zz_IBusCachedPlugin_decodePc_pcPlus_1 = (decode_IS_RVC ? 3'b010 : 3'b100);
  assign _zz_IBusCachedPlugin_decodePc_pcPlus = {29'd0, _zz_IBusCachedPlugin_decodePc_pcPlus_1};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_31 = {{_zz_IBusCachedPlugin_decompressor_decompressed_11,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},12'h0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_38 = {{{3'b000,_zz_IBusCachedPlugin_decompressor_decompressed[9 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},3'b000};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_39 = {{{3'b000,_zz_IBusCachedPlugin_decompressor_decompressed[9 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},3'b000};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_40 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_41 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_42 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_43 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[8 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 9]},2'b00};
  assign _zz_io_cpu_flush_payload_lineId = _zz_io_cpu_flush_payload_lineId_1;
  assign _zz_io_cpu_flush_payload_lineId_1 = (execute_RS1 >>> 3'd6);
  assign _zz_DBusCachedPlugin_exceptionBus_payload_code = (writeBack_MEMORY_WR ? 3'b111 : 3'b101);
  assign _zz_DBusCachedPlugin_exceptionBus_payload_code_1 = (writeBack_MEMORY_WR ? 3'b110 : 3'b100);
  assign _zz_writeBack_DBusCachedPlugin_rspRf = (! dataCache_2_io_cpu_writeBack_exclusiveOk);
  assign _zz__zz_decode_SRC1 = (decode_IS_RVC ? 3'b010 : 3'b100);
  assign _zz__zz_decode_SRC1_1 = decode_INSTRUCTION[19 : 15];
  assign _zz__zz_decode_SRC2_2 = {decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]};
  assign _zz_execute_SrcPlugin_addSub = ($signed(_zz_execute_SrcPlugin_addSub_1) + $signed(_zz_execute_SrcPlugin_addSub_4));
  assign _zz_execute_SrcPlugin_addSub_1 = ($signed(_zz_execute_SrcPlugin_addSub_2) + $signed(_zz_execute_SrcPlugin_addSub_3));
  assign _zz_execute_SrcPlugin_addSub_2 = execute_SRC1;
  assign _zz_execute_SrcPlugin_addSub_3 = (execute_SRC_USE_SUB_LESS ? (~ execute_SRC2) : execute_SRC2);
  assign _zz_execute_SrcPlugin_addSub_4 = (execute_SRC_USE_SUB_LESS ? 32'h00000001 : 32'h0);
  assign _zz_CsrPlugin_timeout_counter_valueNext_1 = CsrPlugin_timeout_counter_willIncrement;
  assign _zz_CsrPlugin_timeout_counter_valueNext = {2'd0, _zz_CsrPlugin_timeout_counter_valueNext_1};
  assign _zz__zz_6 = debugBus_dmToHart_payload_address[0:0];
  assign _zz_CsrPlugin_counters_mcycle_1 = ((! debugMode) || (! CsrPlugin_dcsr_stopcount));
  assign _zz_CsrPlugin_counters_mcycle = {63'd0, _zz_CsrPlugin_counters_mcycle_1};
  assign _zz_CsrPlugin_counters_minstret_1 = ((! debugMode) || (! CsrPlugin_dcsr_stopcount));
  assign _zz_CsrPlugin_counters_minstret = {63'd0, _zz_CsrPlugin_counters_minstret_1};
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code & (~ _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1));
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code - 2'b01);
  assign _zz__zz_execute_BranchPlugin_branch_src2 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]};
  assign _zz__zz_execute_BranchPlugin_branch_src2_4 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]};
  assign _zz_writeBack_MulPlugin_result = {{14{writeBack_MUL_LOW[51]}}, writeBack_MUL_LOW};
  assign _zz_writeBack_MulPlugin_result_1 = ({32'd0,writeBack_MUL_HH} <<< 6'd32);
  assign _zz__zz_decode_RS2_2 = writeBack_MUL_LOW[31 : 0];
  assign _zz__zz_decode_RS2_2_1 = writeBack_MulPlugin_result[63 : 32];
  assign _zz_memory_MulDivIterativePlugin_div_counter_valueNext_1 = memory_MulDivIterativePlugin_div_counter_willIncrement;
  assign _zz_memory_MulDivIterativePlugin_div_counter_valueNext = {5'd0, _zz_memory_MulDivIterativePlugin_div_counter_valueNext_1};
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator = {1'd0, memory_MulDivIterativePlugin_rs2};
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder = memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator[31:0];
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder_1 = memory_MulDivIterativePlugin_div_stage_0_remainderShifted[31:0];
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_outNumerator = {_zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted,(! memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator[32])};
  assign _zz_memory_MulDivIterativePlugin_div_result_1 = _zz_memory_MulDivIterativePlugin_div_result_2;
  assign _zz_memory_MulDivIterativePlugin_div_result_2 = _zz_memory_MulDivIterativePlugin_div_result_3;
  assign _zz_memory_MulDivIterativePlugin_div_result_3 = ({memory_MulDivIterativePlugin_div_needRevert,(memory_MulDivIterativePlugin_div_needRevert ? (~ _zz_memory_MulDivIterativePlugin_div_result) : _zz_memory_MulDivIterativePlugin_div_result)} + _zz_memory_MulDivIterativePlugin_div_result_4);
  assign _zz_memory_MulDivIterativePlugin_div_result_5 = memory_MulDivIterativePlugin_div_needRevert;
  assign _zz_memory_MulDivIterativePlugin_div_result_4 = {32'd0, _zz_memory_MulDivIterativePlugin_div_result_5};
  assign _zz_memory_MulDivIterativePlugin_rs1_3 = _zz_memory_MulDivIterativePlugin_rs1;
  assign _zz_memory_MulDivIterativePlugin_rs1_2 = {32'd0, _zz_memory_MulDivIterativePlugin_rs1_3};
  assign _zz_memory_MulDivIterativePlugin_rs2_2 = _zz_memory_MulDivIterativePlugin_rs2;
  assign _zz_memory_MulDivIterativePlugin_rs2_1 = {31'd0, _zz_memory_MulDivIterativePlugin_rs2_2};
  assign _zz_FpuPlugin_pendings = (_zz_FpuPlugin_pendings_1 - _zz_FpuPlugin_pendings_4);
  assign _zz_FpuPlugin_pendings_1 = (FpuPlugin_pendings + _zz_FpuPlugin_pendings_2);
  assign _zz_FpuPlugin_pendings_3 = FpuPlugin_port_cmd_fire;
  assign _zz_FpuPlugin_pendings_2 = {5'd0, _zz_FpuPlugin_pendings_3};
  assign _zz_FpuPlugin_pendings_5 = FpuPlugin_port_completion_valid;
  assign _zz_FpuPlugin_pendings_4 = {5'd0, _zz_FpuPlugin_pendings_5};
  assign _zz_FpuPlugin_pendings_7 = FpuPlugin_port_rsp_fire;
  assign _zz_FpuPlugin_pendings_6 = {5'd0, _zz_FpuPlugin_pendings_7};
  assign _zz_when_CsrPlugin_l1862 = (execute_CsrPlugin_csrAddress >>> 3'd4);
  assign _zz_decode_RegFilePlugin_rs1Data = 1'b1;
  assign _zz_decode_RegFilePlugin_rs2Data = 1'b1;
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_5 = {_zz_IBusCachedPlugin_jump_pcLoad_payload_3,_zz_IBusCachedPlugin_jump_pcLoad_payload_2};
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_1 = dataCache_2_io_cpu_writeBack_address[2 : 0];
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_3 = dataCache_2_io_cpu_writeBack_address[2 : 1];
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_5 = dataCache_2_io_cpu_writeBack_address[2 : 2];
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_7 = dataCache_2_io_cpu_writeBack_address[2 : 2];
  assign _zz_decode_LEGAL_INSTRUCTION = 32'h0000007f;
  assign _zz_decode_LEGAL_INSTRUCTION_1 = (decode_INSTRUCTION & 32'h0000007f);
  assign _zz_decode_LEGAL_INSTRUCTION_2 = 32'h0000000b;
  assign _zz_decode_LEGAL_INSTRUCTION_3 = ((decode_INSTRUCTION & 32'h0000107f) == 32'h00001073);
  assign _zz_decode_LEGAL_INSTRUCTION_4 = ((decode_INSTRUCTION & 32'h0000207f) == 32'h00002073);
  assign _zz_decode_LEGAL_INSTRUCTION_5 = {((decode_INSTRUCTION & 32'h0000407f) == 32'h00004063),{((decode_INSTRUCTION & 32'h0000207f) == 32'h00002013),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_6) == 32'h00002007),{(_zz_decode_LEGAL_INSTRUCTION_7 == _zz_decode_LEGAL_INSTRUCTION_8),{_zz_decode_LEGAL_INSTRUCTION_9,{_zz_decode_LEGAL_INSTRUCTION_10,_zz_decode_LEGAL_INSTRUCTION_11}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_6 = 32'h0000605f;
  assign _zz_decode_LEGAL_INSTRUCTION_7 = (decode_INSTRUCTION & 32'h0000705b);
  assign _zz_decode_LEGAL_INSTRUCTION_8 = 32'h00002003;
  assign _zz_decode_LEGAL_INSTRUCTION_9 = ((decode_INSTRUCTION & 32'h0000107f) == 32'h00000013);
  assign _zz_decode_LEGAL_INSTRUCTION_10 = ((decode_INSTRUCTION & 32'h0000603f) == 32'h00000023);
  assign _zz_decode_LEGAL_INSTRUCTION_11 = {((decode_INSTRUCTION & 32'h0000207f) == 32'h00000003),{((decode_INSTRUCTION & 32'h0000707b) == 32'h00000063),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_12) == 32'h0000000f),{(_zz_decode_LEGAL_INSTRUCTION_13 == _zz_decode_LEGAL_INSTRUCTION_14),{_zz_decode_LEGAL_INSTRUCTION_15,{_zz_decode_LEGAL_INSTRUCTION_16,_zz_decode_LEGAL_INSTRUCTION_17}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_12 = 32'h0000607f;
  assign _zz_decode_LEGAL_INSTRUCTION_13 = (decode_INSTRUCTION & 32'he400007f);
  assign _zz_decode_LEGAL_INSTRUCTION_14 = 32'h00000053;
  assign _zz_decode_LEGAL_INSTRUCTION_15 = ((decode_INSTRUCTION & 32'h1800707f) == 32'h0000202f);
  assign _zz_decode_LEGAL_INSTRUCTION_16 = ((decode_INSTRUCTION & 32'hfc00007f) == 32'h00000033);
  assign _zz_decode_LEGAL_INSTRUCTION_17 = {((decode_INSTRUCTION & 32'he800707f) == 32'h0800202f),{((decode_INSTRUCTION & 32'h7c00607f) == 32'h20000053),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_18) == 32'h20000053),{(_zz_decode_LEGAL_INSTRUCTION_19 == _zz_decode_LEGAL_INSTRUCTION_20),{_zz_decode_LEGAL_INSTRUCTION_21,{_zz_decode_LEGAL_INSTRUCTION_22,_zz_decode_LEGAL_INSTRUCTION_23}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_18 = 32'h7c00507f;
  assign _zz_decode_LEGAL_INSTRUCTION_19 = (decode_INSTRUCTION & 32'hf400607f);
  assign _zz_decode_LEGAL_INSTRUCTION_20 = 32'h20000053;
  assign _zz_decode_LEGAL_INSTRUCTION_21 = ((decode_INSTRUCTION & 32'h01f0707f) == 32'h0000500f);
  assign _zz_decode_LEGAL_INSTRUCTION_22 = ((decode_INSTRUCTION & 32'hbe00705f) == 32'h00005013);
  assign _zz_decode_LEGAL_INSTRUCTION_23 = {((decode_INSTRUCTION & 32'hfe00305f) == 32'h00001013),{((decode_INSTRUCTION & 32'hede0007f) == 32'hc0000053),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_24) == 32'h00000033),{(_zz_decode_LEGAL_INSTRUCTION_25 == _zz_decode_LEGAL_INSTRUCTION_26),{_zz_decode_LEGAL_INSTRUCTION_27,{_zz_decode_LEGAL_INSTRUCTION_28,_zz_decode_LEGAL_INSTRUCTION_29}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_24 = 32'hbe00707f;
  assign _zz_decode_LEGAL_INSTRUCTION_25 = (decode_INSTRUCTION & 32'hfdf0007f);
  assign _zz_decode_LEGAL_INSTRUCTION_26 = 32'h58000053;
  assign _zz_decode_LEGAL_INSTRUCTION_27 = ((decode_INSTRUCTION & 32'h7ff0007f) == 32'h42000053);
  assign _zz_decode_LEGAL_INSTRUCTION_28 = ((decode_INSTRUCTION & 32'h7ff0007f) == 32'h40100053);
  assign _zz_decode_LEGAL_INSTRUCTION_29 = {((decode_INSTRUCTION & 32'hf9f0707f) == 32'h1000202f),{((decode_INSTRUCTION & 32'hfdf0707f) == 32'he0001053),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_30) == 32'he0000053),{(_zz_decode_LEGAL_INSTRUCTION_31 == _zz_decode_LEGAL_INSTRUCTION_32),{_zz_decode_LEGAL_INSTRUCTION_33,_zz_decode_LEGAL_INSTRUCTION_34}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_30 = 32'heff0707f;
  assign _zz_decode_LEGAL_INSTRUCTION_31 = (decode_INSTRUCTION & 32'hdfffffff);
  assign _zz_decode_LEGAL_INSTRUCTION_32 = 32'h10200073;
  assign _zz_decode_LEGAL_INSTRUCTION_33 = ((decode_INSTRUCTION & 32'hffefffff) == 32'h00000073);
  assign _zz_decode_LEGAL_INSTRUCTION_34 = ((decode_INSTRUCTION & 32'hffffffff) == 32'h10500073);
  assign _zz_IBusCachedPlugin_decompressor_decompressed_28 = {_zz_IBusCachedPlugin_decompressor_decompressed_13,_zz_IBusCachedPlugin_decompressor_decompressed[4 : 3]};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_29 = _zz_IBusCachedPlugin_decompressor_decompressed[5];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_30 = _zz_IBusCachedPlugin_decompressor_decompressed[2];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_32 = (_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] == 2'b01);
  assign _zz_IBusCachedPlugin_decompressor_decompressed_33 = ((_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] == 2'b11) && (_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5] == 2'b00));
  assign _zz_IBusCachedPlugin_decompressor_decompressed_34 = 7'h0;
  assign _zz_IBusCachedPlugin_decompressor_decompressed_35 = _zz_IBusCachedPlugin_decompressor_decompressed[6 : 2];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_36 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  assign _zz_IBusCachedPlugin_decompressor_decompressed_37 = _zz_IBusCachedPlugin_decompressor_decompressed[11 : 7];
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE = (decode_INSTRUCTION & 32'h40003054);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_1 = 32'h40001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_2 = (decode_INSTRUCTION & 32'h02007054);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_3 = 32'h00001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_4 = (decode_INSTRUCTION & 32'h00001000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_5 = 32'h00001000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_6 = ((decode_INSTRUCTION & 32'h00003000) == 32'h00002000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_7 = (|_zz_decode_CfuPlugin_CFU_ENABLE_10);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_8 = (|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE_9 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_10),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_11 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_12)});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_13 = {(|{_zz_decode_CfuPlugin_CFU_ENABLE_7,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_14,_zz__zz_decode_CfuPlugin_CFU_ENABLE_17}}),{(|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_22,_zz__zz_decode_CfuPlugin_CFU_ENABLE_25}),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_40),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_49,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_58,_zz__zz_decode_CfuPlugin_CFU_ENABLE_70}}}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_9 = (decode_INSTRUCTION & 32'h00000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_10 = 32'h00000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_11 = (decode_INSTRUCTION & 32'h20002010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_12 = 32'h20002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_14 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_15 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_16);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_17 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_18,_zz__zz_decode_CfuPlugin_CFU_ENABLE_20};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_22 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_23 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_24);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_25 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_26,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_28,_zz__zz_decode_CfuPlugin_CFU_ENABLE_31}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_40 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_41,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_43,_zz__zz_decode_CfuPlugin_CFU_ENABLE_46}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_49 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_50,_zz__zz_decode_CfuPlugin_CFU_ENABLE_53});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_58 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_59);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_70 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_71,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_80,_zz__zz_decode_CfuPlugin_CFU_ENABLE_82}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_15 = (decode_INSTRUCTION & 32'h20001010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_16 = 32'h20001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_18 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_19) == 32'h08000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_20 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_21) == 32'h80000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_23 = (decode_INSTRUCTION & 32'h00001040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_24 = 32'h00001000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_26 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_27) == 32'h82000000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_28 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_29 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_30);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_31 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_32,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_34,_zz__zz_decode_CfuPlugin_CFU_ENABLE_37}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_41 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_42) == 32'h60000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_43 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_44 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_45);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_46 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_47,_zz_decode_CfuPlugin_CFU_ENABLE_13};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_50 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_51 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_52);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_53 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_54,_zz__zz_decode_CfuPlugin_CFU_ENABLE_56};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_59 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_60,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_62,_zz__zz_decode_CfuPlugin_CFU_ENABLE_65}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_71 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_72,_zz__zz_decode_CfuPlugin_CFU_ENABLE_73});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_80 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_81);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_82 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_83,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_90,_zz__zz_decode_CfuPlugin_CFU_ENABLE_94}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_19 = 32'h28000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_21 = 32'ha0100010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_27 = 32'h82000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_29 = (decode_INSTRUCTION & 32'h02000050);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_30 = 32'h02000040;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_32 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_33) == 32'h12000000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_34 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_35 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_36);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_37 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_38 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_39);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_42 = 32'h60000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_44 = (decode_INSTRUCTION & 32'h18000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_45 = 32'h18000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_47 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_48) == 32'h20000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_51 = (decode_INSTRUCTION & 32'h80000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_52 = 32'h80000000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_54 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_55) == 32'h00000040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_56 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_57) == 32'h40000000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_60 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_61) == 32'h00001010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_62 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_63 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_64);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_65 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_66,_zz__zz_decode_CfuPlugin_CFU_ENABLE_68};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_72 = _zz_decode_CfuPlugin_CFU_ENABLE_12;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_73 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_74,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_76,_zz__zz_decode_CfuPlugin_CFU_ENABLE_77}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_81 = {_zz_decode_CfuPlugin_CFU_ENABLE_12,_zz_decode_CfuPlugin_CFU_ENABLE_8};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_83 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_84,_zz__zz_decode_CfuPlugin_CFU_ENABLE_87});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_90 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_91);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_94 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_95,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_96,_zz__zz_decode_CfuPlugin_CFU_ENABLE_98}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_33 = 32'h12000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_35 = (decode_INSTRUCTION & 32'h42000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_36 = 32'h02000000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_38 = (decode_INSTRUCTION & 32'hd2000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_39 = 32'h40000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_48 = 32'ha0000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_55 = 32'h00000050;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_57 = 32'h50000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_61 = 32'h10001010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_63 = (decode_INSTRUCTION & 32'h30000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_64 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_66 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_67) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_68 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_69) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_74 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_75) == 32'h90000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_76 = _zz_decode_CfuPlugin_CFU_ENABLE_13;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_77 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_78,_zz__zz_decode_CfuPlugin_CFU_ENABLE_79};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_84 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_85 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_86);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_87 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_88,_zz__zz_decode_CfuPlugin_CFU_ENABLE_89};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_91 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_92,_zz__zz_decode_CfuPlugin_CFU_ENABLE_93};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_95 = (|_zz_decode_CfuPlugin_CFU_ENABLE_11);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_96 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_97);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_98 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_99,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_102,_zz__zz_decode_CfuPlugin_CFU_ENABLE_104}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_67 = 32'h88000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_69 = 32'h50000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_75 = 32'h90000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_78 = ((decode_INSTRUCTION & 32'h58000010) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_79 = ((decode_INSTRUCTION & 32'hb0000010) == 32'h00000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_85 = (decode_INSTRUCTION & 32'h10000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_86 = 32'h10000000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_88 = ((decode_INSTRUCTION & 32'h80000020) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_89 = ((decode_INSTRUCTION & 32'h00000030) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_92 = ((decode_INSTRUCTION & 32'h00000060) == 32'h00000040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_93 = ((decode_INSTRUCTION & 32'h0000005c) == 32'h00000004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_97 = _zz_decode_CfuPlugin_CFU_ENABLE_11;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_99 = (|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_100 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_101));
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_102 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_103);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_104 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_105),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_108,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_113,_zz__zz_decode_CfuPlugin_CFU_ENABLE_116}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_100 = (decode_INSTRUCTION & 32'h02004064);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_101 = 32'h02004020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_103 = ((decode_INSTRUCTION & 32'h02004074) == 32'h02000030);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_105 = {((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_106) == 32'h00002000),((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_107) == 32'h00001000)};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_108 = (|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE_109 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_110),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_111 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_112)});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_113 = (|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_114 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_115));
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_116 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_117),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_118),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_121,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_126,_zz__zz_decode_CfuPlugin_CFU_ENABLE_129}}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_106 = 32'h00002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_107 = 32'h00005000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_109 = (decode_INSTRUCTION & 32'h00000068);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_110 = 32'h00000068;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_111 = (decode_INSTRUCTION & 32'h00002034);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_112 = 32'h00000024;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_114 = (decode_INSTRUCTION & 32'h00000078);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_115 = 32'h00000060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_117 = ((decode_INSTRUCTION & 32'h10003070) == 32'h00000070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_118 = {((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_119) == 32'h00100070),((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_120) == 32'h10000030)};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_121 = (|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE_122 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_123),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_124 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_125)});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_126 = (|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_127 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_128));
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_129 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_130),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_131),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_136,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_146,_zz__zz_decode_CfuPlugin_CFU_ENABLE_148}}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_119 = 32'h10103070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_120 = 32'h10403034;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_122 = (decode_INSTRUCTION & 32'h00001070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_123 = 32'h00001070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_124 = (decode_INSTRUCTION & 32'h00002070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_125 = 32'h00002070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_127 = (decode_INSTRUCTION & 32'h00003054);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_128 = 32'h00000004;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_130 = ((decode_INSTRUCTION & 32'h00004054) == 32'h00004004);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_131 = {(_zz__zz_decode_CfuPlugin_CFU_ENABLE_132 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_133),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_134 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_135)};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_136 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_137,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_138,_zz__zz_decode_CfuPlugin_CFU_ENABLE_139}});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_146 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_147);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_148 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_149),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_151,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_166,_zz__zz_decode_CfuPlugin_CFU_ENABLE_175}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_132 = (decode_INSTRUCTION & 32'h00000034);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_133 = 32'h00000034;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_134 = (decode_INSTRUCTION & 32'h00000068);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_135 = 32'h00000028;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_137 = ((decode_INSTRUCTION & 32'h00000034) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_138 = _zz_decode_CfuPlugin_CFU_ENABLE_10;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_139 = {(_zz__zz_decode_CfuPlugin_CFU_ENABLE_140 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_141),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_142,_zz__zz_decode_CfuPlugin_CFU_ENABLE_144}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_147 = ((decode_INSTRUCTION & 32'h10000008) == 32'h00000008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_149 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_150) == 32'h10000008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_151 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_152,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_154,_zz__zz_decode_CfuPlugin_CFU_ENABLE_157}});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_166 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_167,_zz__zz_decode_CfuPlugin_CFU_ENABLE_170});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_175 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_176),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_189,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_202,_zz__zz_decode_CfuPlugin_CFU_ENABLE_220}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_140 = (decode_INSTRUCTION & 32'h00000064);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_141 = 32'h00000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_142 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_143) == 32'h08002008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_144 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_145) == 32'h00002008);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_150 = 32'h10000008;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_152 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_153) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_154 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_155 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_156);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_157 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_158,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_160,_zz__zz_decode_CfuPlugin_CFU_ENABLE_163}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_167 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_168 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_169);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_170 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_171,_zz__zz_decode_CfuPlugin_CFU_ENABLE_173};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_176 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_177,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_179,_zz__zz_decode_CfuPlugin_CFU_ENABLE_182}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_189 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_190,_zz__zz_decode_CfuPlugin_CFU_ENABLE_191});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_202 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_203);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_220 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_221,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_226,_zz__zz_decode_CfuPlugin_CFU_ENABLE_232}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_143 = 32'h08002048;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_145 = 32'h10002048;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_153 = 32'h00000030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_155 = (decode_INSTRUCTION & 32'h00001060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_156 = 32'h00001060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_158 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_159) == 32'h00002060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_160 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_161 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_162);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_163 = {_zz_decode_CfuPlugin_CFU_ENABLE_4,_zz__zz_decode_CfuPlugin_CFU_ENABLE_164};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_168 = (decode_INSTRUCTION & 32'h08000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_169 = 32'h08000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_171 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_172) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_173 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_174) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_177 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_178) == 32'h00004020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_179 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_180 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_181);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_182 = {_zz_decode_CfuPlugin_CFU_ENABLE_9,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_183,_zz__zz_decode_CfuPlugin_CFU_ENABLE_186}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_190 = _zz_decode_CfuPlugin_CFU_ENABLE_9;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_191 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_192,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_194,_zz__zz_decode_CfuPlugin_CFU_ENABLE_197}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_203 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_204,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_206,_zz__zz_decode_CfuPlugin_CFU_ENABLE_209}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_221 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_222,_zz__zz_decode_CfuPlugin_CFU_ENABLE_223});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_226 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_227);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_232 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_233,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_236,_zz__zz_decode_CfuPlugin_CFU_ENABLE_240}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_159 = 32'h00002060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_161 = (decode_INSTRUCTION & 32'h10000060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_162 = 32'h00000060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_164 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_165) == 32'h10000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_172 = 32'h10000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_174 = 32'h00000028;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_178 = 32'h00004020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_180 = (decode_INSTRUCTION & 32'h00000060);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_181 = 32'h00000060;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_183 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_184 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_185);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_186 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_187 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_188);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_192 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_193) == 32'h00002010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_194 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_195 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_196);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_197 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_198,_zz__zz_decode_CfuPlugin_CFU_ENABLE_200};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_204 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_205) == 32'h00000028);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_206 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_207 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_208);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_209 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_210,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_212,_zz__zz_decode_CfuPlugin_CFU_ENABLE_215}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_222 = _zz_decode_CfuPlugin_CFU_ENABLE_7;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_223 = {_zz_decode_CfuPlugin_CFU_ENABLE_3,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_224,_zz__zz_decode_CfuPlugin_CFU_ENABLE_225}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_227 = {_zz_decode_CfuPlugin_CFU_ENABLE_7,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_228,_zz__zz_decode_CfuPlugin_CFU_ENABLE_231}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_233 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_234);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_236 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_237);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_240 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_241,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_256,_zz__zz_decode_CfuPlugin_CFU_ENABLE_258}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_165 = 32'h10400024;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_184 = (decode_INSTRUCTION & 32'h82000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_185 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_187 = (decode_INSTRUCTION & 32'h00000070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_188 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_193 = 32'h00002070;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_195 = (decode_INSTRUCTION & 32'h00001070);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_196 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_198 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_199) == 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_200 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_201) == 32'h00002020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_205 = 32'h00000028;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_207 = (decode_INSTRUCTION & 32'h00000050);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_208 = 32'h00000010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_210 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_211) == 32'h00001030);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_212 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_213 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_214);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_215 = {_zz_decode_CfuPlugin_CFU_ENABLE_8,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_216,_zz__zz_decode_CfuPlugin_CFU_ENABLE_218}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_224 = _zz_decode_CfuPlugin_CFU_ENABLE_6;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_225 = _zz_decode_CfuPlugin_CFU_ENABLE_5;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_228 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_229 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_230);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_231 = _zz_decode_CfuPlugin_CFU_ENABLE_6;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_234 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_235) == 32'h00004010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_237 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_238 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_239);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_241 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_242,_zz__zz_decode_CfuPlugin_CFU_ENABLE_244});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_256 = (|_zz__zz_decode_CfuPlugin_CFU_ENABLE_257);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_258 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_259,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_268,_zz__zz_decode_CfuPlugin_CFU_ENABLE_274}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_199 = 32'h02003020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_201 = 32'h02002068;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_211 = 32'h00001030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_213 = (decode_INSTRUCTION & 32'h00002030);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_214 = 32'h00002030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_216 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_217) == 32'h00000024);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_218 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_219) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_229 = (decode_INSTRUCTION & 32'h00000020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_230 = 32'h0;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_235 = 32'h00004014;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_238 = (decode_INSTRUCTION & 32'h00006014);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_239 = 32'h00002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_242 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_243) == 32'h0);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_244 = {(_zz__zz_decode_CfuPlugin_CFU_ENABLE_245 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_246),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_247,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_249,_zz__zz_decode_CfuPlugin_CFU_ENABLE_252}}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_257 = {_zz_decode_CfuPlugin_CFU_ENABLE_5,_zz_decode_CfuPlugin_CFU_ENABLE_4};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_259 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_260,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_262,_zz__zz_decode_CfuPlugin_CFU_ENABLE_265}});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_268 = (|{_zz__zz_decode_CfuPlugin_CFU_ENABLE_269,_zz__zz_decode_CfuPlugin_CFU_ENABLE_272});
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_274 = {(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_275),{_zz__zz_decode_CfuPlugin_CFU_ENABLE_276,_zz__zz_decode_CfuPlugin_CFU_ENABLE_277}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_217 = 32'h00002024;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_219 = 32'h00000064;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_243 = 32'h00000044;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_245 = (decode_INSTRUCTION & 32'h00000038);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_246 = 32'h00000020;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_247 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_248) == 32'h00004000);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_249 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_250 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_251);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_252 = {_zz__zz_decode_CfuPlugin_CFU_ENABLE_253,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_254,_zz__zz_decode_CfuPlugin_CFU_ENABLE_255}};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_260 = ((decode_INSTRUCTION & _zz__zz_decode_CfuPlugin_CFU_ENABLE_261) == 32'h00000040);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_262 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_263 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_264);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_265 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_266 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_267);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_269 = (_zz__zz_decode_CfuPlugin_CFU_ENABLE_270 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_271);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_272 = {_zz_decode_CfuPlugin_CFU_ENABLE_2,_zz__zz_decode_CfuPlugin_CFU_ENABLE_273};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_275 = {_zz_decode_CfuPlugin_CFU_ENABLE_3,_zz_decode_CfuPlugin_CFU_ENABLE_2};
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_276 = (|_zz_decode_CfuPlugin_CFU_ENABLE_1);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_277 = (|_zz_decode_CfuPlugin_CFU_ENABLE_1);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_248 = 32'h00004050;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_250 = (decode_INSTRUCTION & 32'h00002050);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_251 = 32'h00002000;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_253 = ((decode_INSTRUCTION & 32'h00006024) == 32'h00002020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_254 = ((decode_INSTRUCTION & 32'h00005024) == 32'h00001020);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_255 = ((decode_INSTRUCTION & 32'h90000034) == 32'h90000010);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_261 = 32'h00000044;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_263 = (decode_INSTRUCTION & 32'h00002014);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_264 = 32'h00002010;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_266 = (decode_INSTRUCTION & 32'h40000034);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_267 = 32'h40000030;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_270 = (decode_INSTRUCTION & 32'h00000048);
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_271 = 32'h00000048;
  assign _zz__zz_decode_CfuPlugin_CFU_ENABLE_273 = ((decode_INSTRUCTION & 32'h00002014) == 32'h00000004);
  assign _zz_CsrPlugin_csrMapping_readDataInit_16 = 32'h0;
  assign _zz_CsrPlugin_csrMapping_readDataInit_17 = 32'h0;
  assign _zz_CsrPlugin_csrMapping_readDataInit_18 = 32'h0;
  assign _zz_CsrPlugin_csrMapping_readDataInit_19 = 32'h0;
  always @(posedge io_systemClk) begin
    if(_zz_decode_RegFilePlugin_rs1Data) begin
      RegFilePlugin_regFile_spinal_port0 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress1];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_decode_RegFilePlugin_rs2Data) begin
      RegFilePlugin_regFile_spinal_port1 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress2];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      RegFilePlugin_regFile[lastStageRegFileWrite_payload_address] <= lastStageRegFileWrite_payload_data;
    end
  end

  InstructionCache IBusCachedPlugin_cache (
    .io_flush                              (IBusCachedPlugin_cache_io_flush                           ), //i
    .io_cpu_prefetch_isValid               (IBusCachedPlugin_cache_io_cpu_prefetch_isValid            ), //i
    .io_cpu_prefetch_haltIt                (IBusCachedPlugin_cache_io_cpu_prefetch_haltIt             ), //o
    .io_cpu_prefetch_pc                    (IBusCachedPlugin_iBusRsp_stages_0_input_payload[31:0]     ), //i
    .io_cpu_fetch_isValid                  (IBusCachedPlugin_cache_io_cpu_fetch_isValid               ), //i
    .io_cpu_fetch_isStuck                  (IBusCachedPlugin_cache_io_cpu_fetch_isStuck               ), //i
    .io_cpu_fetch_isRemoved                (IBusCachedPlugin_cache_io_cpu_fetch_isRemoved             ), //i
    .io_cpu_fetch_pc                       (IBusCachedPlugin_iBusRsp_stages_1_input_payload[31:0]     ), //i
    .io_cpu_fetch_data                     (IBusCachedPlugin_cache_io_cpu_fetch_data[31:0]            ), //o
    .io_cpu_fetch_mmuRsp_physicalAddress   (IBusCachedPlugin_mmuBus_rsp_physicalAddress[31:0]         ), //i
    .io_cpu_fetch_mmuRsp_isIoAccess        (IBusCachedPlugin_mmuBus_rsp_isIoAccess                    ), //i
    .io_cpu_fetch_mmuRsp_isPaging          (IBusCachedPlugin_mmuBus_rsp_isPaging                      ), //i
    .io_cpu_fetch_mmuRsp_allowRead         (IBusCachedPlugin_mmuBus_rsp_allowRead                     ), //i
    .io_cpu_fetch_mmuRsp_allowWrite        (IBusCachedPlugin_mmuBus_rsp_allowWrite                    ), //i
    .io_cpu_fetch_mmuRsp_allowExecute      (IBusCachedPlugin_mmuBus_rsp_allowExecute                  ), //i
    .io_cpu_fetch_mmuRsp_exception         (IBusCachedPlugin_mmuBus_rsp_exception                     ), //i
    .io_cpu_fetch_mmuRsp_refilling         (IBusCachedPlugin_mmuBus_rsp_refilling                     ), //i
    .io_cpu_fetch_mmuRsp_bypassTranslation (IBusCachedPlugin_mmuBus_rsp_bypassTranslation             ), //i
    .io_cpu_fetch_physicalAddress          (IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress[31:0] ), //o
    .io_cpu_decode_isValid                 (IBusCachedPlugin_cache_io_cpu_decode_isValid              ), //i
    .io_cpu_decode_isStuck                 (IBusCachedPlugin_cache_io_cpu_decode_isStuck              ), //i
    .io_cpu_decode_pc                      (IBusCachedPlugin_iBusRsp_stages_2_input_payload[31:0]     ), //i
    .io_cpu_decode_physicalAddress         (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31:0]), //o
    .io_cpu_decode_data                    (IBusCachedPlugin_cache_io_cpu_decode_data[31:0]           ), //o
    .io_cpu_decode_cacheMiss               (IBusCachedPlugin_cache_io_cpu_decode_cacheMiss            ), //o
    .io_cpu_decode_error                   (IBusCachedPlugin_cache_io_cpu_decode_error                ), //o
    .io_cpu_decode_mmuRefilling            (IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling         ), //o
    .io_cpu_decode_mmuException            (IBusCachedPlugin_cache_io_cpu_decode_mmuException         ), //o
    .io_cpu_decode_isUser                  (IBusCachedPlugin_cache_io_cpu_decode_isUser               ), //i
    .io_cpu_fill_valid                     (IBusCachedPlugin_cache_io_cpu_fill_valid                  ), //i
    .io_cpu_fill_payload                   (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31:0]), //i
    .io_mem_cmd_valid                      (IBusCachedPlugin_cache_io_mem_cmd_valid                   ), //o
    .io_mem_cmd_ready                      (iBus_cmd_ready                                            ), //i
    .io_mem_cmd_payload_address            (IBusCachedPlugin_cache_io_mem_cmd_payload_address[31:0]   ), //o
    .io_mem_cmd_payload_size               (IBusCachedPlugin_cache_io_mem_cmd_payload_size[2:0]       ), //o
    .io_mem_rsp_valid                      (iBus_rsp_valid                                            ), //i
    .io_mem_rsp_payload_data               (iBus_rsp_payload_data[63:0]                               ), //i
    .io_mem_rsp_payload_error              (iBus_rsp_payload_error                                    ), //i
    .io_systemClk                          (io_systemClk                                              ), //i
    .systemCd_logic_outputReset            (systemCd_logic_outputReset                                )  //i
  );
  DataCache dataCache_2 (
    .io_cpu_execute_isValid                 (dataCache_2_io_cpu_execute_isValid               ), //i
    .io_cpu_execute_address                 (dataCache_2_io_cpu_execute_address[31:0]         ), //i
    .io_cpu_execute_haltIt                  (dataCache_2_io_cpu_execute_haltIt                ), //o
    .io_cpu_execute_args_wr                 (execute_MEMORY_WR                                ), //i
    .io_cpu_execute_args_size               (execute_DBusCachedPlugin_size[1:0]               ), //i
    .io_cpu_execute_args_isLrsc             (dataCache_2_io_cpu_execute_args_isLrsc           ), //i
    .io_cpu_execute_args_isAmo              (execute_MEMORY_AMO                               ), //i
    .io_cpu_execute_args_amoCtrl_swap       (dataCache_2_io_cpu_execute_args_amoCtrl_swap     ), //i
    .io_cpu_execute_args_amoCtrl_alu        (dataCache_2_io_cpu_execute_args_amoCtrl_alu[2:0] ), //i
    .io_cpu_execute_args_totalyConsistent   (execute_MEMORY_FORCE_CONSTISTENCY                ), //i
    .io_cpu_execute_refilling               (dataCache_2_io_cpu_execute_refilling             ), //o
    .io_cpu_memory_isValid                  (dataCache_2_io_cpu_memory_isValid                ), //i
    .io_cpu_memory_isStuck                  (memory_arbitration_isStuck                       ), //i
    .io_cpu_memory_isWrite                  (dataCache_2_io_cpu_memory_isWrite                ), //o
    .io_cpu_memory_address                  (memory_MEMORY_VIRTUAL_ADDRESS[31:0]              ), //i
    .io_cpu_memory_mmuRsp_physicalAddress   (DBusCachedPlugin_mmuBus_rsp_physicalAddress[31:0]), //i
    .io_cpu_memory_mmuRsp_isIoAccess        (dataCache_2_io_cpu_memory_mmuRsp_isIoAccess      ), //i
    .io_cpu_memory_mmuRsp_isPaging          (DBusCachedPlugin_mmuBus_rsp_isPaging             ), //i
    .io_cpu_memory_mmuRsp_allowRead         (DBusCachedPlugin_mmuBus_rsp_allowRead            ), //i
    .io_cpu_memory_mmuRsp_allowWrite        (DBusCachedPlugin_mmuBus_rsp_allowWrite           ), //i
    .io_cpu_memory_mmuRsp_allowExecute      (DBusCachedPlugin_mmuBus_rsp_allowExecute         ), //i
    .io_cpu_memory_mmuRsp_exception         (DBusCachedPlugin_mmuBus_rsp_exception            ), //i
    .io_cpu_memory_mmuRsp_refilling         (DBusCachedPlugin_mmuBus_rsp_refilling            ), //i
    .io_cpu_memory_mmuRsp_bypassTranslation (DBusCachedPlugin_mmuBus_rsp_bypassTranslation    ), //i
    .io_cpu_writeBack_isValid               (dataCache_2_io_cpu_writeBack_isValid             ), //i
    .io_cpu_writeBack_isStuck               (writeBack_arbitration_isStuck                    ), //i
    .io_cpu_writeBack_isFiring              (writeBack_arbitration_isFiring                   ), //i
    .io_cpu_writeBack_isUser                (dataCache_2_io_cpu_writeBack_isUser              ), //i
    .io_cpu_writeBack_haltIt                (dataCache_2_io_cpu_writeBack_haltIt              ), //o
    .io_cpu_writeBack_isWrite               (dataCache_2_io_cpu_writeBack_isWrite             ), //o
    .io_cpu_writeBack_storeData             (dataCache_2_io_cpu_writeBack_storeData[63:0]     ), //i
    .io_cpu_writeBack_data                  (dataCache_2_io_cpu_writeBack_data[63:0]          ), //o
    .io_cpu_writeBack_address               (dataCache_2_io_cpu_writeBack_address[31:0]       ), //i
    .io_cpu_writeBack_mmuException          (dataCache_2_io_cpu_writeBack_mmuException        ), //o
    .io_cpu_writeBack_unalignedAccess       (dataCache_2_io_cpu_writeBack_unalignedAccess     ), //o
    .io_cpu_writeBack_accessError           (dataCache_2_io_cpu_writeBack_accessError         ), //o
    .io_cpu_writeBack_keepMemRspData        (dataCache_2_io_cpu_writeBack_keepMemRspData      ), //o
    .io_cpu_writeBack_fence_SW              (dataCache_2_io_cpu_writeBack_fence_SW            ), //i
    .io_cpu_writeBack_fence_SR              (dataCache_2_io_cpu_writeBack_fence_SR            ), //i
    .io_cpu_writeBack_fence_SO              (dataCache_2_io_cpu_writeBack_fence_SO            ), //i
    .io_cpu_writeBack_fence_SI              (dataCache_2_io_cpu_writeBack_fence_SI            ), //i
    .io_cpu_writeBack_fence_PW              (dataCache_2_io_cpu_writeBack_fence_PW            ), //i
    .io_cpu_writeBack_fence_PR              (dataCache_2_io_cpu_writeBack_fence_PR            ), //i
    .io_cpu_writeBack_fence_PO              (dataCache_2_io_cpu_writeBack_fence_PO            ), //i
    .io_cpu_writeBack_fence_PI              (dataCache_2_io_cpu_writeBack_fence_PI            ), //i
    .io_cpu_writeBack_fence_FM              (dataCache_2_io_cpu_writeBack_fence_FM[3:0]       ), //i
    .io_cpu_writeBack_exclusiveOk           (dataCache_2_io_cpu_writeBack_exclusiveOk         ), //o
    .io_cpu_redo                            (dataCache_2_io_cpu_redo                          ), //o
    .io_cpu_flush_valid                     (dataCache_2_io_cpu_flush_valid                   ), //i
    .io_cpu_flush_ready                     (dataCache_2_io_cpu_flush_ready                   ), //o
    .io_cpu_flush_payload_singleLine        (dataCache_2_io_cpu_flush_payload_singleLine      ), //i
    .io_cpu_flush_payload_lineId            (dataCache_2_io_cpu_flush_payload_lineId[5:0]     ), //i
    .io_cpu_writesPending                   (dataCache_2_io_cpu_writesPending                 ), //o
    .io_mem_cmd_valid                       (dataCache_2_io_mem_cmd_valid                     ), //o
    .io_mem_cmd_ready                       (dataCache_2_io_mem_cmd_rValidN                   ), //i
    .io_mem_cmd_payload_wr                  (dataCache_2_io_mem_cmd_payload_wr                ), //o
    .io_mem_cmd_payload_uncached            (dataCache_2_io_mem_cmd_payload_uncached          ), //o
    .io_mem_cmd_payload_address             (dataCache_2_io_mem_cmd_payload_address[31:0]     ), //o
    .io_mem_cmd_payload_data                (dataCache_2_io_mem_cmd_payload_data[63:0]        ), //o
    .io_mem_cmd_payload_mask                (dataCache_2_io_mem_cmd_payload_mask[7:0]         ), //o
    .io_mem_cmd_payload_size                (dataCache_2_io_mem_cmd_payload_size[2:0]         ), //o
    .io_mem_cmd_payload_exclusive           (dataCache_2_io_mem_cmd_payload_exclusive         ), //o
    .io_mem_cmd_payload_last                (dataCache_2_io_mem_cmd_payload_last              ), //o
    .io_mem_rsp_valid                       (dBus_rsp_valid_regNext                           ), //i
    .io_mem_rsp_payload_aggregated          (dBus_rsp_payload_aggregated_regNext[3:0]         ), //i
    .io_mem_rsp_payload_last                (dBus_rsp_payload_last_regNext                    ), //i
    .io_mem_rsp_payload_data                (dBus_rsp_payload_data_regNextWhen[63:0]          ), //i
    .io_mem_rsp_payload_error               (dBus_rsp_payload_error_regNext                   ), //i
    .io_mem_rsp_payload_exclusive           (dBus_rsp_payload_exclusive_regNext               ), //i
    .io_mem_inv_valid                       (dBus_inv_valid                                   ), //i
    .io_mem_inv_ready                       (dataCache_2_io_mem_inv_ready                     ), //o
    .io_mem_inv_payload_last                (dBus_inv_payload_last                            ), //i
    .io_mem_inv_payload_fragment_enable     (dBus_inv_payload_fragment_enable                 ), //i
    .io_mem_inv_payload_fragment_address    (dBus_inv_payload_fragment_address[31:0]          ), //i
    .io_mem_ack_valid                       (dataCache_2_io_mem_ack_valid                     ), //o
    .io_mem_ack_ready                       (dBus_ack_ready                                   ), //i
    .io_mem_ack_payload_last                (dataCache_2_io_mem_ack_payload_last              ), //o
    .io_mem_ack_payload_fragment_hit        (dataCache_2_io_mem_ack_payload_fragment_hit      ), //o
    .io_mem_sync_valid                      (dBus_sync_valid                                  ), //i
    .io_mem_sync_ready                      (dataCache_2_io_mem_sync_ready                    ), //o
    .io_mem_sync_payload_aggregated         (dBus_sync_payload_aggregated[3:0]                ), //i
    .io_systemClk                           (io_systemClk                                     ), //i
    .systemCd_logic_outputReset             (systemCd_logic_outputReset                       )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC systemCd_logic_outputReset_buffercc (
    .io_dataIn                  (systemCd_logic_outputReset                    ), //i
    .io_dataOut                 (systemCd_logic_outputReset_buffercc_io_dataOut), //o
    .io_systemClk               (io_systemClk                                  ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                    )  //i
  );
  EfxCPUSp1 EfxCPUSp1_inst (
    .src1    (execute_SRC1[31:0]           ), //i
    .src2    (execute_SRC2[31:0]           ), //i
    .bitCtrl (execute_ALU_BITWISE_CTRL[1:0]), //i
    .ctrl    (execute_ALU_CTRL[1:0]        ), //i
    .less    (execute_SRC_LESS             ), //i
    .addSub  (execute_SRC_ADD_SUB[31:0]    ), //i
    .result  (EfxCPUSp1_inst_result[31:0]  )  //o
  );
  EfxCPUSp2 EfxCPUSp2_inst (
    .ctrl   (execute_SHIFT_CTRL[1:0]    ), //i
    .src1   (execute_SRC1[31:0]         ), //i
    .src2   (execute_SRC2[31:0]         ), //i
    .result (EfxCPUSp2_inst_result[31:0])  //o
  );
  always @(*) begin
    case(_zz_IBusCachedPlugin_jump_pcLoad_payload_5)
      2'b00 : _zz_IBusCachedPlugin_jump_pcLoad_payload_4 = DBusCachedPlugin_redoBranch_payload;
      2'b01 : _zz_IBusCachedPlugin_jump_pcLoad_payload_4 = CsrPlugin_jumpInterface_payload;
      default : _zz_IBusCachedPlugin_jump_pcLoad_payload_4 = BranchPlugin_jumpInterface_payload;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_1)
      3'b000 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_0;
      3'b001 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_1;
      3'b010 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_2;
      3'b011 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_3;
      3'b100 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_4;
      3'b101 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_5;
      3'b110 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_6;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_7;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_3)
      2'b00 : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_1;
      2'b01 : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_3;
      2'b10 : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_5;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_7;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_5)
      1'b0 : _zz_writeBack_DBusCachedPlugin_rspShifted_4 = writeBack_DBusCachedPlugin_rspSplits_2;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted_4 = writeBack_DBusCachedPlugin_rspSplits_6;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_7)
      1'b0 : _zz_writeBack_DBusCachedPlugin_rspShifted_6 = writeBack_DBusCachedPlugin_rspSplits_3;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted_6 = writeBack_DBusCachedPlugin_rspSplits_7;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(_zz_execute_to_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_execute_to_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_execute_to_memory_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : decode_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : decode_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : decode_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : decode_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : decode_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL_1)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : decode_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : decode_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : decode_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1)
      Input2Kind_RS : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string = "IMM_I";
      default : _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(memory_FPU_OPCODE)
      FpuOpcode_LOAD : memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : memory_FPU_OPCODE_string = "FCVT_X_X";
      default : memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_memory_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_memory_to_writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_memory_to_writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_memory_to_writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_memory_to_writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_memory_to_writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_memory_to_writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_memory_to_writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_memory_to_writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_memory_to_writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_memory_to_writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_memory_to_writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_memory_to_writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_memory_to_writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_memory_to_writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_memory_to_writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_memory_to_writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_memory_to_writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_memory_to_writeBack_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_FPU_OPCODE)
      FpuOpcode_LOAD : execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : execute_FPU_OPCODE_string = "FCVT_X_X";
      default : execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_execute_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_execute_to_memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_execute_to_memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_execute_to_memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_execute_to_memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_execute_to_memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_execute_to_memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_execute_to_memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_execute_to_memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_execute_to_memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_execute_to_memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_execute_to_memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_execute_to_memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_execute_to_memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_execute_to_memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_execute_to_memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_execute_to_memory_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_execute_to_memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_execute_to_memory_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_execute_to_memory_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_execute_to_memory_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_execute_to_memory_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_execute_to_memory_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_execute_to_memory_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_execute_to_memory_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_execute_to_memory_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_execute_to_memory_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_execute_to_memory_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_execute_to_memory_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_execute_to_memory_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_execute_to_memory_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_execute_to_memory_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_execute_to_memory_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_execute_to_memory_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_execute_to_memory_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_decode_to_execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_to_execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_to_execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_to_execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_to_execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_to_execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_to_execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_to_execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_to_execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_to_execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_to_execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_to_execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_to_execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_to_execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_to_execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_to_execute_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_decode_to_execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_decode_to_execute_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_to_execute_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_to_execute_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_to_execute_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_to_execute_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_to_execute_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_to_execute_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_to_execute_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_to_execute_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_to_execute_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_to_execute_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_to_execute_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_to_execute_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_to_execute_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_to_execute_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_to_execute_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_decode_to_execute_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_BRANCH_CTRL)
      BranchCtrlEnum_INC : decode_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : decode_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : decode_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : decode_BRANCH_CTRL_string = "JALR";
      default : decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_decode_to_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_to_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_to_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL_1)
      BranchCtrlEnum_INC : _zz_decode_to_execute_BRANCH_CTRL_1_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_to_execute_BRANCH_CTRL_1_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_memory_to_writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_memory_to_writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_memory_to_writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_memory_to_writeBack_ENV_CTRL_string = "EBREAK";
      default : _zz_memory_to_writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_memory_to_writeBack_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_memory_to_writeBack_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_memory_to_writeBack_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_memory_to_writeBack_ENV_CTRL_1_string = "EBREAK";
      default : _zz_memory_to_writeBack_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_execute_to_memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_execute_to_memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_execute_to_memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_execute_to_memory_ENV_CTRL_string = "EBREAK";
      default : _zz_execute_to_memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_execute_to_memory_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_execute_to_memory_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_execute_to_memory_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_execute_to_memory_ENV_CTRL_1_string = "EBREAK";
      default : _zz_execute_to_memory_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_ENV_CTRL)
      EnvCtrlEnum_NONE : decode_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : decode_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : decode_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : decode_ENV_CTRL_string = "EBREAK";
      default : decode_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_ENV_CTRL_string = "EBREAK";
      default : _zz_decode_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_decode_to_execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_to_execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_to_execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_to_execute_ENV_CTRL_string = "EBREAK";
      default : _zz_decode_to_execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_decode_to_execute_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_to_execute_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_to_execute_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_to_execute_ENV_CTRL_1_string = "EBREAK";
      default : _zz_decode_to_execute_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : decode_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : decode_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : decode_ALU_CTRL_string = "BITWISE ";
      default : decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL_1)
      AluCtrlEnum_ADD_SUB : _zz_decode_to_execute_ALU_CTRL_1_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_to_execute_ALU_CTRL_1_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_to_execute_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : memory_SHIFT_CTRL_string = "SRA_1    ";
      default : memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : execute_SHIFT_CTRL_string = "SRA_1    ";
      default : execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : execute_ALU_CTRL_string = "BITWISE ";
      default : execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : _zz_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_FPU_FORMAT)
      FpuFormat_FLOAT : decode_FPU_FORMAT_string = "FLOAT ";
      FpuFormat_DOUBLE : decode_FPU_FORMAT_string = "DOUBLE";
      default : decode_FPU_FORMAT_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_FORMAT)
      FpuFormat_FLOAT : _zz_decode_FPU_FORMAT_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_decode_FPU_FORMAT_string = "DOUBLE";
      default : _zz_decode_FPU_FORMAT_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_FPU_OPCODE)
      FpuOpcode_LOAD : decode_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : decode_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : decode_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : decode_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : decode_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : decode_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : decode_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : decode_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : decode_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : decode_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : decode_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : decode_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : decode_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : decode_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : decode_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : decode_FPU_OPCODE_string = "FCVT_X_X";
      default : decode_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_OPCODE)
      FpuOpcode_LOAD : _zz_decode_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_FPU_OPCODE_string = "FCVT_X_X";
      default : _zz_decode_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : execute_BRANCH_CTRL_string = "JALR";
      default : execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(memory_ENV_CTRL)
      EnvCtrlEnum_NONE : memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : memory_ENV_CTRL_string = "EBREAK";
      default : memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_memory_ENV_CTRL_string = "EBREAK";
      default : _zz_memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_ENV_CTRL)
      EnvCtrlEnum_NONE : execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : execute_ENV_CTRL_string = "EBREAK";
      default : execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_execute_ENV_CTRL_string = "EBREAK";
      default : _zz_execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : writeBack_ENV_CTRL_string = "EBREAK";
      default : writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_writeBack_ENV_CTRL_string = "EBREAK";
      default : _zz_writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_SRC2_CTRL)
      Src2CtrlEnum_RS : decode_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : decode_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : decode_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : decode_SRC2_CTRL_string = "PC ";
      default : decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_string = "PC ";
      default : _zz_decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_SRC1_CTRL)
      Src1CtrlEnum_RS : decode_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : decode_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : decode_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : decode_SRC1_CTRL_string = "URS1        ";
      default : decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_1)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1)
      Input2Kind_RS : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string = "IMM_I";
      default : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_FORMAT_1)
      FpuFormat_FLOAT : _zz_decode_FPU_FORMAT_1_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_decode_FPU_FORMAT_1_string = "DOUBLE";
      default : _zz_decode_FPU_FORMAT_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_OPCODE_1)
      FpuOpcode_LOAD : _zz_decode_FPU_OPCODE_1_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_FPU_OPCODE_1_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_FPU_OPCODE_1_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_FPU_OPCODE_1_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_FPU_OPCODE_1_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_FPU_OPCODE_1_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_FPU_OPCODE_1_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_FPU_OPCODE_1_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_FPU_OPCODE_1_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_FPU_OPCODE_1_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_FPU_OPCODE_1_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_FPU_OPCODE_1_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_FPU_OPCODE_1_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_FPU_OPCODE_1_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_FPU_OPCODE_1_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_FPU_OPCODE_1_string = "FCVT_X_X";
      default : _zz_decode_FPU_OPCODE_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_1)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_1_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_1_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_1_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_1_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_1_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_1_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_ENV_CTRL_1_string = "EBREAK";
      default : _zz_decode_ENV_CTRL_1_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_1)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_1_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_1_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_1_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_1_string = "PC ";
      default : _zz_decode_SRC2_CTRL_1_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_1)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_1_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_1_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_1)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_1_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_1_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_1_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_1_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_1_string = "????????????";
    endcase
  end
  always @(*) begin
    case(debugBus_dmToHart_payload_op)
      DebugDmToHartOp_DATA : debugBus_dmToHart_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : debugBus_dmToHart_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : debugBus_dmToHart_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : debugBus_dmToHart_payload_op_string = "REG_READ ";
      default : debugBus_dmToHart_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_cmd_payload_opcode)
      FpuOpcode_LOAD : FpuPlugin_port_cmd_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_cmd_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_cmd_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_cmd_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_cmd_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_cmd_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_cmd_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_cmd_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_cmd_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_cmd_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_cmd_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_cmd_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_cmd_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_cmd_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_cmd_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_cmd_payload_opcode_string = "FCVT_X_X";
      default : FpuPlugin_port_cmd_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_cmd_payload_format)
      FpuFormat_FLOAT : FpuPlugin_port_cmd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : FpuPlugin_port_cmd_payload_format_string = "DOUBLE";
      default : FpuPlugin_port_cmd_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_cmd_payload_roundMode)
      FpuRoundMode_RNE : FpuPlugin_port_cmd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : FpuPlugin_port_cmd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : FpuPlugin_port_cmd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : FpuPlugin_port_cmd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : FpuPlugin_port_cmd_payload_roundMode_string = "RMM";
      default : FpuPlugin_port_cmd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_port_commit_payload_opcode)
      FpuOpcode_LOAD : FpuPlugin_port_commit_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : FpuPlugin_port_commit_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : FpuPlugin_port_commit_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : FpuPlugin_port_commit_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : FpuPlugin_port_commit_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : FpuPlugin_port_commit_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : FpuPlugin_port_commit_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : FpuPlugin_port_commit_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : FpuPlugin_port_commit_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : FpuPlugin_port_commit_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : FpuPlugin_port_commit_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : FpuPlugin_port_commit_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : FpuPlugin_port_commit_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : FpuPlugin_port_commit_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : FpuPlugin_port_commit_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : FpuPlugin_port_commit_payload_opcode_string = "FCVT_X_X";
      default : FpuPlugin_port_commit_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_2)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_2_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_2_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_2_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_2_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_2_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_2)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_2_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_2_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_2_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_2)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_2_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_2_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_2_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_2_string = "PC ";
      default : _zz_decode_SRC2_CTRL_2_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_2)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_2_string = "NONE  ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_2_string = "XRET  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_2_string = "ECALL ";
      EnvCtrlEnum_EBREAK : _zz_decode_ENV_CTRL_2_string = "EBREAK";
      default : _zz_decode_ENV_CTRL_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_2)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_2_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_2_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_2_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_2_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_OPCODE_2)
      FpuOpcode_LOAD : _zz_decode_FPU_OPCODE_2_string = "LOAD    ";
      FpuOpcode_STORE : _zz_decode_FPU_OPCODE_2_string = "STORE   ";
      FpuOpcode_MUL : _zz_decode_FPU_OPCODE_2_string = "MUL     ";
      FpuOpcode_ADD : _zz_decode_FPU_OPCODE_2_string = "ADD     ";
      FpuOpcode_FMA : _zz_decode_FPU_OPCODE_2_string = "FMA     ";
      FpuOpcode_I2F : _zz_decode_FPU_OPCODE_2_string = "I2F     ";
      FpuOpcode_F2I : _zz_decode_FPU_OPCODE_2_string = "F2I     ";
      FpuOpcode_CMP : _zz_decode_FPU_OPCODE_2_string = "CMP     ";
      FpuOpcode_DIV : _zz_decode_FPU_OPCODE_2_string = "DIV     ";
      FpuOpcode_SQRT : _zz_decode_FPU_OPCODE_2_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_decode_FPU_OPCODE_2_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_decode_FPU_OPCODE_2_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_decode_FPU_OPCODE_2_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_decode_FPU_OPCODE_2_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_decode_FPU_OPCODE_2_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_decode_FPU_OPCODE_2_string = "FCVT_X_X";
      default : _zz_decode_FPU_OPCODE_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_FPU_FORMAT_2)
      FpuFormat_FLOAT : _zz_decode_FPU_FORMAT_2_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_decode_FPU_FORMAT_2_string = "DOUBLE";
      default : _zz_decode_FPU_FORMAT_2_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2)
      Input2Kind_RS : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string = "RS   ";
      Input2Kind_IMM_I : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string = "IMM_I";
      default : _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_2)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_2)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_2_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_2_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_2_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_2_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_2_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_cmd_payload_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_cmd_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_cmd_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_cmd_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_cmd_payload_op_string = "REG_READ ";
      default : CsrPlugin_inject_cmd_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_cmd_toStream_payload_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_cmd_toStream_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_cmd_toStream_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_cmd_toStream_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_cmd_toStream_payload_op_string = "REG_READ ";
      default : CsrPlugin_inject_cmd_toStream_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_buffer_payload_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_buffer_payload_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_buffer_payload_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_buffer_payload_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_buffer_payload_op_string = "REG_READ ";
      default : CsrPlugin_inject_buffer_payload_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_inject_cmd_toStream_rData_op)
      DebugDmToHartOp_DATA : CsrPlugin_inject_cmd_toStream_rData_op_string = "DATA     ";
      DebugDmToHartOp_EXECUTE : CsrPlugin_inject_cmd_toStream_rData_op_string = "EXECUTE  ";
      DebugDmToHartOp_REG_WRITE : CsrPlugin_inject_cmd_toStream_rData_op_string = "REG_WRITE";
      DebugDmToHartOp_REG_READ : CsrPlugin_inject_cmd_toStream_rData_op_string = "REG_READ ";
      default : CsrPlugin_inject_cmd_toStream_rData_op_string = "?????????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_BOOT : CsrPlugin_dcsr_stepLogic_stateReg_string = "BOOT  ";
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : CsrPlugin_dcsr_stepLogic_stateReg_string = "IDLE  ";
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : CsrPlugin_dcsr_stepLogic_stateReg_string = "SINGLE";
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : CsrPlugin_dcsr_stepLogic_stateReg_string = "WAIT_1";
      default : CsrPlugin_dcsr_stepLogic_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(CsrPlugin_dcsr_stepLogic_stateNext)
      CsrPlugin_dcsr_stepLogic_enumDef_BOOT : CsrPlugin_dcsr_stepLogic_stateNext_string = "BOOT  ";
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : CsrPlugin_dcsr_stepLogic_stateNext_string = "IDLE  ";
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : CsrPlugin_dcsr_stepLogic_stateNext_string = "SINGLE";
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : CsrPlugin_dcsr_stepLogic_stateNext_string = "WAIT_1";
      default : CsrPlugin_dcsr_stepLogic_stateNext_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPlugin_port_cmd_payload_roundMode)
      FpuRoundMode_RNE : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "RMM";
      default : _zz_FpuPlugin_port_cmd_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPlugin_port_cmd_payload_roundMode_1)
      FpuRoundMode_RNE : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RNE";
      FpuRoundMode_RTZ : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RTZ";
      FpuRoundMode_RDN : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RDN";
      FpuRoundMode_RUP : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RUP";
      FpuRoundMode_RMM : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "RMM";
      default : _zz_FpuPlugin_port_cmd_payload_roundMode_1_string = "???";
    endcase
  end
  always @(*) begin
    case(writeBack_FpuPlugin_commit_payload_opcode)
      FpuOpcode_LOAD : writeBack_FpuPlugin_commit_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FpuPlugin_commit_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FpuPlugin_commit_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FpuPlugin_commit_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FpuPlugin_commit_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FpuPlugin_commit_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FpuPlugin_commit_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FpuPlugin_commit_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FpuPlugin_commit_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FpuPlugin_commit_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FpuPlugin_commit_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FpuPlugin_commit_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FpuPlugin_commit_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FpuPlugin_commit_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FpuPlugin_commit_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FpuPlugin_commit_payload_opcode_string = "FCVT_X_X";
      default : writeBack_FpuPlugin_commit_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(writeBack_FpuPlugin_commit_s2mPipe_payload_opcode)
      FpuOpcode_LOAD : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCVT_X_X";
      default : writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(writeBack_FpuPlugin_commit_rData_opcode)
      FpuOpcode_LOAD : writeBack_FpuPlugin_commit_rData_opcode_string = "LOAD    ";
      FpuOpcode_STORE : writeBack_FpuPlugin_commit_rData_opcode_string = "STORE   ";
      FpuOpcode_MUL : writeBack_FpuPlugin_commit_rData_opcode_string = "MUL     ";
      FpuOpcode_ADD : writeBack_FpuPlugin_commit_rData_opcode_string = "ADD     ";
      FpuOpcode_FMA : writeBack_FpuPlugin_commit_rData_opcode_string = "FMA     ";
      FpuOpcode_I2F : writeBack_FpuPlugin_commit_rData_opcode_string = "I2F     ";
      FpuOpcode_F2I : writeBack_FpuPlugin_commit_rData_opcode_string = "F2I     ";
      FpuOpcode_CMP : writeBack_FpuPlugin_commit_rData_opcode_string = "CMP     ";
      FpuOpcode_DIV : writeBack_FpuPlugin_commit_rData_opcode_string = "DIV     ";
      FpuOpcode_SQRT : writeBack_FpuPlugin_commit_rData_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : writeBack_FpuPlugin_commit_rData_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : writeBack_FpuPlugin_commit_rData_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : writeBack_FpuPlugin_commit_rData_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : writeBack_FpuPlugin_commit_rData_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : writeBack_FpuPlugin_commit_rData_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : writeBack_FpuPlugin_commit_rData_opcode_string = "FCVT_X_X";
      default : writeBack_FpuPlugin_commit_rData_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode)
      FpuOpcode_LOAD : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "FCVT_X_X";
      default : _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : decode_to_execute_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : decode_to_execute_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : decode_to_execute_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : decode_to_execute_ENV_CTRL_string = "EBREAK";
      default : decode_to_execute_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : execute_to_memory_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : execute_to_memory_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : execute_to_memory_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : execute_to_memory_ENV_CTRL_string = "EBREAK";
      default : execute_to_memory_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(memory_to_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : memory_to_writeBack_ENV_CTRL_string = "NONE  ";
      EnvCtrlEnum_XRET : memory_to_writeBack_ENV_CTRL_string = "XRET  ";
      EnvCtrlEnum_ECALL : memory_to_writeBack_ENV_CTRL_string = "ECALL ";
      EnvCtrlEnum_EBREAK : memory_to_writeBack_ENV_CTRL_string = "EBREAK";
      default : memory_to_writeBack_ENV_CTRL_string = "??????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : decode_to_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : decode_to_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : decode_to_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_FPU_OPCODE)
      FpuOpcode_LOAD : decode_to_execute_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : decode_to_execute_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : decode_to_execute_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : decode_to_execute_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : decode_to_execute_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : decode_to_execute_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : decode_to_execute_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : decode_to_execute_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : decode_to_execute_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : decode_to_execute_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : decode_to_execute_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : decode_to_execute_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : decode_to_execute_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : decode_to_execute_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : decode_to_execute_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : decode_to_execute_FPU_OPCODE_string = "FCVT_X_X";
      default : decode_to_execute_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_FPU_OPCODE)
      FpuOpcode_LOAD : execute_to_memory_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : execute_to_memory_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : execute_to_memory_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : execute_to_memory_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : execute_to_memory_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : execute_to_memory_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : execute_to_memory_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : execute_to_memory_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : execute_to_memory_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : execute_to_memory_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : execute_to_memory_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : execute_to_memory_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : execute_to_memory_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : execute_to_memory_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : execute_to_memory_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : execute_to_memory_FPU_OPCODE_string = "FCVT_X_X";
      default : execute_to_memory_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(memory_to_writeBack_FPU_OPCODE)
      FpuOpcode_LOAD : memory_to_writeBack_FPU_OPCODE_string = "LOAD    ";
      FpuOpcode_STORE : memory_to_writeBack_FPU_OPCODE_string = "STORE   ";
      FpuOpcode_MUL : memory_to_writeBack_FPU_OPCODE_string = "MUL     ";
      FpuOpcode_ADD : memory_to_writeBack_FPU_OPCODE_string = "ADD     ";
      FpuOpcode_FMA : memory_to_writeBack_FPU_OPCODE_string = "FMA     ";
      FpuOpcode_I2F : memory_to_writeBack_FPU_OPCODE_string = "I2F     ";
      FpuOpcode_F2I : memory_to_writeBack_FPU_OPCODE_string = "F2I     ";
      FpuOpcode_CMP : memory_to_writeBack_FPU_OPCODE_string = "CMP     ";
      FpuOpcode_DIV : memory_to_writeBack_FPU_OPCODE_string = "DIV     ";
      FpuOpcode_SQRT : memory_to_writeBack_FPU_OPCODE_string = "SQRT    ";
      FpuOpcode_MIN_MAX : memory_to_writeBack_FPU_OPCODE_string = "MIN_MAX ";
      FpuOpcode_SGNJ : memory_to_writeBack_FPU_OPCODE_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : memory_to_writeBack_FPU_OPCODE_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : memory_to_writeBack_FPU_OPCODE_string = "FMV_W_X ";
      FpuOpcode_FCLASS : memory_to_writeBack_FPU_OPCODE_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : memory_to_writeBack_FPU_OPCODE_string = "FCVT_X_X";
      default : memory_to_writeBack_FPU_OPCODE_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "RS   ";
      Input2Kind_IMM_I : decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "IMM_I";
      default : decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : execute_to_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : execute_to_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : execute_to_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : execute_to_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : execute_to_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_BOOT : FpuPlugin_stateReg_string = "BOOT  ";
      FpuPlugin_enumDef_IDLE : FpuPlugin_stateReg_string = "IDLE  ";
      FpuPlugin_enumDef_CMD : FpuPlugin_stateReg_string = "CMD   ";
      FpuPlugin_enumDef_RSP : FpuPlugin_stateReg_string = "RSP   ";
      FpuPlugin_enumDef_RSP_0 : FpuPlugin_stateReg_string = "RSP_0 ";
      FpuPlugin_enumDef_RSP_1 : FpuPlugin_stateReg_string = "RSP_1 ";
      FpuPlugin_enumDef_COMMIT : FpuPlugin_stateReg_string = "COMMIT";
      FpuPlugin_enumDef_DONE : FpuPlugin_stateReg_string = "DONE  ";
      default : FpuPlugin_stateReg_string = "??????";
    endcase
  end
  always @(*) begin
    case(FpuPlugin_stateNext)
      FpuPlugin_enumDef_BOOT : FpuPlugin_stateNext_string = "BOOT  ";
      FpuPlugin_enumDef_IDLE : FpuPlugin_stateNext_string = "IDLE  ";
      FpuPlugin_enumDef_CMD : FpuPlugin_stateNext_string = "CMD   ";
      FpuPlugin_enumDef_RSP : FpuPlugin_stateNext_string = "RSP   ";
      FpuPlugin_enumDef_RSP_0 : FpuPlugin_stateNext_string = "RSP_0 ";
      FpuPlugin_enumDef_RSP_1 : FpuPlugin_stateNext_string = "RSP_1 ";
      FpuPlugin_enumDef_COMMIT : FpuPlugin_stateNext_string = "COMMIT";
      FpuPlugin_enumDef_DONE : FpuPlugin_stateNext_string = "DONE  ";
      default : FpuPlugin_stateNext_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_FpuPlugin_port_cmd_payload_format)
      FpuFormat_FLOAT : _zz_FpuPlugin_port_cmd_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_FpuPlugin_port_cmd_payload_format_string = "DOUBLE";
      default : _zz_FpuPlugin_port_cmd_payload_format_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    CsrPlugin_running_aheadValue = CsrPlugin_running;
    if(when_CsrPlugin_l1534) begin
      if(!when_CsrPlugin_l1542) begin
        CsrPlugin_running_aheadValue = 1'b0;
      end
    end
    if(CsrPlugin_doResume) begin
      CsrPlugin_running_aheadValue = 1'b1;
    end
  end

  assign writeBack_MEMORY_LOAD_DATA = writeBack_DBusCachedPlugin_rspShifted;
  assign memory_MUL_LOW = ($signed(_zz_memory_MUL_LOW) + $signed(_zz_memory_MUL_LOW_6));
  assign execute_SHIFT_RIGHT = EfxCPUSp2_inst_result;
  assign execute_REGFILE_WRITE_DATA = EfxCPUSp1_inst_result;
  assign memory_CfuPlugin_CFU_IN_FLIGHT = execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
  assign execute_CfuPlugin_CFU_IN_FLIGHT = ((execute_CfuPlugin_schedule || execute_CfuPlugin_hold) || execute_CfuPlugin_fired);
  assign memory_MUL_HH = execute_to_memory_MUL_HH;
  assign execute_MUL_HH = execute_MulPlugin_withOuputBuffer_mul_hh;
  assign execute_MUL_HL = execute_MulPlugin_withOuputBuffer_mul_hl;
  assign execute_MUL_LH = execute_MulPlugin_withOuputBuffer_mul_lh;
  assign execute_MUL_LL = execute_MulPlugin_withOuputBuffer_mul_ll;
  assign execute_BRANCH_CALC = {execute_BranchPlugin_branchAdder[31 : 1],1'b0};
  assign execute_BRANCH_DO = _zz_execute_BRANCH_DO_1;
  assign execute_MEMORY_VIRTUAL_ADDRESS = dataCache_2_io_cpu_execute_address;
  assign execute_MEMORY_STORE_DATA_RF = _zz_execute_MEMORY_STORE_DATA_RF;
  assign memory_FPU_COMMIT_LOAD = execute_to_memory_FPU_COMMIT_LOAD;
  assign execute_FPU_COMMIT_LOAD = decode_to_execute_FPU_COMMIT_LOAD;
  assign decode_FPU_COMMIT_LOAD = (decode_FPU_OPCODE == FpuOpcode_LOAD);
  assign memory_FPU_FORKED = execute_to_memory_FPU_FORKED;
  assign execute_FPU_FORKED = decode_to_execute_FPU_FORKED;
  assign decode_FPU_FORKED = (decode_FpuPlugin_forked || (FpuPlugin_port_cmd_fire && (! _zz_decode_FPU_FORKED)));
  assign decode_CSR_READ_OPCODE = (decode_INSTRUCTION[13 : 7] != 7'h20);
  assign decode_CSR_WRITE_OPCODE = (! (((decode_INSTRUCTION[14 : 13] == 2'b01) && (decode_INSTRUCTION[19 : 15] == 5'h0)) || ((decode_INSTRUCTION[14 : 13] == 2'b11) && (decode_INSTRUCTION[19 : 15] == 5'h0))));
  assign decode_SRC2 = _zz_decode_SRC2_4;
  assign decode_SRC1 = _zz_decode_SRC1;
  assign decode_SRC2_FORCE_ZERO = (decode_SRC_ADD_ZERO && (! decode_SRC_USE_SUB_LESS));
  assign memory_RS1 = execute_to_memory_RS1;
  assign _zz_execute_to_memory_SHIFT_CTRL = _zz_execute_to_memory_SHIFT_CTRL_1;
  assign decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL = _zz_decode_to_execute_SHIFT_CTRL_1;
  assign decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL = _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  assign decode_CfuPlugin_CFU_INPUT_2_KIND = _zz_decode_CfuPlugin_CFU_INPUT_2_KIND;
  assign _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND = _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1;
  assign decode_CfuPlugin_CFU_ENABLE = _zz_decode_CfuPlugin_CFU_ENABLE[42];
  assign memory_FPU_OPCODE = _zz_memory_FPU_OPCODE;
  assign _zz_memory_to_writeBack_FPU_OPCODE = _zz_memory_to_writeBack_FPU_OPCODE_1;
  assign execute_FPU_OPCODE = _zz_execute_FPU_OPCODE;
  assign _zz_execute_to_memory_FPU_OPCODE = _zz_execute_to_memory_FPU_OPCODE_1;
  assign _zz_decode_to_execute_FPU_OPCODE = _zz_decode_to_execute_FPU_OPCODE_1;
  assign memory_FPU_RSP = execute_to_memory_FPU_RSP;
  assign execute_FPU_RSP = decode_to_execute_FPU_RSP;
  assign decode_FPU_RSP = _zz_decode_CfuPlugin_CFU_ENABLE[34];
  assign memory_FPU_COMMIT = execute_to_memory_FPU_COMMIT;
  assign execute_FPU_COMMIT = decode_to_execute_FPU_COMMIT;
  assign decode_FPU_COMMIT = _zz_decode_CfuPlugin_CFU_ENABLE[33];
  assign decode_IS_RS2_SIGNED = _zz_decode_CfuPlugin_CFU_ENABLE[31];
  assign decode_IS_RS1_SIGNED = _zz_decode_CfuPlugin_CFU_ENABLE[30];
  assign decode_IS_DIV = _zz_decode_CfuPlugin_CFU_ENABLE[29];
  assign memory_IS_MUL = execute_to_memory_IS_MUL;
  assign decode_IS_MUL = _zz_decode_CfuPlugin_CFU_ENABLE[28];
  assign decode_SRC_LESS_UNSIGNED = _zz_decode_CfuPlugin_CFU_ENABLE[27];
  assign decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL = _zz_decode_to_execute_BRANCH_CTRL_1;
  assign _zz_memory_to_writeBack_ENV_CTRL = _zz_memory_to_writeBack_ENV_CTRL_1;
  assign _zz_execute_to_memory_ENV_CTRL = _zz_execute_to_memory_ENV_CTRL_1;
  assign decode_ENV_CTRL = _zz_decode_ENV_CTRL;
  assign _zz_decode_to_execute_ENV_CTRL = _zz_decode_to_execute_ENV_CTRL_1;
  assign decode_IS_CSR = _zz_decode_CfuPlugin_CFU_ENABLE[22];
  assign memory_MEMORY_FENCE = execute_to_memory_MEMORY_FENCE;
  assign execute_MEMORY_FENCE = decode_to_execute_MEMORY_FENCE;
  assign decode_MEMORY_FENCE = _zz_decode_CfuPlugin_CFU_ENABLE[21];
  assign decode_MEMORY_MANAGMENT = _zz_decode_CfuPlugin_CFU_ENABLE[20];
  assign memory_MEMORY_AMO = execute_to_memory_MEMORY_AMO;
  assign memory_MEMORY_LRSC = execute_to_memory_MEMORY_LRSC;
  assign execute_HAS_SIDE_EFFECT = decode_to_execute_HAS_SIDE_EFFECT;
  assign decode_HAS_SIDE_EFFECT = _zz_decode_CfuPlugin_CFU_ENABLE[15];
  assign decode_MEMORY_WR = _zz_decode_CfuPlugin_CFU_ENABLE[14];
  assign execute_BYPASSABLE_MEMORY_STAGE = decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  assign decode_BYPASSABLE_MEMORY_STAGE = _zz_decode_CfuPlugin_CFU_ENABLE[13];
  assign decode_BYPASSABLE_EXECUTE_STAGE = _zz_decode_CfuPlugin_CFU_ENABLE[12];
  assign decode_ALU_CTRL = _zz_decode_ALU_CTRL;
  assign _zz_decode_to_execute_ALU_CTRL = _zz_decode_to_execute_ALU_CTRL_1;
  assign decode_MEMORY_FENCE_WR = _zz_decode_CfuPlugin_CFU_ENABLE[1];
  assign decode_MEMORY_FORCE_CONSTISTENCY = _zz_decode_MEMORY_FORCE_CONSTISTENCY;
  assign writeBack_FORMAL_PC_NEXT = memory_to_writeBack_FORMAL_PC_NEXT;
  assign memory_FORMAL_PC_NEXT = execute_to_memory_FORMAL_PC_NEXT;
  assign execute_FORMAL_PC_NEXT = decode_to_execute_FORMAL_PC_NEXT;
  assign decode_FORMAL_PC_NEXT = (decode_PC + _zz_decode_FORMAL_PC_NEXT);
  assign memory_SHIFT_RIGHT = execute_to_memory_SHIFT_RIGHT;
  assign memory_SHIFT_CTRL = _zz_memory_SHIFT_CTRL;
  assign execute_SHIFT_CTRL = _zz_execute_SHIFT_CTRL;
  assign execute_SRC_ADD_SUB = execute_SrcPlugin_addSub;
  assign execute_ALU_CTRL = _zz_execute_ALU_CTRL;
  assign execute_ALU_BITWISE_CTRL = _zz_execute_ALU_BITWISE_CTRL;
  always @(*) begin
    _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT = memory_CfuPlugin_CFU_IN_FLIGHT;
    if(memory_arbitration_isStuck) begin
      _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT = 1'b0;
    end
  end

  always @(*) begin
    _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT = execute_CfuPlugin_CFU_IN_FLIGHT;
    if(execute_arbitration_isStuck) begin
      _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT = 1'b0;
    end
  end

  assign writeBack_CfuPlugin_CFU_IN_FLIGHT = memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
  assign execute_CfuPlugin_CFU_INPUT_2_KIND = _zz_execute_CfuPlugin_CFU_INPUT_2_KIND;
  assign writeBack_HAS_SIDE_EFFECT = memory_to_writeBack_HAS_SIDE_EFFECT;
  assign memory_HAS_SIDE_EFFECT = execute_to_memory_HAS_SIDE_EFFECT;
  assign execute_LEGAL_INSTRUCTION = decode_to_execute_LEGAL_INSTRUCTION;
  always @(*) begin
    execute_CfuPlugin_CFU_ENABLE = decode_to_execute_CfuPlugin_CFU_ENABLE;
    if(when_CfuPlugin_l192) begin
      execute_CfuPlugin_CFU_ENABLE = 1'b0;
    end
  end

  always @(*) begin
    _zz_memory_to_writeBack_FPU_FORKED = memory_FPU_FORKED;
    if(memory_arbitration_isStuck) begin
      _zz_memory_to_writeBack_FPU_FORKED = 1'b0;
    end
  end

  always @(*) begin
    _zz_execute_to_memory_FPU_FORKED = execute_FPU_FORKED;
    if(execute_arbitration_isStuck) begin
      _zz_execute_to_memory_FPU_FORKED = 1'b0;
    end
  end

  always @(*) begin
    _zz_decode_to_execute_FPU_FORKED = decode_FPU_FORKED;
    if(decode_arbitration_isStuck) begin
      _zz_decode_to_execute_FPU_FORKED = 1'b0;
    end
  end

  assign writeBack_FPU_OPCODE = _zz_writeBack_FPU_OPCODE;
  assign writeBack_RS1 = memory_to_writeBack_RS1;
  assign _zz_writeBack_FpuPlugin_commit_payload_value = writeBack_MEMORY_LOAD_DATA;
  assign writeBack_FPU_COMMIT_LOAD = memory_to_writeBack_FPU_COMMIT_LOAD;
  always @(*) begin
    DBusBypass0_cond = 1'b0;
    if(writeBack_FpuPlugin_isRsp) begin
      if(writeBack_arbitration_isValid) begin
        DBusBypass0_cond = 1'b1;
      end
    end
  end

  assign writeBack_FPU_COMMIT = memory_to_writeBack_FPU_COMMIT;
  assign writeBack_FPU_RSP = memory_to_writeBack_FPU_RSP;
  assign writeBack_FPU_FORKED = memory_to_writeBack_FPU_FORKED;
  assign decode_FPU_FORMAT = _zz_decode_FPU_FORMAT;
  assign decode_FPU_ARG = _zz_decode_CfuPlugin_CFU_ENABLE[41 : 40];
  assign decode_FPU_OPCODE = _zz_decode_FPU_OPCODE;
  always @(*) begin
    decode_FPU_ENABLE = _zz_decode_FPU_ENABLE;
    if(when_FpuPlugin_l272) begin
      decode_FPU_ENABLE = 1'b0;
    end
  end

  assign execute_IS_RS1_SIGNED = decode_to_execute_IS_RS1_SIGNED;
  assign execute_IS_DIV = decode_to_execute_IS_DIV;
  assign execute_IS_RS2_SIGNED = decode_to_execute_IS_RS2_SIGNED;
  assign memory_IS_DIV = execute_to_memory_IS_DIV;
  assign writeBack_IS_MUL = memory_to_writeBack_IS_MUL;
  assign writeBack_MUL_HH = memory_to_writeBack_MUL_HH;
  assign writeBack_MUL_LOW = memory_to_writeBack_MUL_LOW;
  assign memory_MUL_HL = execute_to_memory_MUL_HL;
  assign memory_MUL_LH = execute_to_memory_MUL_LH;
  assign memory_MUL_LL = execute_to_memory_MUL_LL;
  assign execute_IS_MUL = decode_to_execute_IS_MUL;
  assign memory_BRANCH_CALC = execute_to_memory_BRANCH_CALC;
  assign memory_BRANCH_DO = execute_to_memory_BRANCH_DO;
  assign execute_PC = decode_to_execute_PC;
  assign execute_BRANCH_CTRL = _zz_execute_BRANCH_CTRL;
  assign execute_SRC_LESS = execute_SrcPlugin_less;
  assign execute_CSR_READ_OPCODE = decode_to_execute_CSR_READ_OPCODE;
  assign execute_CSR_WRITE_OPCODE = decode_to_execute_CSR_WRITE_OPCODE;
  assign execute_IS_CSR = decode_to_execute_IS_CSR;
  assign memory_ENV_CTRL = _zz_memory_ENV_CTRL;
  assign execute_ENV_CTRL = _zz_execute_ENV_CTRL;
  assign writeBack_ENV_CTRL = _zz_writeBack_ENV_CTRL;
  assign decode_RS2_USE = _zz_decode_CfuPlugin_CFU_ENABLE[18];
  assign decode_RS1_USE = _zz_decode_CfuPlugin_CFU_ENABLE[6];
  always @(*) begin
    _zz_decode_RS2 = execute_REGFILE_WRITE_DATA;
    if(when_CsrPlugin_l1731) begin
      _zz_decode_RS2 = CsrPlugin_csrMapping_readDataSignal;
    end
  end

  assign execute_REGFILE_WRITE_VALID = decode_to_execute_REGFILE_WRITE_VALID;
  assign execute_BYPASSABLE_EXECUTE_STAGE = decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  always @(*) begin
    _zz_decode_RS2_1 = memory_REGFILE_WRITE_DATA;
    if(when_MulDivIterativePlugin_l128) begin
      _zz_decode_RS2_1 = memory_MulDivIterativePlugin_div_result;
    end
    if(memory_arbitration_isValid) begin
      case(memory_SHIFT_CTRL)
        ShiftCtrlEnum_SLL_1 : begin
          _zz_decode_RS2_1 = _zz_decode_RS2_3;
        end
        ShiftCtrlEnum_SRL_1, ShiftCtrlEnum_SRA_1 : begin
          _zz_decode_RS2_1 = memory_SHIFT_RIGHT;
        end
        default : begin
        end
      endcase
    end
  end

  assign memory_REGFILE_WRITE_VALID = execute_to_memory_REGFILE_WRITE_VALID;
  assign memory_BYPASSABLE_MEMORY_STAGE = execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  assign writeBack_REGFILE_WRITE_VALID = memory_to_writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    decode_RS2 = decode_RegFilePlugin_rs2Data;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr1Match) begin
        decode_RS2 = HazardSimplePlugin_writeBackBuffer_payload_data;
      end
    end
    if(when_HazardSimplePlugin_l45) begin
      if(when_HazardSimplePlugin_l47) begin
        if(when_HazardSimplePlugin_l51) begin
          decode_RS2 = _zz_decode_RS2_2;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_1) begin
      if(memory_BYPASSABLE_MEMORY_STAGE) begin
        if(when_HazardSimplePlugin_l51_1) begin
          decode_RS2 = _zz_decode_RS2_1;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_2) begin
      if(execute_BYPASSABLE_EXECUTE_STAGE) begin
        if(when_HazardSimplePlugin_l51_2) begin
          decode_RS2 = _zz_decode_RS2;
        end
      end
    end
  end

  always @(*) begin
    decode_RS1 = decode_RegFilePlugin_rs1Data;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr0Match) begin
        decode_RS1 = HazardSimplePlugin_writeBackBuffer_payload_data;
      end
    end
    if(when_HazardSimplePlugin_l45) begin
      if(when_HazardSimplePlugin_l47) begin
        if(when_HazardSimplePlugin_l48) begin
          decode_RS1 = _zz_decode_RS2_2;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_1) begin
      if(memory_BYPASSABLE_MEMORY_STAGE) begin
        if(when_HazardSimplePlugin_l48_1) begin
          decode_RS1 = _zz_decode_RS2_1;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_2) begin
      if(execute_BYPASSABLE_EXECUTE_STAGE) begin
        if(when_HazardSimplePlugin_l48_2) begin
          decode_RS1 = _zz_decode_RS2;
        end
      end
    end
  end

  assign execute_SRC_LESS_UNSIGNED = decode_to_execute_SRC_LESS_UNSIGNED;
  assign execute_SRC2_FORCE_ZERO = decode_to_execute_SRC2_FORCE_ZERO;
  assign execute_SRC2 = decode_to_execute_SRC2;
  assign execute_SRC_USE_SUB_LESS = decode_to_execute_SRC_USE_SUB_LESS;
  assign execute_SRC1 = decode_to_execute_SRC1;
  assign _zz_decode_to_execute_PC = decode_PC;
  assign _zz_decode_to_execute_RS2 = decode_RS2;
  assign decode_SRC2_CTRL = _zz_decode_SRC2_CTRL;
  assign _zz_decode_to_execute_RS1 = decode_RS1;
  assign decode_SRC1_CTRL = _zz_decode_SRC1_CTRL;
  assign decode_SRC_USE_SUB_LESS = _zz_decode_CfuPlugin_CFU_ENABLE[4];
  assign decode_SRC_ADD_ZERO = _zz_decode_CfuPlugin_CFU_ENABLE[19];
  assign _zz_lastStageRegFileWrite_payload_address = writeBack_INSTRUCTION;
  assign _zz_lastStageRegFileWrite_valid = writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    _zz_1 = 1'b0;
    if(lastStageRegFileWrite_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign decode_INSTRUCTION_ANTICIPATED = (decode_arbitration_isStuck ? decode_INSTRUCTION : IBusCachedPlugin_decompressor_output_payload_rsp_inst);
  always @(*) begin
    decode_REGFILE_WRITE_VALID = _zz_decode_CfuPlugin_CFU_ENABLE[11];
    if(when_RegFilePlugin_l63) begin
      decode_REGFILE_WRITE_VALID = 1'b0;
    end
  end

  always @(*) begin
    decode_LEGAL_INSTRUCTION = (|{((decode_INSTRUCTION & 32'h0000005f) == 32'h00000017),{((decode_INSTRUCTION & 32'h04000073) == 32'h00000043),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION) == 32'h0000006f),{(_zz_decode_LEGAL_INSTRUCTION_1 == _zz_decode_LEGAL_INSTRUCTION_2),{_zz_decode_LEGAL_INSTRUCTION_3,{_zz_decode_LEGAL_INSTRUCTION_4,_zz_decode_LEGAL_INSTRUCTION_5}}}}}});
    if(decode_FpuPlugin_trap) begin
      decode_LEGAL_INSTRUCTION = 1'b0;
    end
  end

  always @(*) begin
    _zz_decode_RS2_2 = writeBack_REGFILE_WRITE_DATA;
    if(when_DBusCachedPlugin_l599) begin
      _zz_decode_RS2_2 = writeBack_DBusCachedPlugin_rspFormated;
    end
    if(when_MulPlugin_l147) begin
      case(switch_MulPlugin_l148)
        2'b00 : begin
          _zz_decode_RS2_2 = _zz__zz_decode_RS2_2;
        end
        default : begin
          _zz_decode_RS2_2 = _zz__zz_decode_RS2_2_1;
        end
      endcase
    end
    if(writeBack_FpuPlugin_isRsp) begin
      if(writeBack_arbitration_isValid) begin
        _zz_decode_RS2_2 = FpuPlugin_port_rsp_payload_value[31 : 0];
      end
    end
    if(writeBack_CfuPlugin_CFU_IN_FLIGHT) begin
      _zz_decode_RS2_2 = writeBack_CfuPlugin_rsp_payload_outputs_0;
    end
  end

  assign writeBack_MEMORY_WR = memory_to_writeBack_MEMORY_WR;
  assign writeBack_MEMORY_FENCE = memory_to_writeBack_MEMORY_FENCE;
  assign writeBack_MEMORY_AMO = memory_to_writeBack_MEMORY_AMO;
  assign writeBack_MEMORY_LRSC = memory_to_writeBack_MEMORY_LRSC;
  assign writeBack_MEMORY_STORE_DATA_RF = memory_to_writeBack_MEMORY_STORE_DATA_RF;
  assign writeBack_REGFILE_WRITE_DATA = memory_to_writeBack_REGFILE_WRITE_DATA;
  assign writeBack_MEMORY_ENABLE = memory_to_writeBack_MEMORY_ENABLE;
  assign memory_PC = execute_to_memory_PC;
  assign memory_MEMORY_STORE_DATA_RF = execute_to_memory_MEMORY_STORE_DATA_RF;
  assign memory_REGFILE_WRITE_DATA = execute_to_memory_REGFILE_WRITE_DATA;
  assign memory_INSTRUCTION = execute_to_memory_INSTRUCTION;
  assign memory_MEMORY_WR = execute_to_memory_MEMORY_WR;
  assign memory_MEMORY_ENABLE = execute_to_memory_MEMORY_ENABLE;
  assign execute_MEMORY_FENCE_WR = decode_to_execute_MEMORY_FENCE_WR;
  assign memory_MEMORY_VIRTUAL_ADDRESS = execute_to_memory_MEMORY_VIRTUAL_ADDRESS;
  assign execute_MEMORY_AMO = decode_to_execute_MEMORY_AMO;
  assign execute_MEMORY_LRSC = decode_to_execute_MEMORY_LRSC;
  assign execute_MEMORY_FORCE_CONSTISTENCY = decode_to_execute_MEMORY_FORCE_CONSTISTENCY;
  assign execute_RS1 = decode_to_execute_RS1;
  assign execute_MEMORY_MANAGMENT = decode_to_execute_MEMORY_MANAGMENT;
  assign execute_RS2 = decode_to_execute_RS2;
  assign execute_MEMORY_WR = decode_to_execute_MEMORY_WR;
  assign execute_SRC_ADD = execute_SrcPlugin_addSub;
  assign execute_MEMORY_ENABLE = decode_to_execute_MEMORY_ENABLE;
  assign execute_INSTRUCTION = decode_to_execute_INSTRUCTION;
  assign decode_MEMORY_AMO = _zz_decode_CfuPlugin_CFU_ENABLE[17];
  assign decode_MEMORY_LRSC = _zz_decode_CfuPlugin_CFU_ENABLE[16];
  assign decode_MEMORY_ENABLE = _zz_decode_CfuPlugin_CFU_ENABLE[5];
  assign decode_FLUSH_ALL = _zz_decode_CfuPlugin_CFU_ENABLE[0];
  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_4 = IBusCachedPlugin_rsp_issueDetected_3;
    if(when_IBusCachedPlugin_l262) begin
      IBusCachedPlugin_rsp_issueDetected_4 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_3 = IBusCachedPlugin_rsp_issueDetected_2;
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_rsp_issueDetected_3 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_2 = IBusCachedPlugin_rsp_issueDetected_1;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_issueDetected_2 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_1 = IBusCachedPlugin_rsp_issueDetected;
    if(when_IBusCachedPlugin_l245) begin
      IBusCachedPlugin_rsp_issueDetected_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_memory_to_writeBack_FORMAL_PC_NEXT = memory_FORMAL_PC_NEXT;
    if(BranchPlugin_jumpInterface_valid) begin
      _zz_memory_to_writeBack_FORMAL_PC_NEXT = BranchPlugin_jumpInterface_payload;
    end
  end

  assign decode_PC = IBusCachedPlugin_decodePc_pcReg;
  assign decode_INSTRUCTION = IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  assign decode_IS_RVC = IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  assign writeBack_PC = memory_to_writeBack_PC;
  assign writeBack_INSTRUCTION = memory_to_writeBack_INSTRUCTION;
  always @(*) begin
    decode_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l356) begin
      decode_arbitration_haltItself = 1'b1;
    end
    if(when_FpuPlugin_l273) begin
      decode_arbitration_haltItself = 1'b1;
    end
    if(FpuPlugin_port_cmd_isStall) begin
      decode_arbitration_haltItself = 1'b1;
    end
    case(IBusCachedPlugin_injector_port_state)
      3'b010 : begin
        decode_arbitration_haltItself = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    decode_arbitration_haltByOther = 1'b0;
    if(when_HazardSimplePlugin_l113) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
        if(decode_arbitration_isValid) begin
          decode_arbitration_haltByOther = 1'b1;
        end
      end
      default : begin
      end
    endcase
    if(CsrPlugin_pipelineLiberator_active) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(when_CsrPlugin_l1671) begin
      decode_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    decode_arbitration_removeIt = 1'b0;
    if(_zz_when) begin
      decode_arbitration_removeIt = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      decode_arbitration_removeIt = 1'b1;
    end
  end

  assign decode_arbitration_flushIt = 1'b0;
  always @(*) begin
    decode_arbitration_flushNext = 1'b0;
    if(_zz_when) begin
      decode_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l398) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_DBusCachedPlugin_l427) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_CsrPlugin_l1735) begin
      if(execute_CsrPlugin_blockedBySideEffects) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
    if(when_MulPlugin_l65) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_CfuPlugin_l196) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_CfuPlugin_l203) begin
      execute_arbitration_haltItself = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_haltByOther = 1'b0;
    if(when_DBusCachedPlugin_l414) begin
      execute_arbitration_haltByOther = 1'b1;
    end
    if(when_FpuPlugin_l229) begin
      execute_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_removeIt = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_removeIt = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      execute_arbitration_removeIt = 1'b1;
    end
  end

  assign execute_arbitration_flushIt = 1'b0;
  always @(*) begin
    execute_arbitration_flushNext = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    memory_arbitration_haltItself = 1'b0;
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l129) begin
        memory_arbitration_haltItself = 1'b1;
      end
    end
  end

  always @(*) begin
    memory_arbitration_haltByOther = 1'b0;
    if(when_DBusCachedPlugin_l535) begin
      memory_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    memory_arbitration_removeIt = 1'b0;
    if(DBusCachedPlugin_trigger_hitBefore) begin
      memory_arbitration_removeIt = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      memory_arbitration_removeIt = 1'b1;
    end
  end

  assign memory_arbitration_flushIt = 1'b0;
  always @(*) begin
    memory_arbitration_flushNext = 1'b0;
    if(DBusCachedPlugin_trigger_hitBefore) begin
      memory_arbitration_flushNext = 1'b1;
    end
    if(BranchPlugin_jumpInterface_valid) begin
      memory_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l572) begin
      writeBack_arbitration_haltItself = 1'b1;
    end
    if(writeBack_CfuPlugin_CFU_IN_FLIGHT) begin
      if(when_CfuPlugin_l239) begin
        writeBack_arbitration_haltItself = 1'b1;
      end
    end
  end

  always @(*) begin
    writeBack_arbitration_haltByOther = 1'b0;
    if(writeBack_FpuPlugin_isRsp) begin
      if(when_FpuPlugin_l323) begin
        writeBack_arbitration_haltByOther = 1'b1;
      end
    end
    if(when_FpuPlugin_l339) begin
      writeBack_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_removeIt = 1'b0;
    if(DBusCachedPlugin_exceptionBus_valid) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
    if(writeBack_arbitration_isFlushed) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_flushIt = 1'b0;
    if(DBusCachedPlugin_redoBranch_valid) begin
      writeBack_arbitration_flushIt = 1'b1;
    end
    if(CsrPlugin_doResume) begin
      writeBack_arbitration_flushIt = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_flushNext = 1'b0;
    if(DBusCachedPlugin_redoBranch_valid) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(DBusCachedPlugin_exceptionBus_valid) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1534) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1600) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
  end

  assign lastStageInstruction = writeBack_INSTRUCTION;
  assign lastStagePc = writeBack_PC;
  assign lastStageIsValid = writeBack_arbitration_isValid;
  assign lastStageIsFiring = writeBack_arbitration_isFiring;
  always @(*) begin
    IBusCachedPlugin_fetcherHalt = 1'b0;
    if(when_CsrPlugin_l729) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1416) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1534) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1600) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
  end

  assign IBusCachedPlugin_forceNoDecodeCond = 1'b0;
  always @(*) begin
    IBusCachedPlugin_incomingInstruction = 1'b0;
    if(when_Fetcher_l242) begin
      IBusCachedPlugin_incomingInstruction = 1'b1;
    end
    if(IBusCachedPlugin_injector_decodeInput_valid) begin
      IBusCachedPlugin_incomingInstruction = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_csrMapping_allowCsrSignal = 1'b0;
    if(when_CsrPlugin_l1846) begin
      CsrPlugin_csrMapping_allowCsrSignal = 1'b1;
    end
    if(when_CsrPlugin_l1853) begin
      CsrPlugin_csrMapping_allowCsrSignal = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_csrMapping_doForceFailCsr = 1'b0;
    if(when_FpuPlugin_l253) begin
      CsrPlugin_csrMapping_doForceFailCsr = 1'b1;
    end
  end

  assign CsrPlugin_csrMapping_readDataSignal = CsrPlugin_csrMapping_readDataInit;
  assign CsrPlugin_inWfi = 1'b0;
  always @(*) begin
    CsrPlugin_thirdPartyWake = 1'b0;
    if(when_CsrPlugin_l880) begin
      CsrPlugin_thirdPartyWake = 1'b1;
    end
    if(decode_FpuPlugin_forked) begin
      CsrPlugin_thirdPartyWake = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_valid = 1'b0;
    if(when_CsrPlugin_l1534) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
    if(when_CsrPlugin_l1600) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
    if(CsrPlugin_doResume) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CsrPlugin_l1534) begin
      CsrPlugin_jumpInterface_payload = {CsrPlugin_xtvec_base,2'b00};
    end
    if(when_CsrPlugin_l1600) begin
      case(switch_CsrPlugin_l1604)
        2'b11 : begin
          CsrPlugin_jumpInterface_payload = CsrPlugin_mepc;
        end
        default : begin
        end
      endcase
    end
    if(CsrPlugin_doResume) begin
      CsrPlugin_jumpInterface_payload = CsrPlugin_dpc;
    end
  end

  assign CsrPlugin_forceMachineWire = 1'b0;
  always @(*) begin
    CsrPlugin_allowInterrupts = 1'b1;
    if(debugMode) begin
      CsrPlugin_allowInterrupts = 1'b0;
    end
  end

  assign CsrPlugin_allowException = 1'b1;
  assign CsrPlugin_allowEbreakException = 1'b1;
  always @(*) begin
    CsrPlugin_xretAwayFromMachine = 1'b0;
    if(when_CsrPlugin_l1600) begin
      case(switch_CsrPlugin_l1604)
        2'b11 : begin
          if(when_CsrPlugin_l1612) begin
            CsrPlugin_xretAwayFromMachine = 1'b1;
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    BranchPlugin_inDebugNoFetchFlag = 1'b0;
    if(debugMode) begin
      BranchPlugin_inDebugNoFetchFlag = 1'b1;
    end
  end

  assign IBusCachedPlugin_mmuBus_rsp_physicalAddress = IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign IBusCachedPlugin_mmuBus_rsp_allowRead = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowWrite = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_allowExecute = 1'b1;
  assign IBusCachedPlugin_mmuBus_rsp_isIoAccess = (((IBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'hf8000000) || ((IBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'he1000000));
  assign IBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign IBusCachedPlugin_mmuBus_busy = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_physicalAddress = DBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign DBusCachedPlugin_mmuBus_rsp_allowRead = 1'b1;
  assign DBusCachedPlugin_mmuBus_rsp_allowWrite = 1'b1;
  assign DBusCachedPlugin_mmuBus_rsp_allowExecute = 1'b1;
  assign DBusCachedPlugin_mmuBus_rsp_isIoAccess = (((DBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'hf8000000) || ((DBusCachedPlugin_mmuBus_rsp_physicalAddress & (~ 32'h00ffffff)) == 32'he1000000));
  assign DBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign DBusCachedPlugin_mmuBus_busy = 1'b0;
  assign IBusCachedPlugin_externalFlush = (|{writeBack_arbitration_flushNext,{memory_arbitration_flushNext,{execute_arbitration_flushNext,decode_arbitration_flushNext}}});
  assign IBusCachedPlugin_jump_pcLoad_valid = (|{BranchPlugin_jumpInterface_valid,{CsrPlugin_jumpInterface_valid,DBusCachedPlugin_redoBranch_valid}});
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload = {BranchPlugin_jumpInterface_valid,{CsrPlugin_jumpInterface_valid,DBusCachedPlugin_redoBranch_valid}};
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload & (~ _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1));
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_2 = _zz_IBusCachedPlugin_jump_pcLoad_payload_1[1];
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_3 = _zz_IBusCachedPlugin_jump_pcLoad_payload_1[2];
  assign IBusCachedPlugin_jump_pcLoad_payload = _zz_IBusCachedPlugin_jump_pcLoad_payload_4;
  always @(*) begin
    IBusCachedPlugin_fetchPc_correction = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
  end

  assign IBusCachedPlugin_fetchPc_output_fire = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign IBusCachedPlugin_fetchPc_corrected = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_correctionReg);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b0;
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b1;
    end
  end

  assign when_Fetcher_l133 = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_pcRegPropagate);
  assign when_Fetcher_l133_1 = ((! IBusCachedPlugin_fetchPc_output_valid) && IBusCachedPlugin_fetchPc_output_ready);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pc = (IBusCachedPlugin_fetchPc_pcReg + _zz_IBusCachedPlugin_fetchPc_pc);
    if(IBusCachedPlugin_fetchPc_inc) begin
      IBusCachedPlugin_fetchPc_pc[1] = 1'b0;
    end
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_fetchPc_redo_payload;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_jump_pcLoad_payload;
    end
    IBusCachedPlugin_fetchPc_pc[0] = 1'b0;
  end

  always @(*) begin
    IBusCachedPlugin_fetchPc_flushed = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
  end

  assign when_Fetcher_l160 = (IBusCachedPlugin_fetchPc_booted && ((IBusCachedPlugin_fetchPc_output_ready || IBusCachedPlugin_fetchPc_correction) || IBusCachedPlugin_fetchPc_pcRegPropagate));
  assign IBusCachedPlugin_fetchPc_output_valid = ((! IBusCachedPlugin_fetcherHalt) && IBusCachedPlugin_fetchPc_booted);
  assign IBusCachedPlugin_fetchPc_output_payload = IBusCachedPlugin_fetchPc_pc;
  always @(*) begin
    IBusCachedPlugin_decodePc_flushed = 1'b0;
    if(when_Fetcher_l194) begin
      IBusCachedPlugin_decodePc_flushed = 1'b1;
    end
  end

  assign IBusCachedPlugin_decodePc_pcPlus = (IBusCachedPlugin_decodePc_pcReg + _zz_IBusCachedPlugin_decodePc_pcPlus);
  always @(*) begin
    IBusCachedPlugin_decodePc_injectedDecode = 1'b0;
    if(when_Fetcher_l373) begin
      IBusCachedPlugin_decodePc_injectedDecode = 1'b1;
    end
  end

  assign when_Fetcher_l182 = (decode_arbitration_isFiring && (! IBusCachedPlugin_decodePc_injectedDecode));
  assign when_Fetcher_l194 = (IBusCachedPlugin_jump_pcLoad_valid && ((! decode_arbitration_isStuck) || decode_arbitration_removeIt));
  always @(*) begin
    IBusCachedPlugin_iBusRsp_redoFetch = 1'b0;
    if(IBusCachedPlugin_rsp_redoFetch) begin
      IBusCachedPlugin_iBusRsp_redoFetch = 1'b1;
    end
  end

  assign IBusCachedPlugin_iBusRsp_stages_0_input_valid = IBusCachedPlugin_fetchPc_output_valid;
  assign IBusCachedPlugin_fetchPc_output_ready = IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_0_input_payload = IBusCachedPlugin_fetchPc_output_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b0;
    if(IBusCachedPlugin_cache_io_cpu_prefetch_haltIt) begin
      IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready = (! IBusCachedPlugin_iBusRsp_stages_0_halt);
  assign IBusCachedPlugin_iBusRsp_stages_0_input_ready = (IBusCachedPlugin_iBusRsp_stages_0_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_valid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_payload = IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b0;
    if(IBusCachedPlugin_mmuBus_busy) begin
      IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready = (! IBusCachedPlugin_iBusRsp_stages_1_halt);
  assign IBusCachedPlugin_iBusRsp_stages_1_input_ready = (IBusCachedPlugin_iBusRsp_stages_1_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_valid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_payload = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b0;
    if(when_IBusCachedPlugin_l273) begin
      IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready = (! IBusCachedPlugin_iBusRsp_stages_2_halt);
  assign IBusCachedPlugin_iBusRsp_stages_2_input_ready = (IBusCachedPlugin_iBusRsp_stages_2_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_valid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_fetchPc_redo_valid = IBusCachedPlugin_iBusRsp_redoFetch;
  always @(*) begin
    IBusCachedPlugin_fetchPc_redo_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
    if(IBusCachedPlugin_decompressor_throw2BytesReg) begin
      IBusCachedPlugin_fetchPc_redo_payload[1] = 1'b1;
    end
  end

  assign IBusCachedPlugin_iBusRsp_flush = (IBusCachedPlugin_externalFlush || IBusCachedPlugin_iBusRsp_redoFetch);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_ready = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready = ((1'b0 && (! _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid)) || IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_payload = IBusCachedPlugin_fetchPc_pcReg;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_ready = ((1'b0 && (! IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid)) || IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_valid = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready = IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_payload = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_readyForError = 1'b1;
    if(IBusCachedPlugin_injector_decodeInput_valid) begin
      IBusCachedPlugin_iBusRsp_readyForError = 1'b0;
    end
  end

  assign when_Fetcher_l242 = (IBusCachedPlugin_iBusRsp_stages_1_input_valid || IBusCachedPlugin_iBusRsp_stages_2_input_valid);
  assign IBusCachedPlugin_decompressor_input_valid = (IBusCachedPlugin_iBusRsp_output_valid && (! IBusCachedPlugin_iBusRsp_redoFetch));
  assign IBusCachedPlugin_decompressor_input_payload_pc = IBusCachedPlugin_iBusRsp_output_payload_pc;
  assign IBusCachedPlugin_decompressor_input_payload_rsp_error = IBusCachedPlugin_iBusRsp_output_payload_rsp_error;
  assign IBusCachedPlugin_decompressor_input_payload_rsp_inst = IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  assign IBusCachedPlugin_decompressor_input_payload_isRvc = IBusCachedPlugin_iBusRsp_output_payload_isRvc;
  assign IBusCachedPlugin_iBusRsp_output_ready = IBusCachedPlugin_decompressor_input_ready;
  assign IBusCachedPlugin_decompressor_flushNext = 1'b0;
  assign IBusCachedPlugin_decompressor_consumeCurrent = 1'b0;
  assign IBusCachedPlugin_decompressor_isInputLowRvc = (IBusCachedPlugin_decompressor_input_payload_rsp_inst[1 : 0] != 2'b11);
  assign IBusCachedPlugin_decompressor_isInputHighRvc = (IBusCachedPlugin_decompressor_input_payload_rsp_inst[17 : 16] != 2'b11);
  assign IBusCachedPlugin_decompressor_throw2Bytes = (IBusCachedPlugin_decompressor_throw2BytesReg || IBusCachedPlugin_decompressor_input_payload_pc[1]);
  assign IBusCachedPlugin_decompressor_unaligned = (IBusCachedPlugin_decompressor_throw2Bytes || IBusCachedPlugin_decompressor_bufferValid);
  assign IBusCachedPlugin_decompressor_bufferValidPatched = (IBusCachedPlugin_decompressor_input_valid ? IBusCachedPlugin_decompressor_bufferValid : IBusCachedPlugin_decompressor_bufferValidLatch);
  assign IBusCachedPlugin_decompressor_throw2BytesPatched = (IBusCachedPlugin_decompressor_input_valid ? IBusCachedPlugin_decompressor_throw2Bytes : IBusCachedPlugin_decompressor_throw2BytesLatch);
  assign IBusCachedPlugin_decompressor_raw = (IBusCachedPlugin_decompressor_bufferValidPatched ? {IBusCachedPlugin_decompressor_input_payload_rsp_inst[15 : 0],IBusCachedPlugin_decompressor_bufferData} : {IBusCachedPlugin_decompressor_input_payload_rsp_inst[31 : 16],(IBusCachedPlugin_decompressor_throw2BytesPatched ? IBusCachedPlugin_decompressor_input_payload_rsp_inst[31 : 16] : IBusCachedPlugin_decompressor_input_payload_rsp_inst[15 : 0])});
  assign IBusCachedPlugin_decompressor_isRvc = (IBusCachedPlugin_decompressor_raw[1 : 0] != 2'b11);
  assign _zz_IBusCachedPlugin_decompressor_decompressed = IBusCachedPlugin_decompressor_raw[15 : 0];
  always @(*) begin
    IBusCachedPlugin_decompressor_decompressed = 32'h0;
    case(switch_Misc_l44)
      5'h0 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{{2'b00,_zz_IBusCachedPlugin_decompressor_decompressed[10 : 7]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 11]},_zz_IBusCachedPlugin_decompressor_decompressed[5]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},2'b00},5'h02},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h13};
        if(when_Misc_l47) begin
          IBusCachedPlugin_decompressor_decompressed = 32'h0;
        end
      end
      5'h01 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_4,_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h07};
      end
      5'h02 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_3,_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h03};
      end
      5'h03 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_3,_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_2},7'h07};
      end
      5'h05 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_4[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed_2},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed_4[4 : 0]},7'h27};
      end
      5'h06 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_3[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed_2},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_3[4 : 0]},7'h23};
      end
      5'h07 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_3[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed_2},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_3[4 : 0]},7'h27};
      end
      5'h08 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_6,_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13};
      end
      5'h09 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_9[20],_zz_IBusCachedPlugin_decompressor_decompressed_9[10 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_9[11]},_zz_IBusCachedPlugin_decompressor_decompressed_9[19 : 12]},_zz_IBusCachedPlugin_decompressor_decompressed_21},7'h6f};
      end
      5'h0a : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{_zz_IBusCachedPlugin_decompressor_decompressed_6,5'h0},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13};
      end
      5'h0b : begin
        IBusCachedPlugin_decompressor_decompressed = ((_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7] == 5'h02) ? {{{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_28,_zz_IBusCachedPlugin_decompressor_decompressed_29},_zz_IBusCachedPlugin_decompressor_decompressed_30},_zz_IBusCachedPlugin_decompressor_decompressed[6]},4'b0000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13} : {{_zz_IBusCachedPlugin_decompressor_decompressed_31[31 : 12],_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h37});
      end
      5'h0c : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{((_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] == 2'b10) ? _zz_IBusCachedPlugin_decompressor_decompressed_27 : {{1'b0,(_zz_IBusCachedPlugin_decompressor_decompressed_32 || _zz_IBusCachedPlugin_decompressor_decompressed_33)},5'h0}),(((! _zz_IBusCachedPlugin_decompressor_decompressed[11]) || _zz_IBusCachedPlugin_decompressor_decompressed_23) ? _zz_IBusCachedPlugin_decompressor_decompressed[6 : 2] : _zz_IBusCachedPlugin_decompressor_decompressed_2)},_zz_IBusCachedPlugin_decompressor_decompressed_1},_zz_IBusCachedPlugin_decompressor_decompressed_25},_zz_IBusCachedPlugin_decompressor_decompressed_1},(_zz_IBusCachedPlugin_decompressor_decompressed_23 ? 7'h13 : 7'h33)};
      end
      5'h0d : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_16[20],_zz_IBusCachedPlugin_decompressor_decompressed_16[10 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_16[11]},_zz_IBusCachedPlugin_decompressor_decompressed_16[19 : 12]},_zz_IBusCachedPlugin_decompressor_decompressed_20},7'h6f};
      end
      5'h0e : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_19[12],_zz_IBusCachedPlugin_decompressor_decompressed_19[10 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed_20},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed_19[4 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_19[11]},7'h63};
      end
      5'h0f : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_19[12],_zz_IBusCachedPlugin_decompressor_decompressed_19[10 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed_20},_zz_IBusCachedPlugin_decompressor_decompressed_1},3'b001},_zz_IBusCachedPlugin_decompressor_decompressed_19[4 : 1]},_zz_IBusCachedPlugin_decompressor_decompressed_19[11]},7'h63};
      end
      5'h10 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{7'h0,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b001},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h13};
      end
      5'h11 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{3'b000,_zz_IBusCachedPlugin_decompressor_decompressed[4 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[12]},_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5]},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h07};
      end
      5'h12 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[3 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[12]},_zz_IBusCachedPlugin_decompressor_decompressed[6 : 4]},2'b00},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h03};
      end
      5'h13 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{{{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[3 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed[12]},_zz_IBusCachedPlugin_decompressor_decompressed[6 : 4]},2'b00},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h07};
      end
      5'h14 : begin
        IBusCachedPlugin_decompressor_decompressed = ((_zz_IBusCachedPlugin_decompressor_decompressed[12 : 2] == 11'h400) ? 32'h00100073 : ((_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2] == 5'h0) ? {{{{12'h0,_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},3'b000},(_zz_IBusCachedPlugin_decompressor_decompressed[12] ? _zz_IBusCachedPlugin_decompressor_decompressed_21 : _zz_IBusCachedPlugin_decompressor_decompressed_20)},7'h67} : {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_34,_zz_IBusCachedPlugin_decompressor_decompressed_35},(_zz_IBusCachedPlugin_decompressor_decompressed_36 ? _zz_IBusCachedPlugin_decompressor_decompressed_37 : _zz_IBusCachedPlugin_decompressor_decompressed_20)},3'b000},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 7]},7'h33}));
      end
      5'h15 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_38[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b011},_zz_IBusCachedPlugin_decompressor_decompressed_39[4 : 0]},7'h27};
      end
      5'h16 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_40[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_41[4 : 0]},7'h23};
      end
      5'h17 : begin
        IBusCachedPlugin_decompressor_decompressed = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_42[11 : 5],_zz_IBusCachedPlugin_decompressor_decompressed[6 : 2]},_zz_IBusCachedPlugin_decompressor_decompressed_22},3'b010},_zz_IBusCachedPlugin_decompressor_decompressed_43[4 : 0]},7'h27};
      end
      default : begin
      end
    endcase
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_1 = {2'b01,_zz_IBusCachedPlugin_decompressor_decompressed[9 : 7]};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_2 = {2'b01,_zz_IBusCachedPlugin_decompressor_decompressed[4 : 2]};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_3 = {{{{5'h0,_zz_IBusCachedPlugin_decompressor_decompressed[5]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},2'b00};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_4 = {{{4'b0000,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed[12 : 10]},3'b000};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_5 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_6[11] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[10] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[9] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[8] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[7] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[6] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[5] = _zz_IBusCachedPlugin_decompressor_decompressed_5;
    _zz_IBusCachedPlugin_decompressor_decompressed_6[4 : 0] = _zz_IBusCachedPlugin_decompressor_decompressed[6 : 2];
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_7 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_8[9] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[8] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[7] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[6] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[5] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[4] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[3] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[2] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[1] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
    _zz_IBusCachedPlugin_decompressor_decompressed_8[0] = _zz_IBusCachedPlugin_decompressor_decompressed_7;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_9 = {{{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_8,_zz_IBusCachedPlugin_decompressor_decompressed[8]},_zz_IBusCachedPlugin_decompressor_decompressed[10 : 9]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},_zz_IBusCachedPlugin_decompressor_decompressed[7]},_zz_IBusCachedPlugin_decompressor_decompressed[2]},_zz_IBusCachedPlugin_decompressor_decompressed[11]},_zz_IBusCachedPlugin_decompressor_decompressed[5 : 3]},1'b0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_10 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_11[14] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[13] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[12] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[11] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[10] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[9] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[8] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[7] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[6] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[5] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[4] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[3] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[2] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[1] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
    _zz_IBusCachedPlugin_decompressor_decompressed_11[0] = _zz_IBusCachedPlugin_decompressor_decompressed_10;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_12 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_13[2] = _zz_IBusCachedPlugin_decompressor_decompressed_12;
    _zz_IBusCachedPlugin_decompressor_decompressed_13[1] = _zz_IBusCachedPlugin_decompressor_decompressed_12;
    _zz_IBusCachedPlugin_decompressor_decompressed_13[0] = _zz_IBusCachedPlugin_decompressor_decompressed_12;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_14 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_15[9] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[8] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[7] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[6] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[5] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[4] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[3] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[2] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[1] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
    _zz_IBusCachedPlugin_decompressor_decompressed_15[0] = _zz_IBusCachedPlugin_decompressor_decompressed_14;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_16 = {{{{{{{{_zz_IBusCachedPlugin_decompressor_decompressed_15,_zz_IBusCachedPlugin_decompressor_decompressed[8]},_zz_IBusCachedPlugin_decompressor_decompressed[10 : 9]},_zz_IBusCachedPlugin_decompressor_decompressed[6]},_zz_IBusCachedPlugin_decompressor_decompressed[7]},_zz_IBusCachedPlugin_decompressor_decompressed[2]},_zz_IBusCachedPlugin_decompressor_decompressed[11]},_zz_IBusCachedPlugin_decompressor_decompressed[5 : 3]},1'b0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_17 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_18[4] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[3] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[2] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[1] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
    _zz_IBusCachedPlugin_decompressor_decompressed_18[0] = _zz_IBusCachedPlugin_decompressor_decompressed_17;
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_19 = {{{{{_zz_IBusCachedPlugin_decompressor_decompressed_18,_zz_IBusCachedPlugin_decompressor_decompressed[6 : 5]},_zz_IBusCachedPlugin_decompressor_decompressed[2]},_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10]},_zz_IBusCachedPlugin_decompressor_decompressed[4 : 3]},1'b0};
  assign _zz_IBusCachedPlugin_decompressor_decompressed_20 = 5'h0;
  assign _zz_IBusCachedPlugin_decompressor_decompressed_21 = 5'h01;
  assign _zz_IBusCachedPlugin_decompressor_decompressed_22 = 5'h02;
  assign switch_Misc_l44 = {_zz_IBusCachedPlugin_decompressor_decompressed[1 : 0],_zz_IBusCachedPlugin_decompressor_decompressed[15 : 13]};
  assign when_Misc_l47 = (_zz_IBusCachedPlugin_decompressor_decompressed[12 : 2] == 11'h0);
  assign _zz_IBusCachedPlugin_decompressor_decompressed_23 = (_zz_IBusCachedPlugin_decompressor_decompressed[11 : 10] != 2'b11);
  assign switch_Misc_l241 = _zz_IBusCachedPlugin_decompressor_decompressed[11 : 10];
  assign switch_Misc_l241_1 = _zz_IBusCachedPlugin_decompressor_decompressed[6 : 5];
  always @(*) begin
    case(switch_Misc_l241_1)
      2'b00 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b000;
      end
      2'b01 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b100;
      end
      2'b10 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b110;
      end
      default : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_24 = 3'b111;
      end
    endcase
  end

  always @(*) begin
    case(switch_Misc_l241)
      2'b00 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = 3'b101;
      end
      2'b01 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = 3'b101;
      end
      2'b10 : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = 3'b111;
      end
      default : begin
        _zz_IBusCachedPlugin_decompressor_decompressed_25 = _zz_IBusCachedPlugin_decompressor_decompressed_24;
      end
    endcase
  end

  assign _zz_IBusCachedPlugin_decompressor_decompressed_26 = _zz_IBusCachedPlugin_decompressor_decompressed[12];
  always @(*) begin
    _zz_IBusCachedPlugin_decompressor_decompressed_27[6] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[5] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[4] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[3] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[2] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[1] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
    _zz_IBusCachedPlugin_decompressor_decompressed_27[0] = _zz_IBusCachedPlugin_decompressor_decompressed_26;
  end

  assign IBusCachedPlugin_decompressor_output_valid = (IBusCachedPlugin_decompressor_input_valid && (! ((IBusCachedPlugin_decompressor_throw2Bytes && (! IBusCachedPlugin_decompressor_bufferValid)) && (! IBusCachedPlugin_decompressor_isInputHighRvc))));
  assign IBusCachedPlugin_decompressor_output_payload_pc = IBusCachedPlugin_decompressor_input_payload_pc;
  assign IBusCachedPlugin_decompressor_output_payload_isRvc = IBusCachedPlugin_decompressor_isRvc;
  assign IBusCachedPlugin_decompressor_output_payload_rsp_inst = (IBusCachedPlugin_decompressor_isRvc ? IBusCachedPlugin_decompressor_decompressed : IBusCachedPlugin_decompressor_raw);
  assign IBusCachedPlugin_decompressor_input_ready = (IBusCachedPlugin_decompressor_output_ready && (((! IBusCachedPlugin_iBusRsp_stages_2_input_valid) || IBusCachedPlugin_decompressor_flushNext) || ((! (IBusCachedPlugin_decompressor_bufferValid && IBusCachedPlugin_decompressor_isInputHighRvc)) && (! (((! IBusCachedPlugin_decompressor_unaligned) && IBusCachedPlugin_decompressor_isInputLowRvc) && IBusCachedPlugin_decompressor_isInputHighRvc)))));
  assign IBusCachedPlugin_decompressor_output_fire = (IBusCachedPlugin_decompressor_output_valid && IBusCachedPlugin_decompressor_output_ready);
  assign IBusCachedPlugin_decompressor_bufferFill = (((((! IBusCachedPlugin_decompressor_unaligned) && IBusCachedPlugin_decompressor_isInputLowRvc) && (! IBusCachedPlugin_decompressor_isInputHighRvc)) || (IBusCachedPlugin_decompressor_bufferValid && (! IBusCachedPlugin_decompressor_isInputHighRvc))) || ((IBusCachedPlugin_decompressor_throw2Bytes && (! IBusCachedPlugin_decompressor_isRvc)) && (! IBusCachedPlugin_decompressor_isInputHighRvc)));
  assign when_Fetcher_l285 = (IBusCachedPlugin_decompressor_output_ready && IBusCachedPlugin_decompressor_input_valid);
  assign when_Fetcher_l288 = (IBusCachedPlugin_decompressor_output_ready && IBusCachedPlugin_decompressor_input_valid);
  assign when_Fetcher_l293 = (IBusCachedPlugin_externalFlush || IBusCachedPlugin_decompressor_consumeCurrent);
  assign IBusCachedPlugin_decompressor_output_ready = ((1'b0 && (! IBusCachedPlugin_injector_decodeInput_valid)) || IBusCachedPlugin_injector_decodeInput_ready);
  assign IBusCachedPlugin_injector_decodeInput_valid = _zz_IBusCachedPlugin_injector_decodeInput_valid;
  assign IBusCachedPlugin_injector_decodeInput_payload_pc = _zz_IBusCachedPlugin_injector_decodeInput_payload_pc;
  assign IBusCachedPlugin_injector_decodeInput_payload_rsp_error = _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_error;
  assign IBusCachedPlugin_injector_decodeInput_payload_rsp_inst = _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst;
  assign IBusCachedPlugin_injector_decodeInput_payload_isRvc = _zz_IBusCachedPlugin_injector_decodeInput_payload_isRvc;
  assign when_Fetcher_l331 = (! 1'b0);
  assign when_Fetcher_l331_1 = (! execute_arbitration_isStuck);
  assign when_Fetcher_l331_2 = (! memory_arbitration_isStuck);
  assign when_Fetcher_l331_3 = (! writeBack_arbitration_isStuck);
  assign IBusCachedPlugin_pcValids_0 = IBusCachedPlugin_injector_nextPcCalc_valids_0;
  assign IBusCachedPlugin_pcValids_1 = IBusCachedPlugin_injector_nextPcCalc_valids_1;
  assign IBusCachedPlugin_pcValids_2 = IBusCachedPlugin_injector_nextPcCalc_valids_2;
  assign IBusCachedPlugin_pcValids_3 = IBusCachedPlugin_injector_nextPcCalc_valids_3;
  assign IBusCachedPlugin_injector_decodeInput_ready = (! decode_arbitration_isStuck);
  always @(*) begin
    decode_arbitration_isValid = IBusCachedPlugin_injector_decodeInput_valid;
    case(IBusCachedPlugin_injector_port_state)
      3'b010 : begin
        decode_arbitration_isValid = 1'b1;
      end
      3'b011 : begin
        decode_arbitration_isValid = 1'b1;
      end
      default : begin
      end
    endcase
    if(IBusCachedPlugin_forceNoDecodeCond) begin
      decode_arbitration_isValid = 1'b0;
    end
  end

  assign iBus_cmd_valid = IBusCachedPlugin_cache_io_mem_cmd_valid;
  always @(*) begin
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  end

  assign iBus_cmd_payload_size = IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  assign IBusCachedPlugin_s0_tightlyCoupledHit = 1'b0;
  assign IBusCachedPlugin_cache_io_cpu_prefetch_isValid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && (! IBusCachedPlugin_s0_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isValid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && (! IBusCachedPlugin_s1_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_isValid = IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  assign IBusCachedPlugin_mmuBus_cmd_0_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_virtualAddress = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  assign IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign IBusCachedPlugin_mmuBus_end = (IBusCachedPlugin_iBusRsp_stages_1_input_ready || IBusCachedPlugin_externalFlush);
  assign IBusCachedPlugin_cache_io_cpu_decode_isValid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && (! IBusCachedPlugin_s2_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_decode_isStuck = (! IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_cache_io_cpu_decode_isUser = (CsrPlugin_privilege == 2'b00);
  assign IBusCachedPlugin_rsp_iBusRspOutputHalt = 1'b0;
  assign IBusCachedPlugin_rsp_issueDetected = 1'b0;
  always @(*) begin
    IBusCachedPlugin_rsp_redoFetch = 1'b0;
    if(when_IBusCachedPlugin_l245) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_cache_io_cpu_fill_valid = (IBusCachedPlugin_rsp_redoFetch && (! IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling));
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_cache_io_cpu_fill_valid = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_valid = 1'b0;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
    if(when_IBusCachedPlugin_l262) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_payload_code = 4'bxxxx;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b1100;
    end
    if(when_IBusCachedPlugin_l262) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b0001;
    end
  end

  assign IBusCachedPlugin_decodeExceptionPort_payload_badAddr = {IBusCachedPlugin_iBusRsp_stages_2_input_payload[31 : 2],2'b00};
  assign when_IBusCachedPlugin_l245 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling) && (! IBusCachedPlugin_rsp_issueDetected));
  assign when_IBusCachedPlugin_l250 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuException) && (! IBusCachedPlugin_rsp_issueDetected_1));
  assign when_IBusCachedPlugin_l256 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_cacheMiss) && (! IBusCachedPlugin_rsp_issueDetected_2));
  assign when_IBusCachedPlugin_l262 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_error) && (! IBusCachedPlugin_rsp_issueDetected_3));
  assign when_IBusCachedPlugin_l273 = (IBusCachedPlugin_rsp_issueDetected_4 || IBusCachedPlugin_rsp_iBusRspOutputHalt);
  assign IBusCachedPlugin_iBusRsp_output_valid = IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  assign IBusCachedPlugin_iBusRsp_stages_2_output_ready = IBusCachedPlugin_iBusRsp_output_ready;
  assign IBusCachedPlugin_iBusRsp_output_payload_rsp_inst = IBusCachedPlugin_cache_io_cpu_decode_data;
  assign IBusCachedPlugin_iBusRsp_output_payload_pc = IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  assign IBusCachedPlugin_cache_io_flush = (decode_arbitration_isValid && decode_FLUSH_ALL);
  assign dataCache_2_io_mem_cmd_s2mPipe_valid = (dataCache_2_io_mem_cmd_valid || (! dataCache_2_io_mem_cmd_rValidN));
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_wr = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_wr : dataCache_2_io_mem_cmd_rData_wr);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_uncached = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_uncached : dataCache_2_io_mem_cmd_rData_uncached);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_address = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_address : dataCache_2_io_mem_cmd_rData_address);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_data = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_data : dataCache_2_io_mem_cmd_rData_data);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_mask = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_mask : dataCache_2_io_mem_cmd_rData_mask);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_size = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_size : dataCache_2_io_mem_cmd_rData_size);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_exclusive = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_exclusive : dataCache_2_io_mem_cmd_rData_exclusive);
  assign dataCache_2_io_mem_cmd_s2mPipe_payload_last = (dataCache_2_io_mem_cmd_rValidN ? dataCache_2_io_mem_cmd_payload_last : dataCache_2_io_mem_cmd_rData_last);
  always @(*) begin
    dataCache_2_io_mem_cmd_s2mPipe_ready = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l375) begin
      dataCache_2_io_mem_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid);
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid = dataCache_2_io_mem_cmd_s2mPipe_rValid;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_wr = dataCache_2_io_mem_cmd_s2mPipe_rData_wr;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached = dataCache_2_io_mem_cmd_s2mPipe_rData_uncached;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_address = dataCache_2_io_mem_cmd_s2mPipe_rData_address;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_data = dataCache_2_io_mem_cmd_s2mPipe_rData_data;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_mask = dataCache_2_io_mem_cmd_s2mPipe_rData_mask;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_size = dataCache_2_io_mem_cmd_s2mPipe_rData_size;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_exclusive = dataCache_2_io_mem_cmd_s2mPipe_rData_exclusive;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_last = dataCache_2_io_mem_cmd_s2mPipe_rData_last;
  assign dBus_cmd_valid = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_valid;
  assign dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_ready = dBus_cmd_ready;
  assign dBus_cmd_payload_wr = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_wr;
  assign dBus_cmd_payload_uncached = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached;
  assign dBus_cmd_payload_address = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_address;
  assign dBus_cmd_payload_data = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_data;
  assign dBus_cmd_payload_mask = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_mask;
  assign dBus_cmd_payload_size = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_size;
  assign dBus_cmd_payload_exclusive = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_exclusive;
  assign dBus_cmd_payload_last = dataCache_2_io_mem_cmd_s2mPipe_m2sPipe_payload_last;
  assign when_DBusCachedPlugin_l334 = (dBus_rsp_valid && (! dataCache_2_io_cpu_writeBack_keepMemRspData));
  assign dBus_inv_ready = dataCache_2_io_mem_inv_ready;
  assign dBus_ack_valid = dataCache_2_io_mem_ack_valid;
  assign dBus_ack_payload_last = dataCache_2_io_mem_ack_payload_last;
  assign dBus_ack_payload_fragment_hit = dataCache_2_io_mem_ack_payload_fragment_hit;
  assign dBus_sync_ready = dataCache_2_io_mem_sync_ready;
  assign when_DBusCachedPlugin_l356 = ((DBusCachedPlugin_mmuBus_busy && decode_arbitration_isValid) && decode_MEMORY_ENABLE);
  always @(*) begin
    _zz_decode_MEMORY_FORCE_CONSTISTENCY = 1'b0;
    if(when_DBusCachedPlugin_l364) begin
      if(decode_MEMORY_LRSC) begin
        _zz_decode_MEMORY_FORCE_CONSTISTENCY = 1'b1;
      end
      if(decode_MEMORY_AMO) begin
        _zz_decode_MEMORY_FORCE_CONSTISTENCY = 1'b1;
      end
    end
  end

  assign when_DBusCachedPlugin_l364 = decode_INSTRUCTION[25];
  assign execute_DBusCachedPlugin_size = execute_INSTRUCTION[13 : 12];
  assign dataCache_2_io_cpu_execute_isValid = (execute_arbitration_isValid && execute_MEMORY_ENABLE);
  assign dataCache_2_io_cpu_execute_address = execute_SRC_ADD;
  always @(*) begin
    case(execute_DBusCachedPlugin_size)
      2'b00 : begin
        _zz_execute_MEMORY_STORE_DATA_RF = {{{execute_RS2[7 : 0],execute_RS2[7 : 0]},execute_RS2[7 : 0]},execute_RS2[7 : 0]};
      end
      2'b01 : begin
        _zz_execute_MEMORY_STORE_DATA_RF = {execute_RS2[15 : 0],execute_RS2[15 : 0]};
      end
      default : begin
        _zz_execute_MEMORY_STORE_DATA_RF = execute_RS2[31 : 0];
      end
    endcase
  end

  assign dataCache_2_io_cpu_flush_valid = (execute_arbitration_isValid && execute_MEMORY_MANAGMENT);
  assign dataCache_2_io_cpu_flush_payload_singleLine = (execute_INSTRUCTION[19 : 15] != 5'h0);
  assign dataCache_2_io_cpu_flush_payload_lineId = _zz_io_cpu_flush_payload_lineId[5:0];
  assign dataCache_2_io_cpu_flush_isStall = (dataCache_2_io_cpu_flush_valid && (! dataCache_2_io_cpu_flush_ready));
  assign when_DBusCachedPlugin_l398 = (dataCache_2_io_cpu_flush_isStall || dataCache_2_io_cpu_execute_haltIt);
  always @(*) begin
    dataCache_2_io_cpu_execute_args_isLrsc = 1'b0;
    if(execute_MEMORY_LRSC) begin
      dataCache_2_io_cpu_execute_args_isLrsc = 1'b1;
    end
  end

  assign dataCache_2_io_cpu_execute_args_amoCtrl_alu = execute_INSTRUCTION[31 : 29];
  assign dataCache_2_io_cpu_execute_args_amoCtrl_swap = execute_INSTRUCTION[27];
  assign when_DBusCachedPlugin_l414 = (dataCache_2_io_cpu_execute_refilling && execute_arbitration_isValid);
  assign when_DBusCachedPlugin_l427 = ((execute_arbitration_isValid && execute_MEMORY_FENCE_WR) && dataCache_2_io_cpu_writesPending);
  assign DBusCachedPlugin_writesPending = dataCache_2_io_cpu_writesPending;
  assign dataCache_2_io_cpu_memory_isValid = (memory_arbitration_isValid && memory_MEMORY_ENABLE);
  assign DBusCachedPlugin_mmuBus_cmd_0_isValid = dataCache_2_io_cpu_memory_isValid;
  assign DBusCachedPlugin_mmuBus_cmd_0_isStuck = memory_arbitration_isStuck;
  assign DBusCachedPlugin_mmuBus_cmd_0_virtualAddress = memory_MEMORY_VIRTUAL_ADDRESS;
  assign DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign DBusCachedPlugin_mmuBus_end = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  always @(*) begin
    dataCache_2_io_cpu_memory_mmuRsp_isIoAccess = DBusCachedPlugin_mmuBus_rsp_isIoAccess;
    if(when_DBusCachedPlugin_l476) begin
      dataCache_2_io_cpu_memory_mmuRsp_isIoAccess = 1'b1;
    end
  end

  assign when_DBusCachedPlugin_l476 = (1'b0 && (! dataCache_2_io_cpu_memory_isWrite));
  assign DBusCachedPlugin_trigger_valid = (((memory_arbitration_isValid && (! memory_arbitration_isStuck)) && (! memory_arbitration_isFlushed)) && memory_MEMORY_ENABLE);
  assign DBusCachedPlugin_trigger_load = (! memory_MEMORY_WR);
  assign DBusCachedPlugin_trigger_store = memory_MEMORY_WR;
  assign DBusCachedPlugin_trigger_size = memory_INSTRUCTION[13 : 12];
  assign DBusCachedPlugin_trigger_virtual = memory_REGFILE_WRITE_DATA;
  assign DBusCachedPlugin_trigger_writeData = memory_MEMORY_STORE_DATA_RF;
  assign DBusCachedPlugin_trigger_readData = 32'h0;
  assign DBusCachedPlugin_trigger_readDataValid = 1'b0;
  assign DBusCachedPlugin_trigger_dpc = memory_PC;
  always @(*) begin
    dataCache_2_io_cpu_writeBack_isValid = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
    if(writeBack_arbitration_haltByOther) begin
      dataCache_2_io_cpu_writeBack_isValid = 1'b0;
    end
  end

  assign dataCache_2_io_cpu_writeBack_isUser = (CsrPlugin_privilege == 2'b00);
  assign dataCache_2_io_cpu_writeBack_address = writeBack_REGFILE_WRITE_DATA;
  always @(*) begin
    dataCache_2_io_cpu_writeBack_storeData[31 : 0] = writeBack_MEMORY_STORE_DATA_RF;
    dataCache_2_io_cpu_writeBack_storeData[63 : 32] = writeBack_MEMORY_STORE_DATA_RF;
    if(DBusBypass0_cond) begin
      dataCache_2_io_cpu_writeBack_storeData[63 : 0] = DBusBypass0_value;
    end
  end

  assign _zz_io_cpu_writeBack_fence_SW = writeBack_INSTRUCTION[31 : 20];
  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SW = _zz_io_cpu_writeBack_fence_SW[0];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SW = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SW = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SR = _zz_io_cpu_writeBack_fence_SW[1];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SR = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SR = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SO = _zz_io_cpu_writeBack_fence_SW[2];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SO = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SO = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_SI = _zz_io_cpu_writeBack_fence_SW[3];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_SI = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_SI = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PW = _zz_io_cpu_writeBack_fence_SW[4];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PW = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PW = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PR = _zz_io_cpu_writeBack_fence_SW[5];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PR = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PR = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PO = _zz_io_cpu_writeBack_fence_SW[6];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PO = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PO = 1'b0;
    end
  end

  always @(*) begin
    dataCache_2_io_cpu_writeBack_fence_PI = _zz_io_cpu_writeBack_fence_SW[7];
    if(writeBack_DBusCachedPlugin_fence_aquire) begin
      dataCache_2_io_cpu_writeBack_fence_PI = 1'b1;
    end
    if(when_DBusCachedPlugin_l531) begin
      dataCache_2_io_cpu_writeBack_fence_PI = 1'b0;
    end
  end

  assign dataCache_2_io_cpu_writeBack_fence_FM = _zz_io_cpu_writeBack_fence_SW[11 : 8];
  always @(*) begin
    writeBack_DBusCachedPlugin_fence_aquire = 1'b0;
    if(when_DBusCachedPlugin_l518) begin
      if(writeBack_MEMORY_LRSC) begin
        writeBack_DBusCachedPlugin_fence_aquire = 1'b1;
      end
      if(writeBack_MEMORY_AMO) begin
        writeBack_DBusCachedPlugin_fence_aquire = 1'b1;
      end
    end
  end

  assign when_DBusCachedPlugin_l518 = (writeBack_MEMORY_ENABLE && writeBack_INSTRUCTION[26]);
  assign when_DBusCachedPlugin_l531 = ((! writeBack_MEMORY_FENCE) || (! writeBack_arbitration_isFiring));
  assign when_DBusCachedPlugin_l535 = (writeBack_arbitration_isValid && (writeBack_MEMORY_FENCE || writeBack_DBusCachedPlugin_fence_aquire));
  always @(*) begin
    DBusCachedPlugin_redoBranch_valid = 1'b0;
    if(when_DBusCachedPlugin_l552) begin
      if(dataCache_2_io_cpu_redo) begin
        DBusCachedPlugin_redoBranch_valid = 1'b1;
      end
    end
  end

  assign DBusCachedPlugin_redoBranch_payload = writeBack_PC;
  always @(*) begin
    DBusCachedPlugin_exceptionBus_valid = 1'b0;
    if(when_DBusCachedPlugin_l552) begin
      if(dataCache_2_io_cpu_writeBack_accessError) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_2_io_cpu_writeBack_mmuException) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_2_io_cpu_writeBack_unalignedAccess) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_2_io_cpu_redo) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b0;
      end
    end
  end

  assign DBusCachedPlugin_exceptionBus_payload_badAddr = writeBack_REGFILE_WRITE_DATA;
  always @(*) begin
    DBusCachedPlugin_exceptionBus_payload_code = 4'bxxxx;
    if(when_DBusCachedPlugin_l552) begin
      if(dataCache_2_io_cpu_writeBack_accessError) begin
        DBusCachedPlugin_exceptionBus_payload_code = {1'd0, _zz_DBusCachedPlugin_exceptionBus_payload_code};
      end
      if(dataCache_2_io_cpu_writeBack_mmuException) begin
        DBusCachedPlugin_exceptionBus_payload_code = (writeBack_MEMORY_WR ? 4'b1111 : 4'b1101);
      end
      if(dataCache_2_io_cpu_writeBack_unalignedAccess) begin
        DBusCachedPlugin_exceptionBus_payload_code = {1'd0, _zz_DBusCachedPlugin_exceptionBus_payload_code_1};
      end
    end
  end

  assign when_DBusCachedPlugin_l552 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign when_DBusCachedPlugin_l572 = (dataCache_2_io_cpu_writeBack_isValid && dataCache_2_io_cpu_writeBack_haltIt);
  assign writeBack_DBusCachedPlugin_rspData = dataCache_2_io_cpu_writeBack_data;
  assign writeBack_DBusCachedPlugin_rspSplits_0 = writeBack_DBusCachedPlugin_rspData[7 : 0];
  assign writeBack_DBusCachedPlugin_rspSplits_1 = writeBack_DBusCachedPlugin_rspData[15 : 8];
  assign writeBack_DBusCachedPlugin_rspSplits_2 = writeBack_DBusCachedPlugin_rspData[23 : 16];
  assign writeBack_DBusCachedPlugin_rspSplits_3 = writeBack_DBusCachedPlugin_rspData[31 : 24];
  assign writeBack_DBusCachedPlugin_rspSplits_4 = writeBack_DBusCachedPlugin_rspData[39 : 32];
  assign writeBack_DBusCachedPlugin_rspSplits_5 = writeBack_DBusCachedPlugin_rspData[47 : 40];
  assign writeBack_DBusCachedPlugin_rspSplits_6 = writeBack_DBusCachedPlugin_rspData[55 : 48];
  assign writeBack_DBusCachedPlugin_rspSplits_7 = writeBack_DBusCachedPlugin_rspData[63 : 56];
  always @(*) begin
    writeBack_DBusCachedPlugin_rspShifted[7 : 0] = _zz_writeBack_DBusCachedPlugin_rspShifted;
    writeBack_DBusCachedPlugin_rspShifted[15 : 8] = _zz_writeBack_DBusCachedPlugin_rspShifted_2;
    writeBack_DBusCachedPlugin_rspShifted[23 : 16] = _zz_writeBack_DBusCachedPlugin_rspShifted_4;
    writeBack_DBusCachedPlugin_rspShifted[31 : 24] = _zz_writeBack_DBusCachedPlugin_rspShifted_6;
    writeBack_DBusCachedPlugin_rspShifted[39 : 32] = writeBack_DBusCachedPlugin_rspSplits_4;
    writeBack_DBusCachedPlugin_rspShifted[47 : 40] = writeBack_DBusCachedPlugin_rspSplits_5;
    writeBack_DBusCachedPlugin_rspShifted[55 : 48] = writeBack_DBusCachedPlugin_rspSplits_6;
    writeBack_DBusCachedPlugin_rspShifted[63 : 56] = writeBack_DBusCachedPlugin_rspSplits_7;
  end

  always @(*) begin
    writeBack_DBusCachedPlugin_rspRf = writeBack_DBusCachedPlugin_rspShifted[31 : 0];
    if(when_DBusCachedPlugin_l589) begin
      writeBack_DBusCachedPlugin_rspRf = {31'd0, _zz_writeBack_DBusCachedPlugin_rspRf};
    end
  end

  assign when_DBusCachedPlugin_l589 = (writeBack_MEMORY_LRSC && writeBack_MEMORY_WR);
  assign switch_Misc_l241_2 = writeBack_INSTRUCTION[13 : 12];
  assign _zz_writeBack_DBusCachedPlugin_rspFormated = (writeBack_DBusCachedPlugin_rspRf[7] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[31] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[30] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[29] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[28] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[27] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[26] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[25] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[24] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[23] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[22] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[21] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[20] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[19] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[18] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[17] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[16] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[15] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[14] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[13] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[12] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[11] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[10] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[9] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[8] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[7 : 0] = writeBack_DBusCachedPlugin_rspRf[7 : 0];
  end

  assign _zz_writeBack_DBusCachedPlugin_rspFormated_2 = (writeBack_DBusCachedPlugin_rspRf[15] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[31] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[30] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[29] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[28] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[27] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[26] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[25] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[24] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[23] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[22] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[21] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[20] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[19] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[18] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[17] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[16] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[15 : 0] = writeBack_DBusCachedPlugin_rspRf[15 : 0];
  end

  always @(*) begin
    case(switch_Misc_l241_2)
      2'b00 : begin
        writeBack_DBusCachedPlugin_rspFormated = _zz_writeBack_DBusCachedPlugin_rspFormated_1;
      end
      2'b01 : begin
        writeBack_DBusCachedPlugin_rspFormated = _zz_writeBack_DBusCachedPlugin_rspFormated_3;
      end
      default : begin
        writeBack_DBusCachedPlugin_rspFormated = writeBack_DBusCachedPlugin_rspRf;
      end
    endcase
  end

  assign when_DBusCachedPlugin_l599 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_1 = ((decode_INSTRUCTION & 32'h00007054) == 32'h00001004);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_2 = ((decode_INSTRUCTION & 32'h00004050) == 32'h00004050);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_3 = ((decode_INSTRUCTION & 32'h00000014) == 32'h00000014);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_4 = ((decode_INSTRUCTION & 32'h00000058) == 32'h0);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_5 = ((decode_INSTRUCTION & 32'h00000070) == 32'h00000020);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_6 = ((decode_INSTRUCTION & 32'h00002004) == 32'h00000004);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_7 = ((decode_INSTRUCTION & 32'h00000008) == 32'h00000008);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_8 = ((decode_INSTRUCTION & 32'h90000010) == 32'h80000010);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_9 = ((decode_INSTRUCTION & 32'h0000000c) == 32'h00000004);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_10 = ((decode_INSTRUCTION & 32'h0000004c) == 32'h00000008);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_11 = ((decode_INSTRUCTION & 32'h00001000) == 32'h0);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_12 = ((decode_INSTRUCTION & 32'h00000020) == 32'h00000020);
  assign _zz_decode_CfuPlugin_CFU_ENABLE_13 = ((decode_INSTRUCTION & 32'hc0000010) == 32'h40000010);
  assign _zz_decode_CfuPlugin_CFU_ENABLE = {(|((decode_INSTRUCTION & 32'h02007054) == 32'h00005010)),{(|{(_zz__zz_decode_CfuPlugin_CFU_ENABLE == _zz__zz_decode_CfuPlugin_CFU_ENABLE_1),(_zz__zz_decode_CfuPlugin_CFU_ENABLE_2 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_3)}),{(|(_zz__zz_decode_CfuPlugin_CFU_ENABLE_4 == _zz__zz_decode_CfuPlugin_CFU_ENABLE_5)),{(|_zz__zz_decode_CfuPlugin_CFU_ENABLE_6),{1'b0,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_7,{_zz__zz_decode_CfuPlugin_CFU_ENABLE_8,_zz__zz_decode_CfuPlugin_CFU_ENABLE_13}}}}}}};
  assign _zz_decode_SRC1_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[3 : 2];
  assign _zz_decode_SRC1_CTRL_1 = _zz_decode_SRC1_CTRL_2;
  assign _zz_decode_ALU_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[8 : 7];
  assign _zz_decode_ALU_CTRL_1 = _zz_decode_ALU_CTRL_2;
  assign _zz_decode_SRC2_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[10 : 9];
  assign _zz_decode_SRC2_CTRL_1 = _zz_decode_SRC2_CTRL_2;
  assign _zz_decode_ENV_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[24 : 23];
  assign _zz_decode_ENV_CTRL_1 = _zz_decode_ENV_CTRL_2;
  assign _zz_decode_BRANCH_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[26 : 25];
  assign _zz_decode_BRANCH_CTRL_1 = _zz_decode_BRANCH_CTRL_2;
  assign _zz_decode_FPU_ENABLE = _zz_decode_CfuPlugin_CFU_ENABLE[32];
  assign _zz_decode_FPU_OPCODE_2 = _zz_decode_CfuPlugin_CFU_ENABLE[38 : 35];
  assign _zz_decode_FPU_OPCODE_1 = _zz_decode_FPU_OPCODE_2;
  assign _zz_decode_FPU_FORMAT_2 = _zz_decode_CfuPlugin_CFU_ENABLE[39 : 39];
  assign _zz_decode_FPU_FORMAT_1 = _zz_decode_FPU_FORMAT_2;
  assign _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2 = _zz_decode_CfuPlugin_CFU_ENABLE[43 : 43];
  assign _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1 = _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_2;
  assign _zz_decode_ALU_BITWISE_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[45 : 44];
  assign _zz_decode_ALU_BITWISE_CTRL_1 = _zz_decode_ALU_BITWISE_CTRL_2;
  assign _zz_decode_SHIFT_CTRL_2 = _zz_decode_CfuPlugin_CFU_ENABLE[47 : 46];
  assign _zz_decode_SHIFT_CTRL_1 = _zz_decode_SHIFT_CTRL_2;
  assign decodeExceptionPort_valid = (decode_arbitration_isValid && (! decode_LEGAL_INSTRUCTION));
  assign decodeExceptionPort_payload_code = 4'b0010;
  assign decodeExceptionPort_payload_badAddr = decode_INSTRUCTION;
  assign when_RegFilePlugin_l63 = (decode_INSTRUCTION[11 : 7] == 5'h0);
  assign decode_RegFilePlugin_regFileReadAddress1 = decode_INSTRUCTION_ANTICIPATED[19 : 15];
  assign decode_RegFilePlugin_regFileReadAddress2 = decode_INSTRUCTION_ANTICIPATED[24 : 20];
  assign decode_RegFilePlugin_rs1Data = RegFilePlugin_regFile_spinal_port0;
  assign decode_RegFilePlugin_rs2Data = RegFilePlugin_regFile_spinal_port1;
  always @(*) begin
    lastStageRegFileWrite_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
    if(_zz_5) begin
      lastStageRegFileWrite_valid = 1'b1;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
    if(_zz_5) begin
      lastStageRegFileWrite_payload_address = 5'h0;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_data = _zz_decode_RS2_2;
    if(_zz_5) begin
      lastStageRegFileWrite_payload_data = 32'h0;
    end
  end

  always @(*) begin
    case(decode_SRC1_CTRL)
      Src1CtrlEnum_RS : begin
        _zz_decode_SRC1 = _zz_decode_to_execute_RS1;
      end
      Src1CtrlEnum_PC_INCREMENT : begin
        _zz_decode_SRC1 = {29'd0, _zz__zz_decode_SRC1};
      end
      Src1CtrlEnum_IMU : begin
        _zz_decode_SRC1 = {decode_INSTRUCTION[31 : 12],12'h0};
      end
      default : begin
        _zz_decode_SRC1 = {27'd0, _zz__zz_decode_SRC1_1};
      end
    endcase
  end

  assign _zz_decode_SRC2 = decode_INSTRUCTION[31];
  always @(*) begin
    _zz_decode_SRC2_1[19] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[18] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[17] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[16] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[15] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[14] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[13] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[12] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[11] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[10] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[9] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[8] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[7] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[6] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[5] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[4] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[3] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[2] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[1] = _zz_decode_SRC2;
    _zz_decode_SRC2_1[0] = _zz_decode_SRC2;
  end

  assign _zz_decode_SRC2_2 = _zz__zz_decode_SRC2_2[11];
  always @(*) begin
    _zz_decode_SRC2_3[19] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[18] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[17] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[16] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[15] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[14] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[13] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[12] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[11] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[10] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[9] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[8] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[7] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[6] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[5] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[4] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[3] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[2] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[1] = _zz_decode_SRC2_2;
    _zz_decode_SRC2_3[0] = _zz_decode_SRC2_2;
  end

  always @(*) begin
    case(decode_SRC2_CTRL)
      Src2CtrlEnum_RS : begin
        _zz_decode_SRC2_4 = _zz_decode_to_execute_RS2;
      end
      Src2CtrlEnum_IMI : begin
        _zz_decode_SRC2_4 = {_zz_decode_SRC2_1,decode_INSTRUCTION[31 : 20]};
      end
      Src2CtrlEnum_IMS : begin
        _zz_decode_SRC2_4 = {_zz_decode_SRC2_3,{decode_INSTRUCTION[31 : 25],decode_INSTRUCTION[11 : 7]}};
      end
      default : begin
        _zz_decode_SRC2_4 = _zz_decode_to_execute_PC;
      end
    endcase
  end

  always @(*) begin
    execute_SrcPlugin_addSub = _zz_execute_SrcPlugin_addSub;
    if(execute_SRC2_FORCE_ZERO) begin
      execute_SrcPlugin_addSub = execute_SRC1;
    end
  end

  assign execute_SrcPlugin_less = ((execute_SRC1[31] == execute_SRC2[31]) ? execute_SrcPlugin_addSub[31] : (execute_SRC_LESS_UNSIGNED ? execute_SRC2[31] : execute_SRC1[31]));
  always @(*) begin
    HazardSimplePlugin_src0Hazard = 1'b0;
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l48) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l48_1) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l48_2) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l105) begin
      HazardSimplePlugin_src0Hazard = 1'b0;
    end
  end

  always @(*) begin
    HazardSimplePlugin_src1Hazard = 1'b0;
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l51) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l51_1) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l51_2) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l108) begin
      HazardSimplePlugin_src1Hazard = 1'b0;
    end
  end

  assign HazardSimplePlugin_writeBackWrites_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
  assign HazardSimplePlugin_writeBackWrites_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
  assign HazardSimplePlugin_writeBackWrites_payload_data = _zz_decode_RS2_2;
  assign HazardSimplePlugin_addr0Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[19 : 15]);
  assign HazardSimplePlugin_addr1Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l47 = 1'b1;
  assign when_HazardSimplePlugin_l48 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58 = (1'b0 || (! when_HazardSimplePlugin_l47));
  assign when_HazardSimplePlugin_l48_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_1 = (1'b0 || (! memory_BYPASSABLE_MEMORY_STAGE));
  assign when_HazardSimplePlugin_l48_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_2 = (1'b0 || (! execute_BYPASSABLE_EXECUTE_STAGE));
  assign when_HazardSimplePlugin_l105 = (! decode_RS1_USE);
  assign when_HazardSimplePlugin_l108 = (! decode_RS2_USE);
  assign when_HazardSimplePlugin_l113 = (decode_arbitration_isValid && (HazardSimplePlugin_src0Hazard || HazardSimplePlugin_src1Hazard));
  always @(*) begin
    when_CsrPlugin_l836 = 1'b0;
    if(when_CsrPlugin_l1534) begin
      when_CsrPlugin_l836 = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_privilege = _zz_CsrPlugin_privilege;
    if(CsrPlugin_forceMachineWire) begin
      CsrPlugin_privilege = 2'b11;
    end
  end

  assign debugMode = (! CsrPlugin_running);
  assign when_CsrPlugin_l729 = (! CsrPlugin_running);
  always @(*) begin
    debugBus_resume_rsp_valid = 1'b0;
    if(CsrPlugin_doResume) begin
      debugBus_resume_rsp_valid = 1'b1;
    end
  end

  assign debugBus_running = CsrPlugin_running;
  assign debugBus_halted = (! CsrPlugin_running);
  assign debugBus_unavailable = systemCd_logic_outputReset_buffercc_io_dataOut;
  assign debugBus_haveReset = _zz_debugBus_haveReset;
  assign CsrPlugin_enterHalt = ((! CsrPlugin_running_aheadValue) && CsrPlugin_running_aheadValue_regNext);
  assign when_CsrPlugin_l747 = ((debugBus_haltReq && debugBus_running) && (! debugMode));
  assign CsrPlugin_forceResume = 1'b0;
  assign CsrPlugin_doResume = (CsrPlugin_forceResume || _zz_CsrPlugin_doResume);
  always @(*) begin
    CsrPlugin_timeout_stateRise = 1'b0;
    if(CsrPlugin_timeout_counter_willOverflow) begin
      CsrPlugin_timeout_stateRise = (! CsrPlugin_timeout_state);
    end
    if(when_CsrPlugin_l753) begin
      CsrPlugin_timeout_stateRise = 1'b0;
    end
    if(CsrPlugin_inject_cmd_valid) begin
      CsrPlugin_timeout_stateRise = 1'b0;
    end
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
        CsrPlugin_timeout_stateRise = 1'b0;
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_timeout_counter_willClear = 1'b0;
    if(when_CsrPlugin_l753) begin
      CsrPlugin_timeout_counter_willClear = 1'b1;
    end
    if(CsrPlugin_inject_cmd_valid) begin
      CsrPlugin_timeout_counter_willClear = 1'b1;
    end
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
        CsrPlugin_timeout_counter_willClear = 1'b1;
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
      end
      default : begin
      end
    endcase
  end

  assign CsrPlugin_timeout_counter_willOverflowIfInc = (CsrPlugin_timeout_counter_value == 3'b110);
  assign CsrPlugin_timeout_counter_willOverflow = (CsrPlugin_timeout_counter_willOverflowIfInc && CsrPlugin_timeout_counter_willIncrement);
  always @(*) begin
    if(CsrPlugin_timeout_counter_willOverflow) begin
      CsrPlugin_timeout_counter_valueNext = 3'b000;
    end else begin
      CsrPlugin_timeout_counter_valueNext = (CsrPlugin_timeout_counter_value + _zz_CsrPlugin_timeout_counter_valueNext);
    end
    if(CsrPlugin_timeout_counter_willClear) begin
      CsrPlugin_timeout_counter_valueNext = 3'b000;
    end
  end

  assign CsrPlugin_timeout_counter_willIncrement = 1'b1;
  assign when_CsrPlugin_l753 = (|{writeBack_arbitration_isValid,{memory_arbitration_isValid,execute_arbitration_isValid}});
  always @(*) begin
    _zz_debugBus_hartToDm_valid = 1'b0;
    if(execute_CsrPlugin_csr_1972) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_debugBus_hartToDm_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    debugBus_hartToDm_valid = _zz_debugBus_hartToDm_valid;
    if(fpuAccess_readDataValid) begin
      debugBus_hartToDm_valid = 1'b1;
    end
  end

  always @(*) begin
    debugBus_hartToDm_payload_address = 4'b0000;
    if(fpuAccess_readDataValid) begin
      debugBus_hartToDm_payload_address = {3'd0, fpuAccess_readDataChunk};
    end
  end

  always @(*) begin
    debugBus_hartToDm_payload_data = execute_SRC1;
    if(fpuAccess_readDataValid) begin
      debugBus_hartToDm_payload_data = fpuAccess_readData;
    end
  end

  assign when_CsrPlugin_l768 = (debugBus_dmToHart_valid && (debugBus_dmToHart_payload_op == DebugDmToHartOp_DATA));
  assign _zz_6 = ({1'd0,1'b1} <<< _zz__zz_6);
  assign CsrPlugin_inject_cmd_valid = (debugBus_dmToHart_valid && (((debugBus_dmToHart_payload_op == DebugDmToHartOp_EXECUTE) || (debugBus_dmToHart_payload_op == DebugDmToHartOp_REG_READ)) || (debugBus_dmToHart_payload_op == DebugDmToHartOp_REG_WRITE)));
  assign CsrPlugin_inject_cmd_payload_op = debugBus_dmToHart_payload_op;
  assign CsrPlugin_inject_cmd_payload_address = debugBus_dmToHart_payload_address;
  assign CsrPlugin_inject_cmd_payload_data = debugBus_dmToHart_payload_data;
  assign CsrPlugin_inject_cmd_payload_size = debugBus_dmToHart_payload_size;
  assign CsrPlugin_inject_cmd_toStream_valid = CsrPlugin_inject_cmd_valid;
  assign CsrPlugin_inject_cmd_toStream_payload_op = CsrPlugin_inject_cmd_payload_op;
  assign CsrPlugin_inject_cmd_toStream_payload_address = CsrPlugin_inject_cmd_payload_address;
  assign CsrPlugin_inject_cmd_toStream_payload_data = CsrPlugin_inject_cmd_payload_data;
  assign CsrPlugin_inject_cmd_toStream_payload_size = CsrPlugin_inject_cmd_payload_size;
  always @(*) begin
    CsrPlugin_inject_cmd_toStream_ready = CsrPlugin_inject_buffer_ready;
    if(when_Stream_l375_1) begin
      CsrPlugin_inject_cmd_toStream_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! CsrPlugin_inject_buffer_valid);
  assign CsrPlugin_inject_buffer_valid = CsrPlugin_inject_cmd_toStream_rValid;
  assign CsrPlugin_inject_buffer_payload_op = CsrPlugin_inject_cmd_toStream_rData_op;
  assign CsrPlugin_inject_buffer_payload_address = CsrPlugin_inject_cmd_toStream_rData_address;
  assign CsrPlugin_inject_buffer_payload_data = CsrPlugin_inject_cmd_toStream_rData_data;
  assign CsrPlugin_inject_buffer_payload_size = CsrPlugin_inject_cmd_toStream_rData_size;
  assign CsrPlugin_injectionPort_valid = (CsrPlugin_inject_buffer_valid && (CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_EXECUTE));
  assign CsrPlugin_injectionPort_payload = CsrPlugin_inject_buffer_payload_data;
  assign CsrPlugin_injectionPort_fire = (CsrPlugin_injectionPort_valid && CsrPlugin_injectionPort_ready);
  always @(*) begin
    CsrPlugin_inject_buffer_ready = CsrPlugin_injectionPort_fire;
    if(fpuAccess_done) begin
      CsrPlugin_inject_buffer_ready = 1'b1;
    end
  end

  assign fpuAccess_start = (CsrPlugin_inject_buffer_valid && ((CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_REG_READ) || (CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_REG_WRITE)));
  assign fpuAccess_regId = CsrPlugin_inject_buffer_payload_address;
  assign fpuAccess_write = (CsrPlugin_inject_buffer_payload_op == DebugDmToHartOp_REG_WRITE);
  assign fpuAccess_writeData = {CsrPlugin_dataCsrw_value_1,CsrPlugin_dataCsrw_value_0};
  assign fpuAccess_size = CsrPlugin_inject_buffer_payload_size;
  assign debugBus_regSuccess = fpuAccess_done;
  assign when_CsrPlugin_l804 = (CsrPlugin_inject_cmd_valid && (debugBus_dmToHart_payload_op == DebugDmToHartOp_EXECUTE));
  assign when_CsrPlugin_l804_1 = (((debugBus_exception || debugBus_commit) || debugBus_ebreak) || debugBus_redo);
  assign debugBus_redo = (CsrPlugin_inject_pending && CsrPlugin_timeout_state);
  assign CsrPlugin_dcsr_nmip = 1'b0;
  assign CsrPlugin_dcsr_mprven = 1'b1;
  assign CsrPlugin_dcsr_xdebugver = 4'b0100;
  assign CsrPlugin_dcsr_stepLogic_wantExit = 1'b0;
  always @(*) begin
    CsrPlugin_dcsr_stepLogic_wantStart = 1'b0;
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
      end
      default : begin
        CsrPlugin_dcsr_stepLogic_wantStart = 1'b1;
      end
    endcase
  end

  assign CsrPlugin_dcsr_stepLogic_wantKill = 1'b0;
  always @(*) begin
    CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_stateReg;
    case(CsrPlugin_dcsr_stepLogic_stateReg)
      CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
        if(when_CsrPlugin_l830) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_SINGLE;
        end
      end
      CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
        if(when_CsrPlugin_l836) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1;
        end
        if(decode_arbitration_isFiring) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1;
        end
      end
      CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
        if(when_CsrPlugin_l848) begin
          CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_SINGLE;
        end
      end
      default : begin
      end
    endcase
    if(CsrPlugin_enterHalt) begin
      CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_IDLE;
    end
    if(CsrPlugin_dcsr_stepLogic_wantStart) begin
      CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_IDLE;
    end
    if(CsrPlugin_dcsr_stepLogic_wantKill) begin
      CsrPlugin_dcsr_stepLogic_stateNext = CsrPlugin_dcsr_stepLogic_enumDef_BOOT;
    end
  end

  assign when_CsrPlugin_l830 = (CsrPlugin_dcsr_step && debugBus_resume_rsp_valid);
  assign when_CsrPlugin_l848 = ((! CsrPlugin_doHalt) && CsrPlugin_timeout_state);
  assign when_CsrPlugin_l880 = ((debugMode || CsrPlugin_dcsr_step) || debugBus_haltReq);
  assign CsrPlugin_misa_base = 2'b01;
  assign CsrPlugin_misa_extensions = 26'h000112d;
  assign _zz_when_CsrPlugin_l1446 = (CsrPlugin_mip_MTIP && CsrPlugin_mie_MTIE);
  assign _zz_when_CsrPlugin_l1446_1 = (CsrPlugin_mip_MSIP && CsrPlugin_mie_MSIE);
  assign _zz_when_CsrPlugin_l1446_2 = (CsrPlugin_mip_MEIP && CsrPlugin_mie_MEIE);
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped = 2'b11;
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege = ((CsrPlugin_privilege < CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped) ? CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped : CsrPlugin_privilege);
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code = {decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid};
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1[0];
  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_decode = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_execute = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_memory = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
    if(memory_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
    if(DBusCachedPlugin_exceptionBus_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b1;
    end
    if(writeBack_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b0;
    end
  end

  assign when_CsrPlugin_l1403 = (! decode_arbitration_isStuck);
  assign when_CsrPlugin_l1403_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1403_2 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l1403_3 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l1416 = (|{CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValids_memory,{CsrPlugin_exceptionPortCtrl_exceptionValids_execute,CsrPlugin_exceptionPortCtrl_exceptionValids_decode}}});
  assign CsrPlugin_exceptionPendings_0 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  assign CsrPlugin_exceptionPendings_1 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  assign CsrPlugin_exceptionPendings_2 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  assign CsrPlugin_exceptionPendings_3 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  assign when_CsrPlugin_l1440 = (CsrPlugin_mstatus_MIE || (CsrPlugin_privilege < 2'b11));
  assign when_CsrPlugin_l1446 = ((_zz_when_CsrPlugin_l1446 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l1446_1 = ((_zz_when_CsrPlugin_l1446_1 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l1446_2 = ((_zz_when_CsrPlugin_l1446_2 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l1459 = (CsrPlugin_dcsr_step && (! CsrPlugin_dcsr_stepie));
  assign CsrPlugin_exception = (CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack && CsrPlugin_allowException);
  assign CsrPlugin_lastStageWasWfi = 1'b0;
  assign CsrPlugin_pipelineLiberator_active = ((CsrPlugin_interrupt_valid && CsrPlugin_allowInterrupts) && decode_arbitration_isValid);
  assign when_CsrPlugin_l1479 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1479_1 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l1479_2 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l1484 = ((! CsrPlugin_pipelineLiberator_active) || decode_arbitration_removeIt);
  always @(*) begin
    CsrPlugin_pipelineLiberator_done = CsrPlugin_pipelineLiberator_pcValids_2;
    if(when_CsrPlugin_l1490) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
    if(CsrPlugin_hadException) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
  end

  assign when_CsrPlugin_l1490 = (|{CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory,CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute}});
  assign CsrPlugin_interruptJump = ((CsrPlugin_interrupt_valid && CsrPlugin_pipelineLiberator_done) && CsrPlugin_allowInterrupts);
  assign debugBus_commit = (debugMode && writeBack_arbitration_isFiring);
  always @(*) begin
    debugBus_exception = (debugMode && CsrPlugin_hadException);
    if(when_CsrPlugin_l1534) begin
      if(!when_CsrPlugin_l1542) begin
        if(!when_CsrPlugin_l1572) begin
          debugBus_exception = (! CsrPlugin_trapCauseEbreakDebug);
        end
      end
    end
  end

  always @(*) begin
    debugBus_ebreak = 1'b0;
    if(when_CsrPlugin_l1534) begin
      if(!when_CsrPlugin_l1542) begin
        if(!when_CsrPlugin_l1572) begin
          debugBus_ebreak = CsrPlugin_trapCauseEbreakDebug;
        end
      end
    end
  end

  always @(*) begin
    CsrPlugin_targetPrivilege = CsrPlugin_interrupt_targetPrivilege;
    if(CsrPlugin_hadException) begin
      CsrPlugin_targetPrivilege = CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
    end
  end

  always @(*) begin
    CsrPlugin_trapCause = CsrPlugin_interrupt_code;
    if(CsrPlugin_hadException) begin
      CsrPlugin_trapCause = CsrPlugin_exceptionPortCtrl_exceptionContext_code;
    end
  end

  always @(*) begin
    CsrPlugin_trapCauseEbreakDebug = 1'b0;
    if(CsrPlugin_hadException) begin
      if(when_CsrPlugin_l1517) begin
        if(debugMode) begin
          CsrPlugin_trapCauseEbreakDebug = 1'b1;
        end
        if(when_CsrPlugin_l1519) begin
          CsrPlugin_trapCauseEbreakDebug = 1'b1;
        end
      end
    end
  end

  assign when_CsrPlugin_l1517 = (CsrPlugin_exceptionPortCtrl_exceptionContext_code == 4'b0011);
  assign when_CsrPlugin_l1519 = ((CsrPlugin_privilege == 2'b11) && CsrPlugin_dcsr_ebreakm);
  always @(*) begin
    CsrPlugin_xtvec_mode = 2'bxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_mode = CsrPlugin_mtvec_mode;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_xtvec_base = 30'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_base = CsrPlugin_mtvec_base;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_trapEnterDebug = 1'b0;
    if(when_CsrPlugin_l1533) begin
      CsrPlugin_trapEnterDebug = 1'b1;
    end
  end

  assign when_CsrPlugin_l1533 = (((CsrPlugin_doHalt || CsrPlugin_trapCauseEbreakDebug) || ((! CsrPlugin_hadException) && CsrPlugin_doHalt)) || (! CsrPlugin_running));
  assign when_CsrPlugin_l1534 = (CsrPlugin_hadException || CsrPlugin_interruptJump);
  assign when_CsrPlugin_l1542 = (! CsrPlugin_trapEnterDebug);
  assign when_CsrPlugin_l1572 = (! debugMode);
  assign when_CsrPlugin_l1600 = (writeBack_arbitration_isValid && (writeBack_ENV_CTRL == EnvCtrlEnum_XRET));
  assign switch_CsrPlugin_l1604 = writeBack_INSTRUCTION[29 : 28];
  assign when_CsrPlugin_l1612 = (CsrPlugin_mstatus_MPP < 2'b11);
  assign contextSwitching = CsrPlugin_jumpInterface_valid;
  assign when_CsrPlugin_l1671 = (|{(writeBack_arbitration_isValid && (writeBack_ENV_CTRL == EnvCtrlEnum_XRET)),{(memory_arbitration_isValid && (memory_ENV_CTRL == EnvCtrlEnum_XRET)),(execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_XRET))}});
  assign execute_CsrPlugin_blockedBySideEffects = ((|{writeBack_arbitration_isValid,memory_arbitration_isValid}) || 1'b0);
  always @(*) begin
    execute_CsrPlugin_illegalAccess = 1'b1;
    if(execute_CsrPlugin_csr_1972) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_1969) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_1968) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_3857) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3858) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3859) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3860) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_769) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_768) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_836) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_772) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_773) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_833) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_832) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_834) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_835) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_2) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_1) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_256) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(CsrPlugin_csrMapping_allowCsrSignal) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(when_CsrPlugin_l1863) begin
      execute_CsrPlugin_illegalAccess = 1'b1;
    end
    if(when_CsrPlugin_l1869) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_illegalInstruction = 1'b0;
    if(when_CsrPlugin_l1691) begin
      if(when_CsrPlugin_l1692) begin
        execute_CsrPlugin_illegalInstruction = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrPlugin_selfException_valid = 1'b0;
    if(when_CsrPlugin_l1684) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
    if(when_CsrPlugin_l1699) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
    if(when_CsrPlugin_l1709) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_selfException_payload_code = 4'bxxxx;
    if(when_CsrPlugin_l1684) begin
      CsrPlugin_selfException_payload_code = 4'b0010;
    end
    if(when_CsrPlugin_l1699) begin
      case(CsrPlugin_privilege)
        2'b00 : begin
          CsrPlugin_selfException_payload_code = 4'b1000;
        end
        default : begin
          CsrPlugin_selfException_payload_code = 4'b1011;
        end
      endcase
    end
    if(when_CsrPlugin_l1709) begin
      CsrPlugin_selfException_payload_code = 4'b0011;
    end
  end

  assign CsrPlugin_selfException_payload_badAddr = execute_INSTRUCTION;
  assign when_CsrPlugin_l1684 = (execute_CsrPlugin_illegalAccess || execute_CsrPlugin_illegalInstruction);
  assign when_CsrPlugin_l1691 = (execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_XRET));
  assign when_CsrPlugin_l1692 = (CsrPlugin_privilege < execute_INSTRUCTION[29 : 28]);
  assign when_CsrPlugin_l1699 = (execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_ECALL));
  assign when_CsrPlugin_l1709 = ((execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_EBREAK)) && CsrPlugin_allowEbreakException);
  always @(*) begin
    execute_CsrPlugin_writeInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_WRITE_OPCODE);
    if(when_CsrPlugin_l1863) begin
      execute_CsrPlugin_writeInstruction = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_readInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_READ_OPCODE);
    if(when_CsrPlugin_l1863) begin
      execute_CsrPlugin_readInstruction = 1'b0;
    end
  end

  assign execute_CsrPlugin_writeEnable = (execute_CsrPlugin_writeInstruction && (! execute_arbitration_isStuck));
  assign execute_CsrPlugin_readEnable = (execute_CsrPlugin_readInstruction && (! execute_arbitration_isStuck));
  assign CsrPlugin_csrMapping_hazardFree = (! execute_CsrPlugin_blockedBySideEffects);
  assign execute_CsrPlugin_readToWriteData = CsrPlugin_csrMapping_readDataSignal;
  assign switch_Misc_l241_3 = execute_INSTRUCTION[13];
  always @(*) begin
    case(switch_Misc_l241_3)
      1'b0 : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = execute_SRC1;
      end
      default : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = (execute_INSTRUCTION[12] ? (execute_CsrPlugin_readToWriteData & (~ execute_SRC1)) : (execute_CsrPlugin_readToWriteData | execute_SRC1));
      end
    endcase
  end

  assign CsrPlugin_csrMapping_writeDataSignal = _zz_CsrPlugin_csrMapping_writeDataSignal;
  assign when_CsrPlugin_l1731 = (execute_arbitration_isValid && execute_IS_CSR);
  assign when_CsrPlugin_l1735 = (execute_arbitration_isValid && (execute_IS_CSR || 1'b0));
  assign execute_CsrPlugin_csrAddress = execute_INSTRUCTION[31 : 20];
  assign execute_BranchPlugin_eq = (execute_SRC1 == execute_SRC2);
  assign switch_Misc_l241_4 = execute_INSTRUCTION[14 : 12];
  always @(*) begin
    case(switch_Misc_l241_4)
      3'b000 : begin
        _zz_execute_BRANCH_DO = execute_BranchPlugin_eq;
      end
      3'b001 : begin
        _zz_execute_BRANCH_DO = (! execute_BranchPlugin_eq);
      end
      3'b101 : begin
        _zz_execute_BRANCH_DO = (! execute_SRC_LESS);
      end
      3'b111 : begin
        _zz_execute_BRANCH_DO = (! execute_SRC_LESS);
      end
      default : begin
        _zz_execute_BRANCH_DO = execute_SRC_LESS;
      end
    endcase
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : begin
        _zz_execute_BRANCH_DO_1 = 1'b0;
      end
      BranchCtrlEnum_JAL : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      BranchCtrlEnum_JALR : begin
        _zz_execute_BRANCH_DO_1 = 1'b1;
      end
      default : begin
        _zz_execute_BRANCH_DO_1 = _zz_execute_BRANCH_DO;
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src1 = ((execute_BRANCH_CTRL == BranchCtrlEnum_JALR) ? execute_RS1 : execute_PC);
  assign _zz_execute_BranchPlugin_branch_src2 = _zz__zz_execute_BranchPlugin_branch_src2[19];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_1[10] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[9] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[8] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[7] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[6] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[5] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[4] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[3] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[2] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[1] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[0] = _zz_execute_BranchPlugin_branch_src2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_2 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_3[19] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[18] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[17] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[16] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[15] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[14] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[13] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[12] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[11] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[10] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[9] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[8] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[7] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[6] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[5] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[4] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[3] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[2] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[1] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[0] = _zz_execute_BranchPlugin_branch_src2_2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_4 = _zz__zz_execute_BranchPlugin_branch_src2_4[11];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_5[18] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[17] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[16] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[15] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[14] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[13] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[12] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[11] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[10] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[9] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[8] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[7] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[6] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[5] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[4] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[3] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[2] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[1] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[0] = _zz_execute_BranchPlugin_branch_src2_4;
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_JAL : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_1,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]}},1'b0};
      end
      BranchCtrlEnum_JALR : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {_zz_execute_BranchPlugin_branch_src2_3,execute_INSTRUCTION[31 : 20]};
      end
      default : begin
        _zz_execute_BranchPlugin_branch_src2_6 = {{_zz_execute_BranchPlugin_branch_src2_5,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]}},1'b0};
      end
    endcase
  end

  assign execute_BranchPlugin_branch_src2 = _zz_execute_BranchPlugin_branch_src2_6;
  assign execute_BranchPlugin_branchAdder = (execute_BranchPlugin_branch_src1 + execute_BranchPlugin_branch_src2);
  assign BranchPlugin_jumpInterface_valid = ((memory_arbitration_isValid && memory_BRANCH_DO) && (! 1'b0));
  assign BranchPlugin_jumpInterface_payload = memory_BRANCH_CALC;
  assign when_MulPlugin_l65 = ((execute_arbitration_isValid && execute_IS_MUL) && (execute_MulPlugin_delayLogic_counter != 1'b1));
  assign when_MulPlugin_l70 = ((! execute_arbitration_isStuck) || execute_arbitration_isStuckByOthers);
  assign execute_MulPlugin_a = execute_RS1;
  assign execute_MulPlugin_b = execute_RS2;
  assign switch_MulPlugin_l87 = execute_INSTRUCTION[13 : 12];
  always @(*) begin
    case(switch_MulPlugin_l87)
      2'b01 : begin
        execute_MulPlugin_aSigned = 1'b1;
      end
      2'b10 : begin
        execute_MulPlugin_aSigned = 1'b1;
      end
      default : begin
        execute_MulPlugin_aSigned = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(switch_MulPlugin_l87)
      2'b01 : begin
        execute_MulPlugin_bSigned = 1'b1;
      end
      2'b10 : begin
        execute_MulPlugin_bSigned = 1'b0;
      end
      default : begin
        execute_MulPlugin_bSigned = 1'b0;
      end
    endcase
  end

  assign execute_MulPlugin_aULow = execute_MulPlugin_a[15 : 0];
  assign execute_MulPlugin_bULow = execute_MulPlugin_b[15 : 0];
  assign execute_MulPlugin_aSLow = {1'b0,execute_MulPlugin_a[15 : 0]};
  assign execute_MulPlugin_bSLow = {1'b0,execute_MulPlugin_b[15 : 0]};
  assign execute_MulPlugin_aHigh = {(execute_MulPlugin_aSigned && execute_MulPlugin_a[31]),execute_MulPlugin_a[31 : 16]};
  assign execute_MulPlugin_bHigh = {(execute_MulPlugin_bSigned && execute_MulPlugin_b[31]),execute_MulPlugin_b[31 : 16]};
  assign writeBack_MulPlugin_result = ($signed(_zz_writeBack_MulPlugin_result) + $signed(_zz_writeBack_MulPlugin_result_1));
  assign when_MulPlugin_l147 = (writeBack_arbitration_isValid && writeBack_IS_MUL);
  assign switch_MulPlugin_l148 = writeBack_INSTRUCTION[13 : 12];
  assign memory_MulDivIterativePlugin_frontendOk = 1'b1;
  always @(*) begin
    memory_MulDivIterativePlugin_div_counter_willIncrement = 1'b0;
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l132) begin
        memory_MulDivIterativePlugin_div_counter_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    memory_MulDivIterativePlugin_div_counter_willClear = 1'b0;
    if(when_MulDivIterativePlugin_l162) begin
      memory_MulDivIterativePlugin_div_counter_willClear = 1'b1;
    end
  end

  assign memory_MulDivIterativePlugin_div_counter_willOverflowIfInc = (memory_MulDivIterativePlugin_div_counter_value == 6'h21);
  assign memory_MulDivIterativePlugin_div_counter_willOverflow = (memory_MulDivIterativePlugin_div_counter_willOverflowIfInc && memory_MulDivIterativePlugin_div_counter_willIncrement);
  always @(*) begin
    if(memory_MulDivIterativePlugin_div_counter_willOverflow) begin
      memory_MulDivIterativePlugin_div_counter_valueNext = 6'h0;
    end else begin
      memory_MulDivIterativePlugin_div_counter_valueNext = (memory_MulDivIterativePlugin_div_counter_value + _zz_memory_MulDivIterativePlugin_div_counter_valueNext);
    end
    if(memory_MulDivIterativePlugin_div_counter_willClear) begin
      memory_MulDivIterativePlugin_div_counter_valueNext = 6'h0;
    end
  end

  assign when_MulDivIterativePlugin_l126 = (memory_MulDivIterativePlugin_div_counter_value == 6'h20);
  assign when_MulDivIterativePlugin_l126_1 = (! memory_arbitration_isStuck);
  assign when_MulDivIterativePlugin_l128 = (memory_arbitration_isValid && memory_IS_DIV);
  assign when_MulDivIterativePlugin_l129 = ((! memory_MulDivIterativePlugin_frontendOk) || (! memory_MulDivIterativePlugin_div_done));
  assign when_MulDivIterativePlugin_l132 = (memory_MulDivIterativePlugin_frontendOk && (! memory_MulDivIterativePlugin_div_done));
  assign _zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted = memory_MulDivIterativePlugin_rs1[31 : 0];
  assign memory_MulDivIterativePlugin_div_stage_0_remainderShifted = {memory_MulDivIterativePlugin_accumulator[31 : 0],_zz_memory_MulDivIterativePlugin_div_stage_0_remainderShifted[31]};
  assign memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator = (memory_MulDivIterativePlugin_div_stage_0_remainderShifted - _zz_memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator);
  assign memory_MulDivIterativePlugin_div_stage_0_outRemainder = ((! memory_MulDivIterativePlugin_div_stage_0_remainderMinusDenominator[32]) ? _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder : _zz_memory_MulDivIterativePlugin_div_stage_0_outRemainder_1);
  assign memory_MulDivIterativePlugin_div_stage_0_outNumerator = _zz_memory_MulDivIterativePlugin_div_stage_0_outNumerator[31:0];
  assign when_MulDivIterativePlugin_l151 = (memory_MulDivIterativePlugin_div_counter_value == 6'h20);
  assign _zz_memory_MulDivIterativePlugin_div_result = (memory_INSTRUCTION[13] ? memory_MulDivIterativePlugin_accumulator[31 : 0] : memory_MulDivIterativePlugin_rs1[31 : 0]);
  assign when_MulDivIterativePlugin_l162 = (! memory_arbitration_isStuck);
  assign _zz_memory_MulDivIterativePlugin_rs2 = (execute_RS2[31] && execute_IS_RS2_SIGNED);
  assign _zz_memory_MulDivIterativePlugin_rs1 = (1'b0 || ((execute_IS_DIV && execute_RS1[31]) && execute_IS_RS1_SIGNED));
  always @(*) begin
    _zz_memory_MulDivIterativePlugin_rs1_1[32] = (execute_IS_RS1_SIGNED && execute_RS1[31]);
    _zz_memory_MulDivIterativePlugin_rs1_1[31 : 0] = execute_RS1;
  end

  assign FpuPlugin_port_cmd_fire = (FpuPlugin_port_cmd_valid && FpuPlugin_port_cmd_ready);
  assign FpuPlugin_port_rsp_fire = (FpuPlugin_port_rsp_valid && FpuPlugin_port_rsp_ready);
  assign FpuPlugin_hasPending = (FpuPlugin_pendings != 6'h0);
  assign when_FpuPlugin_l215 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_NV);
  assign when_FpuPlugin_l216 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_DZ);
  assign when_FpuPlugin_l217 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_OF);
  assign when_FpuPlugin_l218 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_UF);
  assign when_FpuPlugin_l219 = (FpuPlugin_port_completion_valid && FpuPlugin_port_completion_payload_flags_NX);
  assign FpuPlugin_csrActive = (execute_arbitration_isValid && execute_IS_CSR);
  assign when_FpuPlugin_l229 = (FpuPlugin_csrActive && FpuPlugin_hasPending);
  assign FpuPlugin_sd = (FpuPlugin_fs == 2'b11);
  assign when_FpuPlugin_l234 = (FpuPlugin_port_completion_valid && (FpuPlugin_port_completion_payload_written || (|{FpuPlugin_port_completion_payload_flags_NV,{FpuPlugin_port_completion_payload_flags_DZ,{FpuPlugin_port_completion_payload_flags_OF,{FpuPlugin_port_completion_payload_flags_UF,FpuPlugin_port_completion_payload_flags_NX}}}})));
  always @(*) begin
    _zz_when_FpuPlugin_l237 = 1'b0;
    if(execute_CsrPlugin_csr_2) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_when_FpuPlugin_l237 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_when_FpuPlugin_l237_1 = 1'b0;
    if(execute_CsrPlugin_csr_3) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_when_FpuPlugin_l237_1 = 1'b1;
      end
    end
  end

  always @(*) begin
    _zz_when_FpuPlugin_l237_2 = 1'b0;
    if(execute_CsrPlugin_csr_1) begin
      if(execute_CsrPlugin_writeEnable) begin
        _zz_when_FpuPlugin_l237_2 = 1'b1;
      end
    end
  end

  assign when_FpuPlugin_l237 = (|{_zz_when_FpuPlugin_l237_2,{_zz_when_FpuPlugin_l237_1,_zz_when_FpuPlugin_l237}});
  always @(*) begin
    FpuPlugin_accessFpuCsr = 1'b0;
    if(execute_CsrPlugin_csr_3) begin
      FpuPlugin_accessFpuCsr = 1'b1;
    end
    if(execute_CsrPlugin_csr_2) begin
      FpuPlugin_accessFpuCsr = 1'b1;
    end
    if(execute_CsrPlugin_csr_1) begin
      FpuPlugin_accessFpuCsr = 1'b1;
    end
  end

  assign when_FpuPlugin_l253 = ((FpuPlugin_accessFpuCsr && (FpuPlugin_fs == 2'b00)) && (! debugMode));
  always @(*) begin
    _zz_decode_FPU_FORKED = 1'b0;
    if(when_FpuPlugin_l350) begin
      _zz_decode_FPU_FORKED = 1'b1;
    end
  end

  assign decode_FpuPlugin_trap = (((_zz_decode_FPU_ENABLE && (FpuPlugin_fs == 2'b00)) && (! debugMode)) && (! (|{writeBack_arbitration_isValid,{memory_arbitration_isValid,execute_arbitration_isValid}})));
  assign when_FpuPlugin_l268 = (FpuPlugin_port_cmd_fire && (! _zz_decode_FPU_FORKED));
  assign when_FpuPlugin_l268_1 = (! decode_arbitration_isStuck);
  assign decode_FpuPlugin_hazard = ((FpuPlugin_pendings[5] || FpuPlugin_csrActive) || ((FpuPlugin_fs == 2'b00) && (! debugMode)));
  assign when_FpuPlugin_l272 = (! decode_LEGAL_INSTRUCTION);
  assign when_FpuPlugin_l273 = ((decode_arbitration_isValid && decode_FPU_ENABLE) && decode_FpuPlugin_hazard);
  assign FpuPlugin_port_cmd_isStall = (FpuPlugin_port_cmd_valid && (! FpuPlugin_port_cmd_ready));
  assign decode_FpuPlugin_iRoundMode = decode_INSTRUCTION[14 : 12];
  assign decode_FpuPlugin_roundMode = ((decode_INSTRUCTION[14 : 12] == 3'b111) ? FpuPlugin_rm : decode_INSTRUCTION[14 : 12]);
  always @(*) begin
    FpuPlugin_port_cmd_valid = (((decode_arbitration_isValid && decode_FPU_ENABLE) && (! decode_FpuPlugin_forked)) && (! decode_FpuPlugin_hazard));
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_valid = 1'b1;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_cmd_payload_opcode = decode_FPU_OPCODE;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        if(fpuAccess_write) begin
          FpuPlugin_port_cmd_payload_opcode = FpuOpcode_LOAD;
        end else begin
          FpuPlugin_port_cmd_payload_opcode = FpuOpcode_STORE;
        end
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign FpuPlugin_port_cmd_payload_arg = decode_FPU_ARG;
  assign FpuPlugin_port_cmd_payload_rs1 = decode_INSTRUCTION[19 : 15];
  always @(*) begin
    FpuPlugin_port_cmd_payload_rs2 = decode_INSTRUCTION[24 : 20];
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_payload_rs2 = fpuAccess_regId;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign FpuPlugin_port_cmd_payload_rs3 = decode_INSTRUCTION[31 : 27];
  always @(*) begin
    FpuPlugin_port_cmd_payload_rd = decode_INSTRUCTION[11 : 7];
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_payload_rd = fpuAccess_regId;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_cmd_payload_format = decode_FPU_FORMAT;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
        FpuPlugin_port_cmd_payload_format = _zz_FpuPlugin_port_cmd_payload_format;
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign _zz_FpuPlugin_port_cmd_payload_roundMode_1 = decode_FpuPlugin_roundMode;
  assign _zz_FpuPlugin_port_cmd_payload_roundMode = _zz_FpuPlugin_port_cmd_payload_roundMode_1;
  assign FpuPlugin_port_cmd_payload_roundMode = _zz_FpuPlugin_port_cmd_payload_roundMode;
  assign writeBack_FpuPlugin_isRsp = (writeBack_FPU_FORKED && writeBack_FPU_RSP);
  assign writeBack_FpuPlugin_isCommit = (writeBack_FPU_FORKED && writeBack_FPU_COMMIT);
  always @(*) begin
    writeBack_FpuPlugin_storeFormated = FpuPlugin_port_rsp_payload_value;
    if(when_FpuPlugin_l306) begin
      writeBack_FpuPlugin_storeFormated[63 : 32] = FpuPlugin_port_rsp_payload_value[31 : 0];
    end
  end

  assign when_FpuPlugin_l306 = (! writeBack_INSTRUCTION[12]);
  always @(*) begin
    FpuPlugin_port_rsp_ready = 1'b0;
    if(writeBack_FpuPlugin_isRsp) begin
      if(!when_FpuPlugin_l323) begin
        if(when_FpuPlugin_l325) begin
          FpuPlugin_port_rsp_ready = 1'b1;
        end
      end
    end
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
        FpuPlugin_port_rsp_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign DBusBypass0_value = writeBack_FpuPlugin_storeFormated;
  assign when_FpuPlugin_l315 = ((! writeBack_arbitration_isStuck) && (! writeBack_arbitration_removeIt));
  assign when_FpuPlugin_l318 = (FpuPlugin_port_rsp_payload_NV || FpuPlugin_port_rsp_payload_NX);
  assign when_FpuPlugin_l323 = (! FpuPlugin_port_rsp_valid);
  assign when_FpuPlugin_l325 = (! writeBack_arbitration_haltItself);
  assign writeBack_FpuPlugin_commit_valid = (writeBack_FpuPlugin_isCommit && (! writeBack_arbitration_isStuck));
  always @(*) begin
    writeBack_FpuPlugin_commit_payload_value[31 : 0] = (writeBack_FPU_COMMIT_LOAD ? _zz_writeBack_FpuPlugin_commit_payload_value[31 : 0] : writeBack_RS1);
    writeBack_FpuPlugin_commit_payload_value[63 : 32] = _zz_writeBack_FpuPlugin_commit_payload_value[63 : 32];
  end

  assign writeBack_FpuPlugin_commit_payload_write = (writeBack_arbitration_isValid && (! writeBack_arbitration_removeIt));
  assign writeBack_FpuPlugin_commit_payload_opcode = writeBack_FPU_OPCODE;
  assign writeBack_FpuPlugin_commit_payload_rd = writeBack_INSTRUCTION[11 : 7];
  assign when_FpuPlugin_l339 = (writeBack_FpuPlugin_isCommit && (! writeBack_FpuPlugin_commit_ready));
  assign writeBack_FpuPlugin_commit_ready = writeBack_FpuPlugin_commit_rValidN;
  assign writeBack_FpuPlugin_commit_s2mPipe_valid = (writeBack_FpuPlugin_commit_valid || (! writeBack_FpuPlugin_commit_rValidN));
  assign _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_opcode : writeBack_FpuPlugin_commit_rData_opcode);
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_opcode = _zz_writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_rd = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_rd : writeBack_FpuPlugin_commit_rData_rd);
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_write = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_write : writeBack_FpuPlugin_commit_rData_write);
  assign writeBack_FpuPlugin_commit_s2mPipe_payload_value = (writeBack_FpuPlugin_commit_rValidN ? writeBack_FpuPlugin_commit_payload_value : writeBack_FpuPlugin_commit_rData_value);
  always @(*) begin
    FpuPlugin_port_commit_valid = writeBack_FpuPlugin_commit_s2mPipe_valid;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_valid = 1'b1;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign writeBack_FpuPlugin_commit_s2mPipe_ready = FpuPlugin_port_commit_ready;
  always @(*) begin
    FpuPlugin_port_commit_payload_opcode = writeBack_FpuPlugin_commit_s2mPipe_payload_opcode;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_opcode = FpuOpcode_LOAD;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_commit_payload_rd = writeBack_FpuPlugin_commit_s2mPipe_payload_rd;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_rd = fpuAccess_regId;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_commit_payload_write = writeBack_FpuPlugin_commit_s2mPipe_payload_write;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_write = 1'b1;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    FpuPlugin_port_commit_payload_value = writeBack_FpuPlugin_commit_s2mPipe_payload_value;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
        FpuPlugin_port_commit_payload_value = fpuAccess_writeData;
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign FpuPlugin_wantExit = 1'b0;
  always @(*) begin
    FpuPlugin_wantStart = 1'b0;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
        FpuPlugin_wantStart = 1'b1;
      end
    endcase
  end

  assign FpuPlugin_wantKill = 1'b0;
  assign when_FpuPlugin_l350 = (! (FpuPlugin_stateReg == FpuPlugin_enumDef_IDLE));
  always @(*) begin
    fpuAccess_done = 1'b0;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
      end
      FpuPlugin_enumDef_RSP_1 : begin
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
        fpuAccess_done = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fpuAccess_readDataValid = 1'b0;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
        fpuAccess_readDataValid = 1'b1;
      end
      FpuPlugin_enumDef_RSP_1 : begin
        fpuAccess_readDataValid = 1'b1;
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fpuAccess_readDataChunk = 1'bx;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
        fpuAccess_readDataChunk = 1'b0;
      end
      FpuPlugin_enumDef_RSP_1 : begin
        fpuAccess_readDataChunk = 1'b1;
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fpuAccess_readData = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
      end
      FpuPlugin_enumDef_CMD : begin
      end
      FpuPlugin_enumDef_RSP : begin
      end
      FpuPlugin_enumDef_RSP_0 : begin
        fpuAccess_readData = FpuPlugin_port_rsp_payload_value[31 : 0];
      end
      FpuPlugin_enumDef_RSP_1 : begin
        fpuAccess_readData = FpuPlugin_port_rsp_payload_value[63 : 32];
      end
      FpuPlugin_enumDef_COMMIT : begin
      end
      FpuPlugin_enumDef_DONE : begin
      end
      default : begin
      end
    endcase
  end

  assign when_CfuPlugin_l192 = (! execute_LEGAL_INSTRUCTION);
  assign execute_CfuPlugin_hazard = (|{(writeBack_arbitration_isValid && writeBack_HAS_SIDE_EFFECT),(memory_arbitration_isValid && memory_HAS_SIDE_EFFECT)});
  assign execute_CfuPlugin_scheduleWish = (execute_arbitration_isValid && execute_CfuPlugin_CFU_ENABLE);
  assign execute_CfuPlugin_schedule = (execute_CfuPlugin_scheduleWish && (! execute_CfuPlugin_hazard));
  assign when_CfuPlugin_l196 = (execute_CfuPlugin_scheduleWish && execute_CfuPlugin_hazard);
  assign CfuPlugin_bus_cmd_fire = (CfuPlugin_bus_cmd_valid && CfuPlugin_bus_cmd_ready);
  assign when_CfuPlugin_l199 = (! execute_arbitration_isStuck);
  assign CfuPlugin_bus_cmd_valid = ((execute_CfuPlugin_schedule || execute_CfuPlugin_hold) && (! execute_CfuPlugin_fired));
  assign when_CfuPlugin_l203 = (CfuPlugin_bus_cmd_valid && (! CfuPlugin_bus_cmd_ready));
  assign execute_CfuPlugin_functionsIds_0 = {execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[14 : 12]};
  assign CfuPlugin_bus_cmd_payload_function_id = execute_CfuPlugin_functionsIds_0;
  assign CfuPlugin_bus_cmd_payload_inputs_0 = execute_RS1;
  assign _zz_CfuPlugin_bus_cmd_payload_inputs_1 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[23] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[22] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[21] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[20] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[19] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[18] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[17] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[16] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[15] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[14] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[13] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[12] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[11] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[10] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[9] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[8] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[7] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[6] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[5] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[4] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[3] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[2] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[1] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
    _zz_CfuPlugin_bus_cmd_payload_inputs_1_1[0] = _zz_CfuPlugin_bus_cmd_payload_inputs_1;
  end

  always @(*) begin
    case(execute_CfuPlugin_CFU_INPUT_2_KIND)
      Input2Kind_RS : begin
        _zz_CfuPlugin_bus_cmd_payload_inputs_1_2 = execute_RS2;
      end
      default : begin
        _zz_CfuPlugin_bus_cmd_payload_inputs_1_2 = {_zz_CfuPlugin_bus_cmd_payload_inputs_1_1,execute_INSTRUCTION[31 : 24]};
      end
    endcase
  end

  assign CfuPlugin_bus_cmd_payload_inputs_1 = _zz_CfuPlugin_bus_cmd_payload_inputs_1_2;
  assign CfuPlugin_bus_rsp_ready = CfuPlugin_bus_rsp_rValidN;
  assign writeBack_CfuPlugin_rsp_valid = (CfuPlugin_bus_rsp_valid || (! CfuPlugin_bus_rsp_rValidN));
  assign writeBack_CfuPlugin_rsp_payload_outputs_0 = (CfuPlugin_bus_rsp_rValidN ? CfuPlugin_bus_rsp_payload_outputs_0 : CfuPlugin_bus_rsp_rData_outputs_0);
  always @(*) begin
    writeBack_CfuPlugin_rsp_ready = 1'b0;
    if(writeBack_CfuPlugin_CFU_IN_FLIGHT) begin
      writeBack_CfuPlugin_rsp_ready = (! writeBack_arbitration_isStuckByOthers);
    end
  end

  assign when_CfuPlugin_l239 = (! writeBack_CfuPlugin_rsp_valid);
  always @(*) begin
    _zz_decode_RS2_3[0] = memory_SHIFT_RIGHT[31];
    _zz_decode_RS2_3[1] = memory_SHIFT_RIGHT[30];
    _zz_decode_RS2_3[2] = memory_SHIFT_RIGHT[29];
    _zz_decode_RS2_3[3] = memory_SHIFT_RIGHT[28];
    _zz_decode_RS2_3[4] = memory_SHIFT_RIGHT[27];
    _zz_decode_RS2_3[5] = memory_SHIFT_RIGHT[26];
    _zz_decode_RS2_3[6] = memory_SHIFT_RIGHT[25];
    _zz_decode_RS2_3[7] = memory_SHIFT_RIGHT[24];
    _zz_decode_RS2_3[8] = memory_SHIFT_RIGHT[23];
    _zz_decode_RS2_3[9] = memory_SHIFT_RIGHT[22];
    _zz_decode_RS2_3[10] = memory_SHIFT_RIGHT[21];
    _zz_decode_RS2_3[11] = memory_SHIFT_RIGHT[20];
    _zz_decode_RS2_3[12] = memory_SHIFT_RIGHT[19];
    _zz_decode_RS2_3[13] = memory_SHIFT_RIGHT[18];
    _zz_decode_RS2_3[14] = memory_SHIFT_RIGHT[17];
    _zz_decode_RS2_3[15] = memory_SHIFT_RIGHT[16];
    _zz_decode_RS2_3[16] = memory_SHIFT_RIGHT[15];
    _zz_decode_RS2_3[17] = memory_SHIFT_RIGHT[14];
    _zz_decode_RS2_3[18] = memory_SHIFT_RIGHT[13];
    _zz_decode_RS2_3[19] = memory_SHIFT_RIGHT[12];
    _zz_decode_RS2_3[20] = memory_SHIFT_RIGHT[11];
    _zz_decode_RS2_3[21] = memory_SHIFT_RIGHT[10];
    _zz_decode_RS2_3[22] = memory_SHIFT_RIGHT[9];
    _zz_decode_RS2_3[23] = memory_SHIFT_RIGHT[8];
    _zz_decode_RS2_3[24] = memory_SHIFT_RIGHT[7];
    _zz_decode_RS2_3[25] = memory_SHIFT_RIGHT[6];
    _zz_decode_RS2_3[26] = memory_SHIFT_RIGHT[5];
    _zz_decode_RS2_3[27] = memory_SHIFT_RIGHT[4];
    _zz_decode_RS2_3[28] = memory_SHIFT_RIGHT[3];
    _zz_decode_RS2_3[29] = memory_SHIFT_RIGHT[2];
    _zz_decode_RS2_3[30] = memory_SHIFT_RIGHT[1];
    _zz_decode_RS2_3[31] = memory_SHIFT_RIGHT[0];
  end

  assign when_Pipeline_l124 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_1 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_2 = ((! writeBack_arbitration_isStuck) && (! CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack));
  assign when_Pipeline_l124_3 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_4 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_5 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_6 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_7 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_8 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_9 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_10 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_11 = (! execute_arbitration_isStuck);
  assign _zz_decode_SRC1_CTRL = _zz_decode_SRC1_CTRL_1;
  assign when_Pipeline_l124_12 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_13 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_14 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_15 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_CTRL_1 = decode_ALU_CTRL;
  assign _zz_decode_ALU_CTRL = _zz_decode_ALU_CTRL_1;
  assign when_Pipeline_l124_16 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_CTRL = decode_to_execute_ALU_CTRL;
  assign _zz_decode_SRC2_CTRL = _zz_decode_SRC2_CTRL_1;
  assign when_Pipeline_l124_17 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_18 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_19 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_20 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_21 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_22 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_23 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_24 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_25 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_26 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_27 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_28 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_29 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_30 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_31 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_32 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_33 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_34 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_35 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_36 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_37 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_38 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_39 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ENV_CTRL_1 = decode_ENV_CTRL;
  assign _zz_execute_to_memory_ENV_CTRL_1 = execute_ENV_CTRL;
  assign _zz_memory_to_writeBack_ENV_CTRL_1 = memory_ENV_CTRL;
  assign _zz_decode_ENV_CTRL = _zz_decode_ENV_CTRL_1;
  assign when_Pipeline_l124_40 = (! execute_arbitration_isStuck);
  assign _zz_execute_ENV_CTRL = decode_to_execute_ENV_CTRL;
  assign when_Pipeline_l124_41 = (! memory_arbitration_isStuck);
  assign _zz_memory_ENV_CTRL = execute_to_memory_ENV_CTRL;
  assign when_Pipeline_l124_42 = (! writeBack_arbitration_isStuck);
  assign _zz_writeBack_ENV_CTRL = memory_to_writeBack_ENV_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL_1 = decode_BRANCH_CTRL;
  assign _zz_decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL_1;
  assign when_Pipeline_l124_43 = (! execute_arbitration_isStuck);
  assign _zz_execute_BRANCH_CTRL = decode_to_execute_BRANCH_CTRL;
  assign when_Pipeline_l124_44 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_45 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_46 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_47 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_48 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_49 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_50 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_51 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_52 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_53 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_54 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_55 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_56 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_57 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_FPU_OPCODE_1 = decode_FPU_OPCODE;
  assign _zz_execute_to_memory_FPU_OPCODE_1 = execute_FPU_OPCODE;
  assign _zz_memory_to_writeBack_FPU_OPCODE_1 = memory_FPU_OPCODE;
  assign _zz_decode_FPU_OPCODE = _zz_decode_FPU_OPCODE_1;
  assign when_Pipeline_l124_58 = (! execute_arbitration_isStuck);
  assign _zz_execute_FPU_OPCODE = decode_to_execute_FPU_OPCODE;
  assign when_Pipeline_l124_59 = (! memory_arbitration_isStuck);
  assign _zz_memory_FPU_OPCODE = execute_to_memory_FPU_OPCODE;
  assign when_Pipeline_l124_60 = (! writeBack_arbitration_isStuck);
  assign _zz_writeBack_FPU_OPCODE = memory_to_writeBack_FPU_OPCODE;
  assign _zz_decode_FPU_FORMAT = _zz_decode_FPU_FORMAT_1;
  assign when_Pipeline_l124_61 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND_1 = decode_CfuPlugin_CFU_INPUT_2_KIND;
  assign _zz_decode_CfuPlugin_CFU_INPUT_2_KIND = _zz_decode_CfuPlugin_CFU_INPUT_2_KIND_1;
  assign when_Pipeline_l124_62 = (! execute_arbitration_isStuck);
  assign _zz_execute_CfuPlugin_CFU_INPUT_2_KIND = decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL_1 = decode_ALU_BITWISE_CTRL;
  assign _zz_decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL_1;
  assign when_Pipeline_l124_63 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_BITWISE_CTRL = decode_to_execute_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL_1 = decode_SHIFT_CTRL;
  assign _zz_execute_to_memory_SHIFT_CTRL_1 = execute_SHIFT_CTRL;
  assign _zz_decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL_1;
  assign when_Pipeline_l124_64 = (! execute_arbitration_isStuck);
  assign _zz_execute_SHIFT_CTRL = decode_to_execute_SHIFT_CTRL;
  assign when_Pipeline_l124_65 = (! memory_arbitration_isStuck);
  assign _zz_memory_SHIFT_CTRL = execute_to_memory_SHIFT_CTRL;
  assign when_Pipeline_l124_66 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_67 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_68 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_69 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_70 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_71 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_72 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_73 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_74 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_75 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_76 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_77 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_78 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_79 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_80 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_81 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_82 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_83 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_84 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_85 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_86 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_87 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_88 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_89 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_90 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_91 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_92 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_93 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_94 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_95 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_96 = (! writeBack_arbitration_isStuck);
  assign decode_arbitration_isFlushed = ((|{writeBack_arbitration_flushNext,{memory_arbitration_flushNext,execute_arbitration_flushNext}}) || (|{writeBack_arbitration_flushIt,{memory_arbitration_flushIt,{execute_arbitration_flushIt,decode_arbitration_flushIt}}}));
  assign execute_arbitration_isFlushed = ((|{writeBack_arbitration_flushNext,memory_arbitration_flushNext}) || (|{writeBack_arbitration_flushIt,{memory_arbitration_flushIt,execute_arbitration_flushIt}}));
  assign memory_arbitration_isFlushed = ((|writeBack_arbitration_flushNext) || (|{writeBack_arbitration_flushIt,memory_arbitration_flushIt}));
  assign writeBack_arbitration_isFlushed = (1'b0 || (|writeBack_arbitration_flushIt));
  assign decode_arbitration_isStuckByOthers = (decode_arbitration_haltByOther || (((1'b0 || execute_arbitration_isStuck) || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign decode_arbitration_isStuck = (decode_arbitration_haltItself || decode_arbitration_isStuckByOthers);
  assign decode_arbitration_isMoving = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign decode_arbitration_isFiring = ((decode_arbitration_isValid && (! decode_arbitration_isStuck)) && (! decode_arbitration_removeIt));
  assign execute_arbitration_isStuckByOthers = (execute_arbitration_haltByOther || ((1'b0 || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign execute_arbitration_isStuck = (execute_arbitration_haltItself || execute_arbitration_isStuckByOthers);
  assign execute_arbitration_isMoving = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign execute_arbitration_isFiring = ((execute_arbitration_isValid && (! execute_arbitration_isStuck)) && (! execute_arbitration_removeIt));
  assign memory_arbitration_isStuckByOthers = (memory_arbitration_haltByOther || (1'b0 || writeBack_arbitration_isStuck));
  assign memory_arbitration_isStuck = (memory_arbitration_haltItself || memory_arbitration_isStuckByOthers);
  assign memory_arbitration_isMoving = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  assign memory_arbitration_isFiring = ((memory_arbitration_isValid && (! memory_arbitration_isStuck)) && (! memory_arbitration_removeIt));
  assign writeBack_arbitration_isStuckByOthers = (writeBack_arbitration_haltByOther || 1'b0);
  assign writeBack_arbitration_isStuck = (writeBack_arbitration_haltItself || writeBack_arbitration_isStuckByOthers);
  assign writeBack_arbitration_isMoving = ((! writeBack_arbitration_isStuck) && (! writeBack_arbitration_removeIt));
  assign writeBack_arbitration_isFiring = ((writeBack_arbitration_isValid && (! writeBack_arbitration_isStuck)) && (! writeBack_arbitration_removeIt));
  assign when_Pipeline_l151 = ((! execute_arbitration_isStuck) || execute_arbitration_removeIt);
  assign when_Pipeline_l154 = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign when_Pipeline_l151_1 = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  assign when_Pipeline_l154_1 = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign when_Pipeline_l151_2 = ((! writeBack_arbitration_isStuck) || writeBack_arbitration_removeIt);
  assign when_Pipeline_l154_2 = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  always @(*) begin
    CsrPlugin_injectionPort_ready = 1'b0;
    case(IBusCachedPlugin_injector_port_state)
      3'b100 : begin
        CsrPlugin_injectionPort_ready = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign when_Fetcher_l373 = (IBusCachedPlugin_injector_port_state != 3'b000);
  assign when_Fetcher_l391 = (! decode_arbitration_isStuck);
  assign when_Fetcher_l411 = (IBusCachedPlugin_injector_port_state != 3'b000);
  assign when_CsrPlugin_l1813 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_2 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_3 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_4 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_5 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_6 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_7 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_8 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_9 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_10 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_11 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_12 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_13 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_14 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_15 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_16 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_17 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_18 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1813_19 = (! execute_arbitration_isStuck);
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit = 32'h0;
    if(execute_CsrPlugin_csr_1972) begin
      _zz_CsrPlugin_csrMapping_readDataInit[31 : 0] = CsrPlugin_dataCsrw_value_0;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_1 = 32'h0;
    if(execute_CsrPlugin_csr_1969) begin
      _zz_CsrPlugin_csrMapping_readDataInit_1[31 : 0] = CsrPlugin_dpc;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_2 = 32'h0;
    if(execute_CsrPlugin_csr_1968) begin
      _zz_CsrPlugin_csrMapping_readDataInit_2[3 : 3] = CsrPlugin_dcsr_nmip;
      _zz_CsrPlugin_csrMapping_readDataInit_2[8 : 6] = CsrPlugin_dcsr_cause;
      _zz_CsrPlugin_csrMapping_readDataInit_2[31 : 28] = CsrPlugin_dcsr_xdebugver;
      _zz_CsrPlugin_csrMapping_readDataInit_2[4 : 4] = CsrPlugin_dcsr_mprven;
      _zz_CsrPlugin_csrMapping_readDataInit_2[1 : 0] = CsrPlugin_dcsr_prv;
      _zz_CsrPlugin_csrMapping_readDataInit_2[2 : 2] = CsrPlugin_dcsr_step;
      _zz_CsrPlugin_csrMapping_readDataInit_2[9 : 9] = CsrPlugin_dcsr_stoptime;
      _zz_CsrPlugin_csrMapping_readDataInit_2[10 : 10] = CsrPlugin_dcsr_stopcount;
      _zz_CsrPlugin_csrMapping_readDataInit_2[11 : 11] = CsrPlugin_dcsr_stepie;
      _zz_CsrPlugin_csrMapping_readDataInit_2[15 : 15] = CsrPlugin_dcsr_ebreakm;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_3 = 32'h0;
    if(execute_CsrPlugin_csr_769) begin
      _zz_CsrPlugin_csrMapping_readDataInit_3[31 : 30] = CsrPlugin_misa_base;
      _zz_CsrPlugin_csrMapping_readDataInit_3[25 : 0] = CsrPlugin_misa_extensions;
    end
  end

  assign switch_CsrPlugin_l1167 = CsrPlugin_csrMapping_writeDataSignal[12 : 11];
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_4 = 32'h0;
    if(execute_CsrPlugin_csr_768) begin
      _zz_CsrPlugin_csrMapping_readDataInit_4[7 : 7] = CsrPlugin_mstatus_MPIE;
      _zz_CsrPlugin_csrMapping_readDataInit_4[3 : 3] = CsrPlugin_mstatus_MIE;
      _zz_CsrPlugin_csrMapping_readDataInit_4[12 : 11] = CsrPlugin_mstatus_MPP;
      _zz_CsrPlugin_csrMapping_readDataInit_4[14 : 13] = FpuPlugin_fs;
      _zz_CsrPlugin_csrMapping_readDataInit_4[31 : 31] = FpuPlugin_sd;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_5 = 32'h0;
    if(execute_CsrPlugin_csr_836) begin
      _zz_CsrPlugin_csrMapping_readDataInit_5[11 : 11] = CsrPlugin_mip_MEIP;
      _zz_CsrPlugin_csrMapping_readDataInit_5[7 : 7] = CsrPlugin_mip_MTIP;
      _zz_CsrPlugin_csrMapping_readDataInit_5[3 : 3] = CsrPlugin_mip_MSIP;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_6 = 32'h0;
    if(execute_CsrPlugin_csr_772) begin
      _zz_CsrPlugin_csrMapping_readDataInit_6[11 : 11] = CsrPlugin_mie_MEIE;
      _zz_CsrPlugin_csrMapping_readDataInit_6[7 : 7] = CsrPlugin_mie_MTIE;
      _zz_CsrPlugin_csrMapping_readDataInit_6[3 : 3] = CsrPlugin_mie_MSIE;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_7 = 32'h0;
    if(execute_CsrPlugin_csr_773) begin
      _zz_CsrPlugin_csrMapping_readDataInit_7[31 : 2] = CsrPlugin_mtvec_base;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_8 = 32'h0;
    if(execute_CsrPlugin_csr_833) begin
      _zz_CsrPlugin_csrMapping_readDataInit_8[31 : 0] = CsrPlugin_mepc;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_9 = 32'h0;
    if(execute_CsrPlugin_csr_832) begin
      _zz_CsrPlugin_csrMapping_readDataInit_9[31 : 0] = CsrPlugin_mscratch;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_10 = 32'h0;
    if(execute_CsrPlugin_csr_834) begin
      _zz_CsrPlugin_csrMapping_readDataInit_10[31 : 31] = CsrPlugin_mcause_interrupt;
      _zz_CsrPlugin_csrMapping_readDataInit_10[3 : 0] = CsrPlugin_mcause_exceptionCode;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_11 = 32'h0;
    if(execute_CsrPlugin_csr_835) begin
      _zz_CsrPlugin_csrMapping_readDataInit_11[31 : 0] = CsrPlugin_mtval;
    end
  end

  assign _zz_FpuPlugin_flags_NX = CsrPlugin_csrMapping_writeDataSignal[4 : 0];
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_12 = 32'h0;
    if(execute_CsrPlugin_csr_3) begin
      _zz_CsrPlugin_csrMapping_readDataInit_12[7 : 5] = FpuPlugin_rm;
      _zz_CsrPlugin_csrMapping_readDataInit_12[4 : 0] = {FpuPlugin_flags_NV,{FpuPlugin_flags_DZ,{FpuPlugin_flags_OF,{FpuPlugin_flags_UF,FpuPlugin_flags_NX}}}};
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_13 = 32'h0;
    if(execute_CsrPlugin_csr_2) begin
      _zz_CsrPlugin_csrMapping_readDataInit_13[2 : 0] = FpuPlugin_rm;
    end
  end

  assign _zz_FpuPlugin_flags_NX_1 = CsrPlugin_csrMapping_writeDataSignal[4 : 0];
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_14 = 32'h0;
    if(execute_CsrPlugin_csr_1) begin
      _zz_CsrPlugin_csrMapping_readDataInit_14[4 : 0] = {FpuPlugin_flags_NV,{FpuPlugin_flags_DZ,{FpuPlugin_flags_OF,{FpuPlugin_flags_UF,FpuPlugin_flags_NX}}}};
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_15 = 32'h0;
    if(execute_CsrPlugin_csr_256) begin
      _zz_CsrPlugin_csrMapping_readDataInit_15[14 : 13] = FpuPlugin_fs;
      _zz_CsrPlugin_csrMapping_readDataInit_15[31 : 31] = FpuPlugin_sd;
    end
  end

  assign CsrPlugin_csrMapping_readDataInit = (((((_zz_CsrPlugin_csrMapping_readDataInit | _zz_CsrPlugin_csrMapping_readDataInit_1) | (_zz_CsrPlugin_csrMapping_readDataInit_2 | _zz_CsrPlugin_csrMapping_readDataInit_16)) | ((_zz_CsrPlugin_csrMapping_readDataInit_17 | _zz_CsrPlugin_csrMapping_readDataInit_18) | (_zz_CsrPlugin_csrMapping_readDataInit_19 | _zz_CsrPlugin_csrMapping_readDataInit_3))) | (((_zz_CsrPlugin_csrMapping_readDataInit_4 | _zz_CsrPlugin_csrMapping_readDataInit_5) | (_zz_CsrPlugin_csrMapping_readDataInit_6 | _zz_CsrPlugin_csrMapping_readDataInit_7)) | ((_zz_CsrPlugin_csrMapping_readDataInit_8 | _zz_CsrPlugin_csrMapping_readDataInit_9) | (_zz_CsrPlugin_csrMapping_readDataInit_10 | _zz_CsrPlugin_csrMapping_readDataInit_11)))) | ((_zz_CsrPlugin_csrMapping_readDataInit_12 | _zz_CsrPlugin_csrMapping_readDataInit_13) | (_zz_CsrPlugin_csrMapping_readDataInit_14 | _zz_CsrPlugin_csrMapping_readDataInit_15)));
  assign when_CsrPlugin_l1846 = ((execute_arbitration_isValid && execute_IS_CSR) && (({execute_CsrPlugin_csrAddress[11 : 2],2'b00} == 12'h3a0) || ({execute_CsrPlugin_csrAddress[11 : 4],4'b0000} == 12'h3b0)));
  assign _zz_when_CsrPlugin_l1853 = (execute_CsrPlugin_csrAddress & 12'hf60);
  assign when_CsrPlugin_l1853 = (((execute_arbitration_isValid && execute_IS_CSR) && (5'h03 <= execute_CsrPlugin_csrAddress[4 : 0])) && (((_zz_when_CsrPlugin_l1853 == 12'hb00) || (((_zz_when_CsrPlugin_l1853 == 12'hc00) && (! execute_CsrPlugin_writeInstruction)) && (CsrPlugin_privilege == 2'b11))) || ((execute_CsrPlugin_csrAddress & 12'hfe0) == 12'h320)));
  always @(*) begin
    when_CsrPlugin_l1863 = CsrPlugin_csrMapping_doForceFailCsr;
    if(when_CsrPlugin_l1861) begin
      when_CsrPlugin_l1863 = 1'b1;
    end
    if(when_CsrPlugin_l1862) begin
      when_CsrPlugin_l1863 = 1'b1;
    end
  end

  assign when_CsrPlugin_l1861 = (CsrPlugin_privilege < execute_CsrPlugin_csrAddress[9 : 8]);
  assign when_CsrPlugin_l1862 = ((! debugMode) && (_zz_when_CsrPlugin_l1862 == 8'h7b));
  assign when_CsrPlugin_l1869 = ((! execute_arbitration_isValid) || (! execute_IS_CSR));
  always @(*) begin
    FpuPlugin_stateNext = FpuPlugin_stateReg;
    case(FpuPlugin_stateReg)
      FpuPlugin_enumDef_IDLE : begin
        if(fpuAccess_start) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_CMD;
        end
      end
      FpuPlugin_enumDef_CMD : begin
        if(fpuAccess_write) begin
          if(FpuPlugin_port_cmd_ready) begin
            FpuPlugin_stateNext = FpuPlugin_enumDef_COMMIT;
          end
        end else begin
          if(FpuPlugin_port_cmd_ready) begin
            FpuPlugin_stateNext = FpuPlugin_enumDef_RSP;
          end
        end
      end
      FpuPlugin_enumDef_RSP : begin
        if(FpuPlugin_port_rsp_valid) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_RSP_0;
        end
      end
      FpuPlugin_enumDef_RSP_0 : begin
        if(when_FpuPlugin_l402) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_RSP_1;
        end else begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_DONE;
        end
      end
      FpuPlugin_enumDef_RSP_1 : begin
        FpuPlugin_stateNext = FpuPlugin_enumDef_DONE;
      end
      FpuPlugin_enumDef_COMMIT : begin
        if(FpuPlugin_port_commit_ready) begin
          FpuPlugin_stateNext = FpuPlugin_enumDef_DONE;
        end
      end
      FpuPlugin_enumDef_DONE : begin
        FpuPlugin_stateNext = FpuPlugin_enumDef_IDLE;
      end
      default : begin
      end
    endcase
    if(FpuPlugin_wantStart) begin
      FpuPlugin_stateNext = FpuPlugin_enumDef_IDLE;
    end
    if(FpuPlugin_wantKill) begin
      FpuPlugin_stateNext = FpuPlugin_enumDef_BOOT;
    end
  end

  always @(*) begin
    _zz_FpuPlugin_port_cmd_payload_format = (1'bx);
    case(fpuAccess_size)
      3'b010 : begin
        _zz_FpuPlugin_port_cmd_payload_format = FpuFormat_FLOAT;
      end
      3'b011 : begin
        _zz_FpuPlugin_port_cmd_payload_format = FpuFormat_DOUBLE;
      end
      default : begin
      end
    endcase
  end

  assign when_FpuPlugin_l402 = (3'b010 < fpuAccess_size);
  assign DBusCachedPlugin_trigger_hitBefore = 1'b0;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      IBusCachedPlugin_fetchPc_pcReg <= 32'hf9000000;
      IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      IBusCachedPlugin_fetchPc_booted <= 1'b0;
      IBusCachedPlugin_fetchPc_inc <= 1'b0;
      IBusCachedPlugin_decodePc_pcReg <= 32'hf9000000;
      _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1 <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      IBusCachedPlugin_decompressor_bufferValid <= 1'b0;
      IBusCachedPlugin_decompressor_throw2BytesReg <= 1'b0;
      _zz_IBusCachedPlugin_injector_decodeInput_valid <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      IBusCachedPlugin_rspCounter <= 32'h0;
      dataCache_2_io_mem_cmd_rValidN <= 1'b1;
      dataCache_2_io_mem_cmd_s2mPipe_rValid <= 1'b0;
      dBus_rsp_valid_regNext <= 1'b0;
      DBusCachedPlugin_rspCounter <= 32'h0;
      _zz_5 <= 1'b1;
      HazardSimplePlugin_writeBackBuffer_valid <= 1'b0;
      _zz_CsrPlugin_privilege <= 2'b11;
      CsrPlugin_running <= 1'b1;
      CsrPlugin_reseting <= 1'b1;
      _zz_debugBus_haveReset <= 1'b0;
      CsrPlugin_running_aheadValue_regNext <= 1'b0;
      CsrPlugin_doHalt <= 1'b0;
      _zz_CsrPlugin_doResume <= 1'b0;
      CsrPlugin_timeout_state <= 1'b0;
      CsrPlugin_timeout_counter_value <= 3'b000;
      CsrPlugin_inject_cmd_toStream_rValid <= 1'b0;
      CsrPlugin_inject_pending <= 1'b0;
      CsrPlugin_dcsr_prv <= 2'b11;
      CsrPlugin_dcsr_step <= 1'b0;
      CsrPlugin_dcsr_cause <= 3'b000;
      CsrPlugin_dcsr_stoptime <= 1'b1;
      CsrPlugin_dcsr_stopcount <= 1'b0;
      CsrPlugin_dcsr_stepie <= 1'b0;
      CsrPlugin_dcsr_ebreakm <= 1'b0;
      CsrPlugin_dcsr_stepLogic_stateReg <= CsrPlugin_dcsr_stepLogic_enumDef_BOOT;
      stoptime <= 1'b0;
      CsrPlugin_mstatus_MIE <= 1'b0;
      CsrPlugin_mstatus_MPIE <= 1'b0;
      CsrPlugin_mstatus_MPP <= 2'b11;
      CsrPlugin_mie_MEIE <= 1'b0;
      CsrPlugin_mie_MTIE <= 1'b0;
      CsrPlugin_mie_MSIE <= 1'b0;
      CsrPlugin_counters_mcycle <= 64'h0;
      CsrPlugin_counters_minstret <= 64'h0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      CsrPlugin_interrupt_valid <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      CsrPlugin_hadException <= 1'b0;
      execute_CsrPlugin_wfiWake <= 1'b0;
      memory_MulDivIterativePlugin_div_counter_value <= 6'h0;
      FpuPlugin_pendings <= 6'h0;
      FpuPlugin_flags_NV <= 1'b0;
      FpuPlugin_flags_DZ <= 1'b0;
      FpuPlugin_flags_OF <= 1'b0;
      FpuPlugin_flags_UF <= 1'b0;
      FpuPlugin_flags_NX <= 1'b0;
      FpuPlugin_rm <= 3'b000;
      FpuPlugin_fs <= 2'b01;
      decode_FpuPlugin_forked <= 1'b0;
      writeBack_FpuPlugin_commit_rValidN <= 1'b1;
      execute_CfuPlugin_hold <= 1'b0;
      execute_CfuPlugin_fired <= 1'b0;
      CfuPlugin_bus_rsp_rValidN <= 1'b1;
      execute_arbitration_isValid <= 1'b0;
      memory_arbitration_isValid <= 1'b0;
      writeBack_arbitration_isValid <= 1'b0;
      IBusCachedPlugin_injector_port_state <= 3'b000;
      FpuPlugin_stateReg <= FpuPlugin_enumDef_BOOT;
      decode_to_execute_FPU_FORKED <= 1'b0;
      execute_to_memory_FPU_FORKED <= 1'b0;
      memory_to_writeBack_FPU_FORKED <= 1'b0;
      memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT <= 1'b0;
      execute_to_memory_CfuPlugin_CFU_IN_FLIGHT <= 1'b0;
    end else begin
      if(IBusCachedPlugin_fetchPc_correction) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_output_fire) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      end
      IBusCachedPlugin_fetchPc_booted <= 1'b1;
      if(when_Fetcher_l133) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_output_fire) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b1;
      end
      if(when_Fetcher_l133_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(when_Fetcher_l160) begin
        IBusCachedPlugin_fetchPc_pcReg <= IBusCachedPlugin_fetchPc_pc;
      end
      if(when_Fetcher_l182) begin
        IBusCachedPlugin_decodePc_pcReg <= IBusCachedPlugin_decodePc_pcPlus;
      end
      if(when_Fetcher_l194) begin
        IBusCachedPlugin_decodePc_pcReg <= IBusCachedPlugin_jump_pcLoad_payload;
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1 <= 1'b0;
      end
      if(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_input_valid_1 <= (IBusCachedPlugin_iBusRsp_stages_0_output_valid && (! 1'b0));
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      end
      if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= (IBusCachedPlugin_iBusRsp_stages_1_output_valid && (! IBusCachedPlugin_iBusRsp_flush));
      end
      if(IBusCachedPlugin_decompressor_output_fire) begin
        IBusCachedPlugin_decompressor_throw2BytesReg <= ((((! IBusCachedPlugin_decompressor_unaligned) && IBusCachedPlugin_decompressor_isInputLowRvc) && IBusCachedPlugin_decompressor_isInputHighRvc) || (IBusCachedPlugin_decompressor_bufferValid && IBusCachedPlugin_decompressor_isInputHighRvc));
      end
      if(when_Fetcher_l285) begin
        IBusCachedPlugin_decompressor_bufferValid <= 1'b0;
      end
      if(when_Fetcher_l288) begin
        if(IBusCachedPlugin_decompressor_bufferFill) begin
          IBusCachedPlugin_decompressor_bufferValid <= 1'b1;
        end
      end
      if(when_Fetcher_l293) begin
        IBusCachedPlugin_decompressor_throw2BytesReg <= 1'b0;
        IBusCachedPlugin_decompressor_bufferValid <= 1'b0;
      end
      if(decode_arbitration_removeIt) begin
        _zz_IBusCachedPlugin_injector_decodeInput_valid <= 1'b0;
      end
      if(IBusCachedPlugin_decompressor_output_ready) begin
        _zz_IBusCachedPlugin_injector_decodeInput_valid <= (IBusCachedPlugin_decompressor_output_valid && (! IBusCachedPlugin_externalFlush));
      end
      if(when_Fetcher_l331) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b1;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      end
      if(when_Fetcher_l331_1) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= IBusCachedPlugin_injector_nextPcCalc_valids_0;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(when_Fetcher_l331_2) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= IBusCachedPlugin_injector_nextPcCalc_valids_1;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(when_Fetcher_l331_3) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= IBusCachedPlugin_injector_nextPcCalc_valids_2;
      end
      if(IBusCachedPlugin_decodePc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(iBus_rsp_valid) begin
        IBusCachedPlugin_rspCounter <= (IBusCachedPlugin_rspCounter + 32'h00000001);
      end
      if(dataCache_2_io_mem_cmd_valid) begin
        dataCache_2_io_mem_cmd_rValidN <= 1'b0;
      end
      if(dataCache_2_io_mem_cmd_s2mPipe_ready) begin
        dataCache_2_io_mem_cmd_rValidN <= 1'b1;
      end
      if(dataCache_2_io_mem_cmd_s2mPipe_ready) begin
        dataCache_2_io_mem_cmd_s2mPipe_rValid <= dataCache_2_io_mem_cmd_s2mPipe_valid;
      end
      dBus_rsp_valid_regNext <= dBus_rsp_valid;
      if(dBus_rsp_valid) begin
        DBusCachedPlugin_rspCounter <= (DBusCachedPlugin_rspCounter + 32'h00000001);
      end
      _zz_5 <= 1'b0;
      HazardSimplePlugin_writeBackBuffer_valid <= HazardSimplePlugin_writeBackWrites_valid;
      CsrPlugin_reseting <= 1'b0;
      if(CsrPlugin_reseting) begin
        _zz_debugBus_haveReset <= 1'b1;
      end
      if(debugBus_ackReset) begin
        _zz_debugBus_haveReset <= 1'b0;
      end
      CsrPlugin_running_aheadValue_regNext <= CsrPlugin_running_aheadValue;
      if(when_CsrPlugin_l747) begin
        CsrPlugin_doHalt <= 1'b1;
      end
      if(CsrPlugin_enterHalt) begin
        CsrPlugin_doHalt <= 1'b0;
      end
      if(debugBus_resume_cmd_valid) begin
        _zz_CsrPlugin_doResume <= 1'b1;
      end
      if(debugBus_resume_rsp_valid) begin
        _zz_CsrPlugin_doResume <= 1'b0;
      end
      CsrPlugin_timeout_counter_value <= CsrPlugin_timeout_counter_valueNext;
      if(CsrPlugin_timeout_counter_willOverflow) begin
        CsrPlugin_timeout_state <= 1'b1;
      end
      if(when_CsrPlugin_l753) begin
        CsrPlugin_timeout_state <= 1'b0;
      end
      if(CsrPlugin_inject_cmd_toStream_ready) begin
        CsrPlugin_inject_cmd_toStream_rValid <= CsrPlugin_inject_cmd_toStream_valid;
      end
      if(when_CsrPlugin_l804) begin
        CsrPlugin_inject_pending <= 1'b1;
      end
      if(when_CsrPlugin_l804_1) begin
        CsrPlugin_inject_pending <= 1'b0;
      end
      if(CsrPlugin_inject_cmd_valid) begin
        CsrPlugin_timeout_state <= 1'b0;
      end
      CsrPlugin_dcsr_stepLogic_stateReg <= CsrPlugin_dcsr_stepLogic_stateNext;
      case(CsrPlugin_dcsr_stepLogic_stateReg)
        CsrPlugin_dcsr_stepLogic_enumDef_IDLE : begin
        end
        CsrPlugin_dcsr_stepLogic_enumDef_SINGLE : begin
          CsrPlugin_timeout_state <= 1'b0;
          if(when_CsrPlugin_l836) begin
            CsrPlugin_doHalt <= 1'b1;
          end
        end
        CsrPlugin_dcsr_stepLogic_enumDef_WAIT_1 : begin
          if(!when_CsrPlugin_l848) begin
            if(writeBack_arbitration_isFiring) begin
              CsrPlugin_doHalt <= 1'b1;
            end
          end
        end
        default : begin
        end
      endcase
      stoptime <= (debugMode && CsrPlugin_dcsr_stoptime);
      CsrPlugin_counters_mcycle <= (CsrPlugin_counters_mcycle + _zz_CsrPlugin_counters_mcycle);
      if(writeBack_arbitration_isFiring) begin
        CsrPlugin_counters_minstret <= (CsrPlugin_counters_minstret + _zz_CsrPlugin_counters_minstret);
      end
      if(when_CsrPlugin_l1403) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
      end
      if(when_CsrPlugin_l1403_1) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= (CsrPlugin_exceptionPortCtrl_exceptionValids_decode && (! decode_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
      end
      if(when_CsrPlugin_l1403_2) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= (CsrPlugin_exceptionPortCtrl_exceptionValids_execute && (! execute_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
      end
      if(when_CsrPlugin_l1403_3) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= (CsrPlugin_exceptionPortCtrl_exceptionValids_memory && (! memory_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      end
      CsrPlugin_interrupt_valid <= 1'b0;
      if(when_CsrPlugin_l1440) begin
        if(when_CsrPlugin_l1446) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l1446_1) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l1446_2) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
      end
      if(when_CsrPlugin_l1459) begin
        CsrPlugin_interrupt_valid <= 1'b0;
      end
      if(CsrPlugin_doHalt) begin
        CsrPlugin_interrupt_valid <= 1'b1;
      end
      if(CsrPlugin_pipelineLiberator_active) begin
        if(when_CsrPlugin_l1479) begin
          CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b1;
        end
        if(when_CsrPlugin_l1479_1) begin
          CsrPlugin_pipelineLiberator_pcValids_1 <= CsrPlugin_pipelineLiberator_pcValids_0;
        end
        if(when_CsrPlugin_l1479_2) begin
          CsrPlugin_pipelineLiberator_pcValids_2 <= CsrPlugin_pipelineLiberator_pcValids_1;
        end
      end
      if(when_CsrPlugin_l1484) begin
        CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      end
      if(CsrPlugin_interruptJump) begin
        CsrPlugin_interrupt_valid <= 1'b0;
      end
      CsrPlugin_hadException <= CsrPlugin_exception;
      if(when_CsrPlugin_l1534) begin
        if(when_CsrPlugin_l1542) begin
          _zz_CsrPlugin_privilege <= CsrPlugin_targetPrivilege;
          case(CsrPlugin_targetPrivilege)
            2'b11 : begin
              CsrPlugin_mstatus_MIE <= 1'b0;
              CsrPlugin_mstatus_MPIE <= CsrPlugin_mstatus_MIE;
              CsrPlugin_mstatus_MPP <= CsrPlugin_privilege;
            end
            default : begin
            end
          endcase
        end else begin
          if(when_CsrPlugin_l1572) begin
            CsrPlugin_dcsr_cause <= 3'b011;
            if(CsrPlugin_dcsr_step) begin
              CsrPlugin_dcsr_cause <= 3'b100;
            end
            if(CsrPlugin_trapCauseEbreakDebug) begin
              CsrPlugin_dcsr_cause <= 3'b001;
            end
            CsrPlugin_dcsr_prv <= CsrPlugin_privilege;
          end
          _zz_CsrPlugin_privilege <= 2'b11;
        end
      end
      if(when_CsrPlugin_l1600) begin
        case(switch_CsrPlugin_l1604)
          2'b11 : begin
            CsrPlugin_mstatus_MPP <= 2'b00;
            CsrPlugin_mstatus_MIE <= CsrPlugin_mstatus_MPIE;
            CsrPlugin_mstatus_MPIE <= 1'b1;
            _zz_CsrPlugin_privilege <= CsrPlugin_mstatus_MPP;
          end
          default : begin
          end
        endcase
      end
      if(CsrPlugin_doResume) begin
        _zz_CsrPlugin_privilege <= CsrPlugin_dcsr_prv;
      end
      execute_CsrPlugin_wfiWake <= ((|{_zz_when_CsrPlugin_l1446_2,{_zz_when_CsrPlugin_l1446_1,_zz_when_CsrPlugin_l1446}}) || CsrPlugin_thirdPartyWake);
      memory_MulDivIterativePlugin_div_counter_value <= memory_MulDivIterativePlugin_div_counter_valueNext;
      FpuPlugin_pendings <= (_zz_FpuPlugin_pendings - _zz_FpuPlugin_pendings_6);
      if(when_FpuPlugin_l215) begin
        FpuPlugin_flags_NV <= 1'b1;
      end
      if(when_FpuPlugin_l216) begin
        FpuPlugin_flags_DZ <= 1'b1;
      end
      if(when_FpuPlugin_l217) begin
        FpuPlugin_flags_OF <= 1'b1;
      end
      if(when_FpuPlugin_l218) begin
        FpuPlugin_flags_UF <= 1'b1;
      end
      if(when_FpuPlugin_l219) begin
        FpuPlugin_flags_NX <= 1'b1;
      end
      if(when_FpuPlugin_l234) begin
        FpuPlugin_fs <= 2'b11;
      end
      if(when_FpuPlugin_l237) begin
        FpuPlugin_fs <= 2'b11;
      end
      if(when_FpuPlugin_l268) begin
        decode_FpuPlugin_forked <= 1'b1;
      end
      if(when_FpuPlugin_l268_1) begin
        decode_FpuPlugin_forked <= 1'b0;
      end
      if(writeBack_FpuPlugin_isRsp) begin
        if(writeBack_arbitration_isValid) begin
          if(when_FpuPlugin_l315) begin
            if(FpuPlugin_port_rsp_payload_NV) begin
              FpuPlugin_flags_NV <= 1'b1;
            end
            if(FpuPlugin_port_rsp_payload_NX) begin
              FpuPlugin_flags_NX <= 1'b1;
            end
            if(when_FpuPlugin_l318) begin
              FpuPlugin_fs <= 2'b11;
            end
          end
        end
      end
      if(writeBack_FpuPlugin_commit_valid) begin
        writeBack_FpuPlugin_commit_rValidN <= 1'b0;
      end
      if(writeBack_FpuPlugin_commit_s2mPipe_ready) begin
        writeBack_FpuPlugin_commit_rValidN <= 1'b1;
      end
      if(execute_CfuPlugin_schedule) begin
        execute_CfuPlugin_hold <= 1'b1;
      end
      if(CfuPlugin_bus_cmd_ready) begin
        execute_CfuPlugin_hold <= 1'b0;
      end
      if(CfuPlugin_bus_cmd_fire) begin
        execute_CfuPlugin_fired <= 1'b1;
      end
      if(when_CfuPlugin_l199) begin
        execute_CfuPlugin_fired <= 1'b0;
      end
      if(CfuPlugin_bus_rsp_valid) begin
        CfuPlugin_bus_rsp_rValidN <= 1'b0;
      end
      if(writeBack_CfuPlugin_rsp_ready) begin
        CfuPlugin_bus_rsp_rValidN <= 1'b1;
      end
      if(when_Pipeline_l124_75) begin
        decode_to_execute_FPU_FORKED <= _zz_decode_to_execute_FPU_FORKED;
      end
      if(when_Pipeline_l124_76) begin
        execute_to_memory_FPU_FORKED <= _zz_execute_to_memory_FPU_FORKED;
      end
      if(when_Pipeline_l124_77) begin
        memory_to_writeBack_FPU_FORKED <= _zz_memory_to_writeBack_FPU_FORKED;
      end
      if(when_Pipeline_l124_91) begin
        execute_to_memory_CfuPlugin_CFU_IN_FLIGHT <= _zz_execute_to_memory_CfuPlugin_CFU_IN_FLIGHT;
      end
      if(when_Pipeline_l124_92) begin
        memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT <= _zz_memory_to_writeBack_CfuPlugin_CFU_IN_FLIGHT;
      end
      if(when_Pipeline_l151) begin
        execute_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154) begin
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end
      if(when_Pipeline_l151_1) begin
        memory_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_1) begin
        memory_arbitration_isValid <= execute_arbitration_isValid;
      end
      if(when_Pipeline_l151_2) begin
        writeBack_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_2) begin
        writeBack_arbitration_isValid <= memory_arbitration_isValid;
      end
      case(IBusCachedPlugin_injector_port_state)
        3'b000 : begin
          if(CsrPlugin_injectionPort_valid) begin
            IBusCachedPlugin_injector_port_state <= 3'b001;
          end
        end
        3'b001 : begin
          IBusCachedPlugin_injector_port_state <= 3'b010;
        end
        3'b010 : begin
          IBusCachedPlugin_injector_port_state <= 3'b011;
        end
        3'b011 : begin
          if(when_Fetcher_l391) begin
            IBusCachedPlugin_injector_port_state <= 3'b100;
          end
        end
        3'b100 : begin
          IBusCachedPlugin_injector_port_state <= 3'b000;
        end
        default : begin
        end
      endcase
      if(execute_CsrPlugin_csr_1968) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_dcsr_prv <= CsrPlugin_csrMapping_writeDataSignal[1 : 0];
          CsrPlugin_dcsr_step <= CsrPlugin_csrMapping_writeDataSignal[2];
          CsrPlugin_dcsr_stoptime <= CsrPlugin_csrMapping_writeDataSignal[9];
          CsrPlugin_dcsr_stopcount <= CsrPlugin_csrMapping_writeDataSignal[10];
          CsrPlugin_dcsr_stepie <= CsrPlugin_csrMapping_writeDataSignal[11];
          CsrPlugin_dcsr_ebreakm <= CsrPlugin_csrMapping_writeDataSignal[15];
        end
      end
      if(execute_CsrPlugin_csr_768) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mstatus_MPIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mstatus_MIE <= CsrPlugin_csrMapping_writeDataSignal[3];
          case(switch_CsrPlugin_l1167)
            2'b11 : begin
              CsrPlugin_mstatus_MPP <= 2'b11;
            end
            default : begin
            end
          endcase
          FpuPlugin_fs <= CsrPlugin_csrMapping_writeDataSignal[14 : 13];
        end
      end
      if(execute_CsrPlugin_csr_772) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mie_MEIE <= CsrPlugin_csrMapping_writeDataSignal[11];
          CsrPlugin_mie_MTIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mie_MSIE <= CsrPlugin_csrMapping_writeDataSignal[3];
        end
      end
      if(execute_CsrPlugin_csr_3) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_rm <= CsrPlugin_csrMapping_writeDataSignal[7 : 5];
          FpuPlugin_flags_NX <= _zz_FpuPlugin_flags_NX[0];
          FpuPlugin_flags_UF <= _zz_FpuPlugin_flags_NX[1];
          FpuPlugin_flags_OF <= _zz_FpuPlugin_flags_NX[2];
          FpuPlugin_flags_DZ <= _zz_FpuPlugin_flags_NX[3];
          FpuPlugin_flags_NV <= _zz_FpuPlugin_flags_NX[4];
        end
      end
      if(execute_CsrPlugin_csr_2) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_rm <= CsrPlugin_csrMapping_writeDataSignal[2 : 0];
        end
      end
      if(execute_CsrPlugin_csr_1) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_flags_NX <= _zz_FpuPlugin_flags_NX_1[0];
          FpuPlugin_flags_UF <= _zz_FpuPlugin_flags_NX_1[1];
          FpuPlugin_flags_OF <= _zz_FpuPlugin_flags_NX_1[2];
          FpuPlugin_flags_DZ <= _zz_FpuPlugin_flags_NX_1[3];
          FpuPlugin_flags_NV <= _zz_FpuPlugin_flags_NX_1[4];
        end
      end
      if(execute_CsrPlugin_csr_256) begin
        if(execute_CsrPlugin_writeEnable) begin
          FpuPlugin_fs <= CsrPlugin_csrMapping_writeDataSignal[14 : 13];
        end
      end
      FpuPlugin_stateReg <= FpuPlugin_stateNext;
      CsrPlugin_running <= CsrPlugin_running_aheadValue;
    end
  end

  always @(posedge io_systemClk) begin
    if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload <= IBusCachedPlugin_iBusRsp_stages_1_output_payload;
    end
    if(IBusCachedPlugin_decompressor_input_valid) begin
      IBusCachedPlugin_decompressor_bufferValidLatch <= IBusCachedPlugin_decompressor_bufferValid;
    end
    if(IBusCachedPlugin_decompressor_input_valid) begin
      IBusCachedPlugin_decompressor_throw2BytesLatch <= IBusCachedPlugin_decompressor_throw2Bytes;
    end
    if(when_Fetcher_l288) begin
      IBusCachedPlugin_decompressor_bufferData <= IBusCachedPlugin_decompressor_input_payload_rsp_inst[31 : 16];
    end
    if(IBusCachedPlugin_decompressor_output_ready) begin
      _zz_IBusCachedPlugin_injector_decodeInput_payload_pc <= IBusCachedPlugin_decompressor_output_payload_pc;
      _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_error <= IBusCachedPlugin_decompressor_output_payload_rsp_error;
      _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst <= IBusCachedPlugin_decompressor_output_payload_rsp_inst;
      _zz_IBusCachedPlugin_injector_decodeInput_payload_isRvc <= IBusCachedPlugin_decompressor_output_payload_isRvc;
    end
    if(IBusCachedPlugin_injector_decodeInput_ready) begin
      IBusCachedPlugin_injector_formal_rawInDecode <= IBusCachedPlugin_decompressor_raw;
    end
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_s1_tightlyCoupledHit <= IBusCachedPlugin_s0_tightlyCoupledHit;
    end
    if(IBusCachedPlugin_iBusRsp_stages_2_input_ready) begin
      IBusCachedPlugin_s2_tightlyCoupledHit <= IBusCachedPlugin_s1_tightlyCoupledHit;
    end
    if(dataCache_2_io_mem_cmd_rValidN) begin
      dataCache_2_io_mem_cmd_rData_wr <= dataCache_2_io_mem_cmd_payload_wr;
      dataCache_2_io_mem_cmd_rData_uncached <= dataCache_2_io_mem_cmd_payload_uncached;
      dataCache_2_io_mem_cmd_rData_address <= dataCache_2_io_mem_cmd_payload_address;
      dataCache_2_io_mem_cmd_rData_data <= dataCache_2_io_mem_cmd_payload_data;
      dataCache_2_io_mem_cmd_rData_mask <= dataCache_2_io_mem_cmd_payload_mask;
      dataCache_2_io_mem_cmd_rData_size <= dataCache_2_io_mem_cmd_payload_size;
      dataCache_2_io_mem_cmd_rData_exclusive <= dataCache_2_io_mem_cmd_payload_exclusive;
      dataCache_2_io_mem_cmd_rData_last <= dataCache_2_io_mem_cmd_payload_last;
    end
    if(dataCache_2_io_mem_cmd_s2mPipe_ready) begin
      dataCache_2_io_mem_cmd_s2mPipe_rData_wr <= dataCache_2_io_mem_cmd_s2mPipe_payload_wr;
      dataCache_2_io_mem_cmd_s2mPipe_rData_uncached <= dataCache_2_io_mem_cmd_s2mPipe_payload_uncached;
      dataCache_2_io_mem_cmd_s2mPipe_rData_address <= dataCache_2_io_mem_cmd_s2mPipe_payload_address;
      dataCache_2_io_mem_cmd_s2mPipe_rData_data <= dataCache_2_io_mem_cmd_s2mPipe_payload_data;
      dataCache_2_io_mem_cmd_s2mPipe_rData_mask <= dataCache_2_io_mem_cmd_s2mPipe_payload_mask;
      dataCache_2_io_mem_cmd_s2mPipe_rData_size <= dataCache_2_io_mem_cmd_s2mPipe_payload_size;
      dataCache_2_io_mem_cmd_s2mPipe_rData_exclusive <= dataCache_2_io_mem_cmd_s2mPipe_payload_exclusive;
      dataCache_2_io_mem_cmd_s2mPipe_rData_last <= dataCache_2_io_mem_cmd_s2mPipe_payload_last;
    end
    dBus_rsp_payload_exclusive_regNext <= dBus_rsp_payload_exclusive;
    dBus_rsp_payload_error_regNext <= dBus_rsp_payload_error;
    dBus_rsp_payload_last_regNext <= dBus_rsp_payload_last;
    dBus_rsp_payload_aggregated_regNext <= dBus_rsp_payload_aggregated;
    if(when_DBusCachedPlugin_l334) begin
      dBus_rsp_payload_data_regNextWhen <= dBus_rsp_payload_data;
    end
    HazardSimplePlugin_writeBackBuffer_payload_address <= HazardSimplePlugin_writeBackWrites_payload_address;
    HazardSimplePlugin_writeBackBuffer_payload_data <= HazardSimplePlugin_writeBackWrites_payload_data;
    if(when_CsrPlugin_l768) begin
      if(_zz_6[0]) begin
        CsrPlugin_dataCsrw_value_0 <= debugBus_dmToHart_payload_data;
      end
      if(_zz_6[1]) begin
        CsrPlugin_dataCsrw_value_1 <= debugBus_dmToHart_payload_data;
      end
    end
    if(CsrPlugin_inject_cmd_toStream_ready) begin
      CsrPlugin_inject_cmd_toStream_rData_op <= CsrPlugin_inject_cmd_toStream_payload_op;
      CsrPlugin_inject_cmd_toStream_rData_address <= CsrPlugin_inject_cmd_toStream_payload_address;
      CsrPlugin_inject_cmd_toStream_rData_data <= CsrPlugin_inject_cmd_toStream_payload_data;
      CsrPlugin_inject_cmd_toStream_rData_size <= CsrPlugin_inject_cmd_toStream_payload_size;
    end
    CsrPlugin_mip_MEIP <= externalInterrupt;
    CsrPlugin_mip_MTIP <= timerInterrupt;
    CsrPlugin_mip_MSIP <= softwareInterrupt;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_code : decodeExceptionPort_payload_code);
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_badAddr : decodeExceptionPort_payload_badAddr);
    end
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= CsrPlugin_selfException_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= CsrPlugin_selfException_payload_badAddr;
    end
    if(DBusCachedPlugin_exceptionBus_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= DBusCachedPlugin_exceptionBus_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= DBusCachedPlugin_exceptionBus_payload_badAddr;
    end
    if(when_CsrPlugin_l1440) begin
      if(when_CsrPlugin_l1446) begin
        CsrPlugin_interrupt_code <= 4'b0111;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l1446_1) begin
        CsrPlugin_interrupt_code <= 4'b0011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l1446_2) begin
        CsrPlugin_interrupt_code <= 4'b1011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
    end
    if(when_CsrPlugin_l1534) begin
      if(when_CsrPlugin_l1542) begin
        case(CsrPlugin_targetPrivilege)
          2'b11 : begin
            CsrPlugin_mcause_interrupt <= (! CsrPlugin_hadException);
            CsrPlugin_mcause_exceptionCode <= CsrPlugin_trapCause;
            CsrPlugin_mepc <= writeBack_PC;
            if(CsrPlugin_hadException) begin
              CsrPlugin_mtval <= CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
            end
          end
          default : begin
          end
        endcase
      end else begin
        if(when_CsrPlugin_l1572) begin
          CsrPlugin_dpc <= writeBack_PC;
        end
      end
    end
    execute_MulPlugin_delayLogic_counter <= (execute_MulPlugin_delayLogic_counter + 1'b1);
    if(when_MulPlugin_l70) begin
      execute_MulPlugin_delayLogic_counter <= 1'b0;
    end
    execute_MulPlugin_withOuputBuffer_mul_ll <= (execute_MulPlugin_aULow * execute_MulPlugin_bULow);
    execute_MulPlugin_withOuputBuffer_mul_lh <= ($signed(execute_MulPlugin_aSLow) * $signed(execute_MulPlugin_bHigh));
    execute_MulPlugin_withOuputBuffer_mul_hl <= ($signed(execute_MulPlugin_aHigh) * $signed(execute_MulPlugin_bSLow));
    execute_MulPlugin_withOuputBuffer_mul_hh <= ($signed(execute_MulPlugin_aHigh) * $signed(execute_MulPlugin_bHigh));
    if(when_MulDivIterativePlugin_l126) begin
      memory_MulDivIterativePlugin_div_done <= 1'b1;
    end
    if(when_MulDivIterativePlugin_l126_1) begin
      memory_MulDivIterativePlugin_div_done <= 1'b0;
    end
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l132) begin
        memory_MulDivIterativePlugin_rs1[31 : 0] <= memory_MulDivIterativePlugin_div_stage_0_outNumerator;
        memory_MulDivIterativePlugin_accumulator[31 : 0] <= memory_MulDivIterativePlugin_div_stage_0_outRemainder;
        if(when_MulDivIterativePlugin_l151) begin
          memory_MulDivIterativePlugin_div_result <= _zz_memory_MulDivIterativePlugin_div_result_1[31:0];
        end
      end
    end
    if(when_MulDivIterativePlugin_l162) begin
      memory_MulDivIterativePlugin_accumulator <= 65'h0;
      memory_MulDivIterativePlugin_rs1 <= ((_zz_memory_MulDivIterativePlugin_rs1 ? (~ _zz_memory_MulDivIterativePlugin_rs1_1) : _zz_memory_MulDivIterativePlugin_rs1_1) + _zz_memory_MulDivIterativePlugin_rs1_2);
      memory_MulDivIterativePlugin_rs2 <= ((_zz_memory_MulDivIterativePlugin_rs2 ? (~ execute_RS2) : execute_RS2) + _zz_memory_MulDivIterativePlugin_rs2_1);
      memory_MulDivIterativePlugin_div_needRevert <= ((_zz_memory_MulDivIterativePlugin_rs1 ^ (_zz_memory_MulDivIterativePlugin_rs2 && (! execute_INSTRUCTION[13]))) && (! (((execute_RS2 == 32'h0) && execute_IS_RS2_SIGNED) && (! execute_INSTRUCTION[13]))));
    end
    if(writeBack_FpuPlugin_commit_ready) begin
      writeBack_FpuPlugin_commit_rData_opcode <= writeBack_FpuPlugin_commit_payload_opcode;
      writeBack_FpuPlugin_commit_rData_rd <= writeBack_FpuPlugin_commit_payload_rd;
      writeBack_FpuPlugin_commit_rData_write <= writeBack_FpuPlugin_commit_payload_write;
      writeBack_FpuPlugin_commit_rData_value <= writeBack_FpuPlugin_commit_payload_value;
    end
    if(CfuPlugin_bus_rsp_ready) begin
      CfuPlugin_bus_rsp_rData_outputs_0 <= CfuPlugin_bus_rsp_payload_outputs_0;
    end
    if(when_Pipeline_l124) begin
      decode_to_execute_PC <= _zz_decode_to_execute_PC;
    end
    if(when_Pipeline_l124_1) begin
      execute_to_memory_PC <= execute_PC;
    end
    if(when_Pipeline_l124_2) begin
      memory_to_writeBack_PC <= memory_PC;
    end
    if(when_Pipeline_l124_3) begin
      decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
    end
    if(when_Pipeline_l124_4) begin
      execute_to_memory_INSTRUCTION <= execute_INSTRUCTION;
    end
    if(when_Pipeline_l124_5) begin
      memory_to_writeBack_INSTRUCTION <= memory_INSTRUCTION;
    end
    if(when_Pipeline_l124_6) begin
      decode_to_execute_FORMAL_PC_NEXT <= decode_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_7) begin
      execute_to_memory_FORMAL_PC_NEXT <= execute_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_8) begin
      memory_to_writeBack_FORMAL_PC_NEXT <= _zz_memory_to_writeBack_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_9) begin
      decode_to_execute_MEMORY_FORCE_CONSTISTENCY <= decode_MEMORY_FORCE_CONSTISTENCY;
    end
    if(when_Pipeline_l124_10) begin
      decode_to_execute_LEGAL_INSTRUCTION <= decode_LEGAL_INSTRUCTION;
    end
    if(when_Pipeline_l124_11) begin
      decode_to_execute_MEMORY_FENCE_WR <= decode_MEMORY_FENCE_WR;
    end
    if(when_Pipeline_l124_12) begin
      decode_to_execute_SRC_USE_SUB_LESS <= decode_SRC_USE_SUB_LESS;
    end
    if(when_Pipeline_l124_13) begin
      decode_to_execute_MEMORY_ENABLE <= decode_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_14) begin
      execute_to_memory_MEMORY_ENABLE <= execute_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_15) begin
      memory_to_writeBack_MEMORY_ENABLE <= memory_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_16) begin
      decode_to_execute_ALU_CTRL <= _zz_decode_to_execute_ALU_CTRL;
    end
    if(when_Pipeline_l124_17) begin
      decode_to_execute_REGFILE_WRITE_VALID <= decode_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_18) begin
      execute_to_memory_REGFILE_WRITE_VALID <= execute_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_19) begin
      memory_to_writeBack_REGFILE_WRITE_VALID <= memory_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_20) begin
      decode_to_execute_BYPASSABLE_EXECUTE_STAGE <= decode_BYPASSABLE_EXECUTE_STAGE;
    end
    if(when_Pipeline_l124_21) begin
      decode_to_execute_BYPASSABLE_MEMORY_STAGE <= decode_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_22) begin
      execute_to_memory_BYPASSABLE_MEMORY_STAGE <= execute_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_23) begin
      decode_to_execute_MEMORY_WR <= decode_MEMORY_WR;
    end
    if(when_Pipeline_l124_24) begin
      execute_to_memory_MEMORY_WR <= execute_MEMORY_WR;
    end
    if(when_Pipeline_l124_25) begin
      memory_to_writeBack_MEMORY_WR <= memory_MEMORY_WR;
    end
    if(when_Pipeline_l124_26) begin
      decode_to_execute_HAS_SIDE_EFFECT <= decode_HAS_SIDE_EFFECT;
    end
    if(when_Pipeline_l124_27) begin
      execute_to_memory_HAS_SIDE_EFFECT <= execute_HAS_SIDE_EFFECT;
    end
    if(when_Pipeline_l124_28) begin
      memory_to_writeBack_HAS_SIDE_EFFECT <= memory_HAS_SIDE_EFFECT;
    end
    if(when_Pipeline_l124_29) begin
      decode_to_execute_MEMORY_LRSC <= decode_MEMORY_LRSC;
    end
    if(when_Pipeline_l124_30) begin
      execute_to_memory_MEMORY_LRSC <= execute_MEMORY_LRSC;
    end
    if(when_Pipeline_l124_31) begin
      memory_to_writeBack_MEMORY_LRSC <= memory_MEMORY_LRSC;
    end
    if(when_Pipeline_l124_32) begin
      decode_to_execute_MEMORY_AMO <= decode_MEMORY_AMO;
    end
    if(when_Pipeline_l124_33) begin
      execute_to_memory_MEMORY_AMO <= execute_MEMORY_AMO;
    end
    if(when_Pipeline_l124_34) begin
      memory_to_writeBack_MEMORY_AMO <= memory_MEMORY_AMO;
    end
    if(when_Pipeline_l124_35) begin
      decode_to_execute_MEMORY_MANAGMENT <= decode_MEMORY_MANAGMENT;
    end
    if(when_Pipeline_l124_36) begin
      decode_to_execute_MEMORY_FENCE <= decode_MEMORY_FENCE;
    end
    if(when_Pipeline_l124_37) begin
      execute_to_memory_MEMORY_FENCE <= execute_MEMORY_FENCE;
    end
    if(when_Pipeline_l124_38) begin
      memory_to_writeBack_MEMORY_FENCE <= memory_MEMORY_FENCE;
    end
    if(when_Pipeline_l124_39) begin
      decode_to_execute_IS_CSR <= decode_IS_CSR;
    end
    if(when_Pipeline_l124_40) begin
      decode_to_execute_ENV_CTRL <= _zz_decode_to_execute_ENV_CTRL;
    end
    if(when_Pipeline_l124_41) begin
      execute_to_memory_ENV_CTRL <= _zz_execute_to_memory_ENV_CTRL;
    end
    if(when_Pipeline_l124_42) begin
      memory_to_writeBack_ENV_CTRL <= _zz_memory_to_writeBack_ENV_CTRL;
    end
    if(when_Pipeline_l124_43) begin
      decode_to_execute_BRANCH_CTRL <= _zz_decode_to_execute_BRANCH_CTRL;
    end
    if(when_Pipeline_l124_44) begin
      decode_to_execute_SRC_LESS_UNSIGNED <= decode_SRC_LESS_UNSIGNED;
    end
    if(when_Pipeline_l124_45) begin
      decode_to_execute_IS_MUL <= decode_IS_MUL;
    end
    if(when_Pipeline_l124_46) begin
      execute_to_memory_IS_MUL <= execute_IS_MUL;
    end
    if(when_Pipeline_l124_47) begin
      memory_to_writeBack_IS_MUL <= memory_IS_MUL;
    end
    if(when_Pipeline_l124_48) begin
      decode_to_execute_IS_DIV <= decode_IS_DIV;
    end
    if(when_Pipeline_l124_49) begin
      execute_to_memory_IS_DIV <= execute_IS_DIV;
    end
    if(when_Pipeline_l124_50) begin
      decode_to_execute_IS_RS1_SIGNED <= decode_IS_RS1_SIGNED;
    end
    if(when_Pipeline_l124_51) begin
      decode_to_execute_IS_RS2_SIGNED <= decode_IS_RS2_SIGNED;
    end
    if(when_Pipeline_l124_52) begin
      decode_to_execute_FPU_COMMIT <= decode_FPU_COMMIT;
    end
    if(when_Pipeline_l124_53) begin
      execute_to_memory_FPU_COMMIT <= execute_FPU_COMMIT;
    end
    if(when_Pipeline_l124_54) begin
      memory_to_writeBack_FPU_COMMIT <= memory_FPU_COMMIT;
    end
    if(when_Pipeline_l124_55) begin
      decode_to_execute_FPU_RSP <= decode_FPU_RSP;
    end
    if(when_Pipeline_l124_56) begin
      execute_to_memory_FPU_RSP <= execute_FPU_RSP;
    end
    if(when_Pipeline_l124_57) begin
      memory_to_writeBack_FPU_RSP <= memory_FPU_RSP;
    end
    if(when_Pipeline_l124_58) begin
      decode_to_execute_FPU_OPCODE <= _zz_decode_to_execute_FPU_OPCODE;
    end
    if(when_Pipeline_l124_59) begin
      execute_to_memory_FPU_OPCODE <= _zz_execute_to_memory_FPU_OPCODE;
    end
    if(when_Pipeline_l124_60) begin
      memory_to_writeBack_FPU_OPCODE <= _zz_memory_to_writeBack_FPU_OPCODE;
    end
    if(when_Pipeline_l124_61) begin
      decode_to_execute_CfuPlugin_CFU_ENABLE <= decode_CfuPlugin_CFU_ENABLE;
    end
    if(when_Pipeline_l124_62) begin
      decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND <= _zz_decode_to_execute_CfuPlugin_CFU_INPUT_2_KIND;
    end
    if(when_Pipeline_l124_63) begin
      decode_to_execute_ALU_BITWISE_CTRL <= _zz_decode_to_execute_ALU_BITWISE_CTRL;
    end
    if(when_Pipeline_l124_64) begin
      decode_to_execute_SHIFT_CTRL <= _zz_decode_to_execute_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_65) begin
      execute_to_memory_SHIFT_CTRL <= _zz_execute_to_memory_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_66) begin
      decode_to_execute_RS1 <= _zz_decode_to_execute_RS1;
    end
    if(when_Pipeline_l124_67) begin
      execute_to_memory_RS1 <= execute_RS1;
    end
    if(when_Pipeline_l124_68) begin
      memory_to_writeBack_RS1 <= memory_RS1;
    end
    if(when_Pipeline_l124_69) begin
      decode_to_execute_RS2 <= _zz_decode_to_execute_RS2;
    end
    if(when_Pipeline_l124_70) begin
      decode_to_execute_SRC2_FORCE_ZERO <= decode_SRC2_FORCE_ZERO;
    end
    if(when_Pipeline_l124_71) begin
      decode_to_execute_SRC1 <= decode_SRC1;
    end
    if(when_Pipeline_l124_72) begin
      decode_to_execute_SRC2 <= decode_SRC2;
    end
    if(when_Pipeline_l124_73) begin
      decode_to_execute_CSR_WRITE_OPCODE <= decode_CSR_WRITE_OPCODE;
    end
    if(when_Pipeline_l124_74) begin
      decode_to_execute_CSR_READ_OPCODE <= decode_CSR_READ_OPCODE;
    end
    if(when_Pipeline_l124_78) begin
      decode_to_execute_FPU_COMMIT_LOAD <= decode_FPU_COMMIT_LOAD;
    end
    if(when_Pipeline_l124_79) begin
      execute_to_memory_FPU_COMMIT_LOAD <= execute_FPU_COMMIT_LOAD;
    end
    if(when_Pipeline_l124_80) begin
      memory_to_writeBack_FPU_COMMIT_LOAD <= memory_FPU_COMMIT_LOAD;
    end
    if(when_Pipeline_l124_81) begin
      execute_to_memory_MEMORY_STORE_DATA_RF <= execute_MEMORY_STORE_DATA_RF;
    end
    if(when_Pipeline_l124_82) begin
      memory_to_writeBack_MEMORY_STORE_DATA_RF <= memory_MEMORY_STORE_DATA_RF;
    end
    if(when_Pipeline_l124_83) begin
      execute_to_memory_MEMORY_VIRTUAL_ADDRESS <= execute_MEMORY_VIRTUAL_ADDRESS;
    end
    if(when_Pipeline_l124_84) begin
      execute_to_memory_BRANCH_DO <= execute_BRANCH_DO;
    end
    if(when_Pipeline_l124_85) begin
      execute_to_memory_BRANCH_CALC <= execute_BRANCH_CALC;
    end
    if(when_Pipeline_l124_86) begin
      execute_to_memory_MUL_LL <= execute_MUL_LL;
    end
    if(when_Pipeline_l124_87) begin
      execute_to_memory_MUL_LH <= execute_MUL_LH;
    end
    if(when_Pipeline_l124_88) begin
      execute_to_memory_MUL_HL <= execute_MUL_HL;
    end
    if(when_Pipeline_l124_89) begin
      execute_to_memory_MUL_HH <= execute_MUL_HH;
    end
    if(when_Pipeline_l124_90) begin
      memory_to_writeBack_MUL_HH <= memory_MUL_HH;
    end
    if(when_Pipeline_l124_93) begin
      execute_to_memory_REGFILE_WRITE_DATA <= _zz_decode_RS2;
    end
    if(when_Pipeline_l124_94) begin
      memory_to_writeBack_REGFILE_WRITE_DATA <= _zz_decode_RS2_1;
    end
    if(when_Pipeline_l124_95) begin
      execute_to_memory_SHIFT_RIGHT <= execute_SHIFT_RIGHT;
    end
    if(when_Pipeline_l124_96) begin
      memory_to_writeBack_MUL_LOW <= memory_MUL_LOW;
    end
    if(when_Fetcher_l411) begin
      _zz_IBusCachedPlugin_injector_decodeInput_payload_rsp_inst <= CsrPlugin_injectionPort_payload;
    end
    if(when_CsrPlugin_l1813) begin
      execute_CsrPlugin_csr_1972 <= (decode_INSTRUCTION[31 : 20] == 12'h7b4);
    end
    if(when_CsrPlugin_l1813_1) begin
      execute_CsrPlugin_csr_1969 <= (decode_INSTRUCTION[31 : 20] == 12'h7b1);
    end
    if(when_CsrPlugin_l1813_2) begin
      execute_CsrPlugin_csr_1968 <= (decode_INSTRUCTION[31 : 20] == 12'h7b0);
    end
    if(when_CsrPlugin_l1813_3) begin
      execute_CsrPlugin_csr_3857 <= (decode_INSTRUCTION[31 : 20] == 12'hf11);
    end
    if(when_CsrPlugin_l1813_4) begin
      execute_CsrPlugin_csr_3858 <= (decode_INSTRUCTION[31 : 20] == 12'hf12);
    end
    if(when_CsrPlugin_l1813_5) begin
      execute_CsrPlugin_csr_3859 <= (decode_INSTRUCTION[31 : 20] == 12'hf13);
    end
    if(when_CsrPlugin_l1813_6) begin
      execute_CsrPlugin_csr_3860 <= (decode_INSTRUCTION[31 : 20] == 12'hf14);
    end
    if(when_CsrPlugin_l1813_7) begin
      execute_CsrPlugin_csr_769 <= (decode_INSTRUCTION[31 : 20] == 12'h301);
    end
    if(when_CsrPlugin_l1813_8) begin
      execute_CsrPlugin_csr_768 <= (decode_INSTRUCTION[31 : 20] == 12'h300);
    end
    if(when_CsrPlugin_l1813_9) begin
      execute_CsrPlugin_csr_836 <= (decode_INSTRUCTION[31 : 20] == 12'h344);
    end
    if(when_CsrPlugin_l1813_10) begin
      execute_CsrPlugin_csr_772 <= (decode_INSTRUCTION[31 : 20] == 12'h304);
    end
    if(when_CsrPlugin_l1813_11) begin
      execute_CsrPlugin_csr_773 <= (decode_INSTRUCTION[31 : 20] == 12'h305);
    end
    if(when_CsrPlugin_l1813_12) begin
      execute_CsrPlugin_csr_833 <= (decode_INSTRUCTION[31 : 20] == 12'h341);
    end
    if(when_CsrPlugin_l1813_13) begin
      execute_CsrPlugin_csr_832 <= (decode_INSTRUCTION[31 : 20] == 12'h340);
    end
    if(when_CsrPlugin_l1813_14) begin
      execute_CsrPlugin_csr_834 <= (decode_INSTRUCTION[31 : 20] == 12'h342);
    end
    if(when_CsrPlugin_l1813_15) begin
      execute_CsrPlugin_csr_835 <= (decode_INSTRUCTION[31 : 20] == 12'h343);
    end
    if(when_CsrPlugin_l1813_16) begin
      execute_CsrPlugin_csr_3 <= (decode_INSTRUCTION[31 : 20] == 12'h003);
    end
    if(when_CsrPlugin_l1813_17) begin
      execute_CsrPlugin_csr_2 <= (decode_INSTRUCTION[31 : 20] == 12'h002);
    end
    if(when_CsrPlugin_l1813_18) begin
      execute_CsrPlugin_csr_1 <= (decode_INSTRUCTION[31 : 20] == 12'h001);
    end
    if(when_CsrPlugin_l1813_19) begin
      execute_CsrPlugin_csr_256 <= (decode_INSTRUCTION[31 : 20] == 12'h100);
    end
    if(execute_CsrPlugin_csr_1969) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_dpc <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    if(execute_CsrPlugin_csr_836) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mip_MSIP <= CsrPlugin_csrMapping_writeDataSignal[3];
      end
    end
    if(execute_CsrPlugin_csr_773) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mtvec_base <= CsrPlugin_csrMapping_writeDataSignal[31 : 2];
      end
    end
    if(execute_CsrPlugin_csr_833) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mepc <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    if(execute_CsrPlugin_csr_832) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mscratch <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
  end


endmodule

//BufferCC_55 replaced by BufferCC_44

//BufferCC_54 replaced by BufferCC_45

//BufferCC_53 replaced by BufferCC_44

//BufferCC_52 replaced by BufferCC_45

//Timer_3 replaced by Timer_2

module Timer_2 (
  input  wire          io_tick,
  input  wire          io_clear,
  input  wire [15:0]   io_limit,
  output wire          io_full,
  output wire [15:0]   io_value,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire       [15:0]   _zz_counter;
  wire       [0:0]    _zz_counter_1;
  reg        [15:0]   counter;
  wire                limitHit;
  reg                 inhibitFull;

  assign _zz_counter_1 = (! limitHit);
  assign _zz_counter = {15'd0, _zz_counter_1};
  assign limitHit = (counter == io_limit);
  assign io_full = ((limitHit && io_tick) && (! inhibitFull));
  assign io_value = counter;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      inhibitFull <= 1'b0;
    end else begin
      if(io_tick) begin
        inhibitFull <= limitHit;
      end
      if(io_clear) begin
        inhibitFull <= 1'b0;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(io_tick) begin
      counter <= (counter + _zz_counter);
    end
    if(io_clear) begin
      counter <= 16'h0;
    end
  end


endmodule

module Prescaler_2 (
  input  wire          io_clear,
  input  wire [23:0]   io_limit,
  output wire          io_overflow,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  reg        [23:0]   counter;
  wire                when_Prescaler_l17;

  assign when_Prescaler_l17 = (io_clear || io_overflow);
  assign io_overflow = (counter == io_limit);
  always @(posedge io_peripheralClk) begin
    counter <= (counter + 24'h000001);
    if(when_Prescaler_l17) begin
      counter <= 24'h0;
    end
  end


endmodule

//Timer_1 replaced by Timer

//Prescaler_1 replaced by Prescaler

module Timer (
  input  wire          io_tick,
  input  wire          io_clear,
  input  wire [11:0]   io_limit,
  output wire          io_full,
  output wire [11:0]   io_value,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  wire       [11:0]   _zz_counter;
  wire       [0:0]    _zz_counter_1;
  reg        [11:0]   counter;
  wire                limitHit;
  reg                 inhibitFull;

  assign _zz_counter_1 = (! limitHit);
  assign _zz_counter = {11'd0, _zz_counter_1};
  assign limitHit = (counter == io_limit);
  assign io_full = ((limitHit && io_tick) && (! inhibitFull));
  assign io_value = counter;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      inhibitFull <= 1'b0;
    end else begin
      if(io_tick) begin
        inhibitFull <= limitHit;
      end
      if(io_clear) begin
        inhibitFull <= 1'b0;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(io_tick) begin
      counter <= (counter + _zz_counter);
    end
    if(io_clear) begin
      counter <= 12'h0;
    end
  end


endmodule

module Prescaler (
  input  wire          io_clear,
  input  wire [7:0]    io_limit,
  output wire          io_overflow,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  reg        [7:0]    counter;
  wire                when_Prescaler_l17;

  assign when_Prescaler_l17 = (io_clear || io_overflow);
  assign io_overflow = (counter == io_limit);
  always @(posedge io_peripheralClk) begin
    counter <= (counter + 8'h01);
    if(when_Prescaler_l17) begin
      counter <= 8'h0;
    end
  end


endmodule

//I2cSlave_2 replaced by I2cSlave

//I2cSlave_1 replaced by I2cSlave

module I2cSlave (
  output wire          io_i2c_sda_write,
  input  wire          io_i2c_sda_read,
  output wire          io_i2c_scl_write,
  input  wire          io_i2c_scl_read,
  input  wire [9:0]    io_config_samplingClockDivider,
  input  wire [19:0]   io_config_timeout,
  input  wire [5:0]    io_config_tsuData,
  input  wire          io_config_timeoutClear,
  output reg  [2:0]    io_bus_cmd_kind,
  output wire          io_bus_cmd_data,
  input  wire          io_bus_rsp_valid,
  input  wire          io_bus_rsp_enable,
  input  wire          io_bus_rsp_data,
  output wire          io_timeout,
  output wire          io_internals_inFrame,
  output wire          io_internals_sdaRead,
  output wire          io_internals_sclRead,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);
  localparam I2cSlaveCmdMode_NONE = 3'd0;
  localparam I2cSlaveCmdMode_START = 3'd1;
  localparam I2cSlaveCmdMode_RESTART = 3'd2;
  localparam I2cSlaveCmdMode_STOP = 3'd3;
  localparam I2cSlaveCmdMode_DROP = 3'd4;
  localparam I2cSlaveCmdMode_DRIVE = 3'd5;
  localparam I2cSlaveCmdMode_READ = 3'd6;

  wire                io_i2c_scl_read_buffercc_io_dataOut;
  wire                io_i2c_sda_read_buffercc_io_dataOut;
  reg        [9:0]    filter_timer_counter;
  wire                filter_timer_tick;
  wire                filter_sampler_sclSync;
  wire                filter_sampler_sdaSync;
  wire                filter_sampler_sclSamples_0;
  wire                filter_sampler_sclSamples_1;
  wire                filter_sampler_sclSamples_2;
  wire                _zz_filter_sampler_sclSamples_0;
  reg                 _zz_filter_sampler_sclSamples_1;
  reg                 _zz_filter_sampler_sclSamples_2;
  wire                filter_sampler_sdaSamples_0;
  wire                filter_sampler_sdaSamples_1;
  wire                filter_sampler_sdaSamples_2;
  wire                _zz_filter_sampler_sdaSamples_0;
  reg                 _zz_filter_sampler_sdaSamples_1;
  reg                 _zz_filter_sampler_sdaSamples_2;
  reg                 filter_sda;
  reg                 filter_scl;
  wire                when_Misc_l82;
  wire                when_Misc_l85;
  wire                sclEdge_rise;
  wire                sclEdge_fall;
  wire                sclEdge_toggle;
  reg                 filter_scl_regNext;
  wire                sdaEdge_rise;
  wire                sdaEdge_fall;
  wire                sdaEdge_toggle;
  reg                 filter_sda_regNext;
  wire                detector_start;
  wire                detector_stop;
  reg        [5:0]    tsuData_counter;
  wire                tsuData_done;
  reg                 tsuData_reset;
  wire                when_I2CSlave_l191;
  reg                 ctrl_inFrame;
  reg                 ctrl_inFrameData;
  reg                 ctrl_sdaWrite;
  reg                 ctrl_sclWrite;
  wire                ctrl_rspBufferIn_valid;
  reg                 ctrl_rspBufferIn_ready;
  wire                ctrl_rspBufferIn_payload_enable;
  wire                ctrl_rspBufferIn_payload_data;
  wire                ctrl_rspBuffer_valid;
  reg                 ctrl_rspBuffer_ready;
  wire                ctrl_rspBuffer_payload_enable;
  wire                ctrl_rspBuffer_payload_data;
  reg                 ctrl_rspBufferIn_rValid;
  reg                 ctrl_rspBufferIn_rData_enable;
  reg                 ctrl_rspBufferIn_rData_data;
  wire                when_Stream_l375;
  wire                ctrl_rspAhead_valid;
  wire                ctrl_rspAhead_payload_enable;
  wire                ctrl_rspAhead_payload_data;
  wire                when_I2CSlave_l241;
  wire                when_I2CSlave_l245;
  wire                when_I2CSlave_l251;
  wire       [2:0]    _zz_io_bus_cmd_kind;
  reg                 timeout_enabled;
  reg        [19:0]   timeout_counter;
  wire                timeout_tick;
  wire                when_I2CSlave_l270;
  wire                when_I2CSlave_l276;
  wire       [2:0]    _zz_io_bus_cmd_kind_1;
  `ifndef SYNTHESIS
  reg [55:0] io_bus_cmd_kind_string;
  reg [55:0] _zz_io_bus_cmd_kind_string;
  reg [55:0] _zz_io_bus_cmd_kind_1_string;
  `endif


  (* keep_hierarchy = "TRUE" *) BufferCC_46 io_i2c_scl_read_buffercc (
    .io_dataIn                      (io_i2c_scl_read                    ), //i
    .io_dataOut                     (io_i2c_scl_read_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                   ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset     )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_46 io_i2c_sda_read_buffercc (
    .io_dataIn                      (io_i2c_sda_read                    ), //i
    .io_dataOut                     (io_i2c_sda_read_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                   ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_bus_cmd_kind)
      I2cSlaveCmdMode_NONE : io_bus_cmd_kind_string = "NONE   ";
      I2cSlaveCmdMode_START : io_bus_cmd_kind_string = "START  ";
      I2cSlaveCmdMode_RESTART : io_bus_cmd_kind_string = "RESTART";
      I2cSlaveCmdMode_STOP : io_bus_cmd_kind_string = "STOP   ";
      I2cSlaveCmdMode_DROP : io_bus_cmd_kind_string = "DROP   ";
      I2cSlaveCmdMode_DRIVE : io_bus_cmd_kind_string = "DRIVE  ";
      I2cSlaveCmdMode_READ : io_bus_cmd_kind_string = "READ   ";
      default : io_bus_cmd_kind_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_io_bus_cmd_kind)
      I2cSlaveCmdMode_NONE : _zz_io_bus_cmd_kind_string = "NONE   ";
      I2cSlaveCmdMode_START : _zz_io_bus_cmd_kind_string = "START  ";
      I2cSlaveCmdMode_RESTART : _zz_io_bus_cmd_kind_string = "RESTART";
      I2cSlaveCmdMode_STOP : _zz_io_bus_cmd_kind_string = "STOP   ";
      I2cSlaveCmdMode_DROP : _zz_io_bus_cmd_kind_string = "DROP   ";
      I2cSlaveCmdMode_DRIVE : _zz_io_bus_cmd_kind_string = "DRIVE  ";
      I2cSlaveCmdMode_READ : _zz_io_bus_cmd_kind_string = "READ   ";
      default : _zz_io_bus_cmd_kind_string = "???????";
    endcase
  end
  always @(*) begin
    case(_zz_io_bus_cmd_kind_1)
      I2cSlaveCmdMode_NONE : _zz_io_bus_cmd_kind_1_string = "NONE   ";
      I2cSlaveCmdMode_START : _zz_io_bus_cmd_kind_1_string = "START  ";
      I2cSlaveCmdMode_RESTART : _zz_io_bus_cmd_kind_1_string = "RESTART";
      I2cSlaveCmdMode_STOP : _zz_io_bus_cmd_kind_1_string = "STOP   ";
      I2cSlaveCmdMode_DROP : _zz_io_bus_cmd_kind_1_string = "DROP   ";
      I2cSlaveCmdMode_DRIVE : _zz_io_bus_cmd_kind_1_string = "DRIVE  ";
      I2cSlaveCmdMode_READ : _zz_io_bus_cmd_kind_1_string = "READ   ";
      default : _zz_io_bus_cmd_kind_1_string = "???????";
    endcase
  end
  `endif

  assign filter_timer_tick = (filter_timer_counter == 10'h0);
  assign filter_sampler_sclSync = io_i2c_scl_read_buffercc_io_dataOut;
  assign filter_sampler_sdaSync = io_i2c_sda_read_buffercc_io_dataOut;
  assign _zz_filter_sampler_sclSamples_0 = filter_sampler_sclSync;
  assign filter_sampler_sclSamples_0 = _zz_filter_sampler_sclSamples_0;
  assign filter_sampler_sclSamples_1 = _zz_filter_sampler_sclSamples_1;
  assign filter_sampler_sclSamples_2 = _zz_filter_sampler_sclSamples_2;
  assign _zz_filter_sampler_sdaSamples_0 = filter_sampler_sdaSync;
  assign filter_sampler_sdaSamples_0 = _zz_filter_sampler_sdaSamples_0;
  assign filter_sampler_sdaSamples_1 = _zz_filter_sampler_sdaSamples_1;
  assign filter_sampler_sdaSamples_2 = _zz_filter_sampler_sdaSamples_2;
  assign when_Misc_l82 = (&{(filter_sampler_sdaSamples_2 != filter_sda),{(filter_sampler_sdaSamples_1 != filter_sda),(filter_sampler_sdaSamples_0 != filter_sda)}});
  assign when_Misc_l85 = (&{(filter_sampler_sclSamples_2 != filter_scl),{(filter_sampler_sclSamples_1 != filter_scl),(filter_sampler_sclSamples_0 != filter_scl)}});
  assign sclEdge_rise = ((! filter_scl_regNext) && filter_scl);
  assign sclEdge_fall = (filter_scl_regNext && (! filter_scl));
  assign sclEdge_toggle = (filter_scl_regNext != filter_scl);
  assign sdaEdge_rise = ((! filter_sda_regNext) && filter_sda);
  assign sdaEdge_fall = (filter_sda_regNext && (! filter_sda));
  assign sdaEdge_toggle = (filter_sda_regNext != filter_sda);
  assign detector_start = (filter_scl && sdaEdge_fall);
  assign detector_stop = (filter_scl && sdaEdge_rise);
  assign tsuData_done = (tsuData_counter == 6'h0);
  always @(*) begin
    tsuData_reset = 1'b0;
    if(ctrl_inFrameData) begin
      tsuData_reset = (! ctrl_rspAhead_valid);
    end
  end

  assign when_I2CSlave_l191 = (! tsuData_done);
  always @(*) begin
    ctrl_sdaWrite = 1'b1;
    if(ctrl_inFrameData) begin
      if(when_I2CSlave_l251) begin
        ctrl_sdaWrite = ctrl_rspAhead_payload_data;
      end
    end
  end

  always @(*) begin
    ctrl_sclWrite = 1'b1;
    if(ctrl_inFrameData) begin
      if(when_I2CSlave_l245) begin
        ctrl_sclWrite = 1'b0;
      end
    end
  end

  always @(*) begin
    ctrl_rspBufferIn_ready = ctrl_rspBuffer_ready;
    if(when_Stream_l375) begin
      ctrl_rspBufferIn_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! ctrl_rspBuffer_valid);
  assign ctrl_rspBuffer_valid = ctrl_rspBufferIn_rValid;
  assign ctrl_rspBuffer_payload_enable = ctrl_rspBufferIn_rData_enable;
  assign ctrl_rspBuffer_payload_data = ctrl_rspBufferIn_rData_data;
  assign ctrl_rspAhead_valid = (ctrl_rspBuffer_valid ? ctrl_rspBuffer_valid : ctrl_rspBufferIn_valid);
  assign ctrl_rspAhead_payload_enable = (ctrl_rspBuffer_valid ? ctrl_rspBuffer_payload_enable : ctrl_rspBufferIn_payload_enable);
  assign ctrl_rspAhead_payload_data = (ctrl_rspBuffer_valid ? ctrl_rspBuffer_payload_data : ctrl_rspBufferIn_payload_data);
  assign ctrl_rspBufferIn_valid = io_bus_rsp_valid;
  assign ctrl_rspBufferIn_payload_enable = io_bus_rsp_enable;
  assign ctrl_rspBufferIn_payload_data = io_bus_rsp_data;
  always @(*) begin
    ctrl_rspBuffer_ready = 1'b0;
    if(ctrl_inFrame) begin
      if(sclEdge_fall) begin
        ctrl_rspBuffer_ready = 1'b1;
      end
    end
  end

  always @(*) begin
    io_bus_cmd_kind = I2cSlaveCmdMode_NONE;
    if(ctrl_inFrame) begin
      if(sclEdge_rise) begin
        io_bus_cmd_kind = I2cSlaveCmdMode_READ;
      end
    end
    if(ctrl_inFrameData) begin
      if(when_I2CSlave_l241) begin
        io_bus_cmd_kind = I2cSlaveCmdMode_DRIVE;
      end
    end
    if(detector_start) begin
      io_bus_cmd_kind = _zz_io_bus_cmd_kind;
    end
    if(when_I2CSlave_l276) begin
      if(ctrl_inFrame) begin
        io_bus_cmd_kind = _zz_io_bus_cmd_kind_1;
      end
    end
  end

  assign io_bus_cmd_data = filter_sda;
  assign when_I2CSlave_l241 = ((! ctrl_rspBuffer_valid) || ctrl_rspBuffer_ready);
  assign when_I2CSlave_l245 = ((! ctrl_rspAhead_valid) || (ctrl_rspAhead_payload_enable && (! tsuData_done)));
  assign when_I2CSlave_l251 = (ctrl_rspAhead_valid && ctrl_rspAhead_payload_enable);
  assign _zz_io_bus_cmd_kind = (ctrl_inFrame ? I2cSlaveCmdMode_RESTART : I2cSlaveCmdMode_START);
  assign timeout_tick = (timeout_enabled && (timeout_counter == 20'h0));
  assign when_I2CSlave_l270 = (((timeout_tick || sclEdge_toggle) || (((! ctrl_inFrame) && filter_scl) && filter_sda)) || io_config_timeoutClear);
  assign io_timeout = timeout_tick;
  assign when_I2CSlave_l276 = (detector_stop || timeout_tick);
  assign _zz_io_bus_cmd_kind_1 = (timeout_tick ? I2cSlaveCmdMode_DROP : I2cSlaveCmdMode_STOP);
  assign io_internals_inFrame = ctrl_inFrame;
  assign io_internals_sdaRead = filter_sda;
  assign io_internals_sclRead = filter_scl;
  assign io_i2c_scl_write = ctrl_sclWrite;
  assign io_i2c_sda_write = ctrl_sdaWrite;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      filter_timer_counter <= 10'h0;
      _zz_filter_sampler_sclSamples_1 <= 1'b1;
      _zz_filter_sampler_sclSamples_2 <= 1'b1;
      _zz_filter_sampler_sdaSamples_1 <= 1'b1;
      _zz_filter_sampler_sdaSamples_2 <= 1'b1;
      filter_sda <= 1'b1;
      filter_scl <= 1'b1;
      filter_scl_regNext <= 1'b1;
      filter_sda_regNext <= 1'b1;
      tsuData_counter <= 6'h0;
      ctrl_inFrame <= 1'b0;
      ctrl_inFrameData <= 1'b0;
      ctrl_rspBufferIn_rValid <= 1'b0;
      timeout_counter <= 20'h0;
    end else begin
      filter_timer_counter <= (filter_timer_counter - 10'h001);
      if(filter_timer_tick) begin
        filter_timer_counter <= io_config_samplingClockDivider;
      end
      if(filter_timer_tick) begin
        _zz_filter_sampler_sclSamples_1 <= _zz_filter_sampler_sclSamples_0;
      end
      if(filter_timer_tick) begin
        _zz_filter_sampler_sclSamples_2 <= _zz_filter_sampler_sclSamples_1;
      end
      if(filter_timer_tick) begin
        _zz_filter_sampler_sdaSamples_1 <= _zz_filter_sampler_sdaSamples_0;
      end
      if(filter_timer_tick) begin
        _zz_filter_sampler_sdaSamples_2 <= _zz_filter_sampler_sdaSamples_1;
      end
      if(filter_timer_tick) begin
        if(when_Misc_l82) begin
          filter_sda <= filter_sampler_sdaSamples_2;
        end
        if(when_Misc_l85) begin
          filter_scl <= filter_sampler_sclSamples_2;
        end
      end
      filter_scl_regNext <= filter_scl;
      filter_sda_regNext <= filter_sda;
      if(when_I2CSlave_l191) begin
        tsuData_counter <= (tsuData_counter - 6'h01);
      end
      if(tsuData_reset) begin
        tsuData_counter <= io_config_tsuData;
      end
      if(ctrl_rspBufferIn_ready) begin
        ctrl_rspBufferIn_rValid <= ctrl_rspBufferIn_valid;
      end
      if(ctrl_inFrame) begin
        if(sclEdge_fall) begin
          ctrl_inFrameData <= 1'b1;
        end
      end
      if(detector_start) begin
        ctrl_inFrame <= 1'b1;
        ctrl_inFrameData <= 1'b0;
      end
      timeout_counter <= (timeout_counter - 20'h00001);
      if(when_I2CSlave_l270) begin
        timeout_counter <= io_config_timeout;
      end
      if(when_I2CSlave_l276) begin
        ctrl_inFrame <= 1'b0;
        ctrl_inFrameData <= 1'b0;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(ctrl_rspBufferIn_ready) begin
      ctrl_rspBufferIn_rData_enable <= ctrl_rspBufferIn_payload_enable;
      ctrl_rspBufferIn_rData_data <= ctrl_rspBufferIn_payload_data;
    end
    timeout_enabled <= (io_config_timeout != 20'h0);
  end


endmodule

//StreamFifo_14 replaced by StreamFifo_12

//StreamFifo_13 replaced by StreamFifo_11

//TopLevel_1 replaced by TopLevel

module StreamFifo_12 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [7:0]    io_push_payload_data,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [7:0]    io_pop_payload_data,
  input  wire          io_flush,
  output wire [8:0]    io_occupancy,
  output wire [8:0]    io_availability,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  reg        [7:0]    logic_ram_spinal_port1;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [8:0]    logic_ptr_push;
  reg        [8:0]    logic_ptr_pop;
  wire       [8:0]    logic_ptr_occupancy;
  wire       [8:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [7:0]    logic_push_onRam_write_payload_address;
  wire       [7:0]    logic_push_onRam_write_payload_data_data;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [7:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [7:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [7:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [7:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [7:0]    logic_pop_sync_readPort_rsp_data;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [7:0]    logic_pop_sync_readArbitation_translated_payload_data;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [8:0]    logic_pop_sync_popReg;
  reg [7:0] logic_ram [0:255];

  always @(posedge io_peripheralClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= logic_push_onRam_write_payload_data_data;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 9'h100) == 9'h0);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[7:0];
  assign logic_push_onRam_write_payload_data_data = io_push_payload_data;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[7:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign logic_pop_sync_readPort_rsp_data = logic_ram_spinal_port1[7 : 0];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_data = logic_pop_sync_readPort_rsp_data;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = logic_pop_sync_readArbitation_translated_payload_data;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (9'h100 - logic_ptr_occupancy);
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      logic_ptr_push <= 9'h0;
      logic_ptr_pop <= 9'h0;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 9'h0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 9'h001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 9'h001);
      end
      if(io_flush) begin
        logic_ptr_push <= 9'h0;
        logic_ptr_pop <= 9'h0;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 9'h0;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module StreamFifo_11 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire          io_push_payload_kind,
  input  wire          io_push_payload_read,
  input  wire          io_push_payload_write,
  input  wire [7:0]    io_push_payload_data,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire          io_pop_payload_kind,
  output wire          io_pop_payload_read,
  output wire          io_pop_payload_write,
  output wire [7:0]    io_pop_payload_data,
  input  wire          io_flush,
  output wire [8:0]    io_occupancy,
  output wire [8:0]    io_availability,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  reg        [10:0]   logic_ram_spinal_port1;
  wire       [10:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [8:0]    logic_ptr_push;
  reg        [8:0]    logic_ptr_pop;
  wire       [8:0]    logic_ptr_occupancy;
  wire       [8:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [7:0]    logic_push_onRam_write_payload_address;
  wire                logic_push_onRam_write_payload_data_kind;
  wire                logic_push_onRam_write_payload_data_read;
  wire                logic_push_onRam_write_payload_data_write;
  wire       [7:0]    logic_push_onRam_write_payload_data_data;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [7:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [7:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [7:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [7:0]    logic_pop_sync_readPort_cmd_payload;
  wire                logic_pop_sync_readPort_rsp_kind;
  wire                logic_pop_sync_readPort_rsp_read;
  wire                logic_pop_sync_readPort_rsp_write;
  wire       [7:0]    logic_pop_sync_readPort_rsp_data;
  wire       [10:0]   _zz_logic_pop_sync_readPort_rsp_kind;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire                logic_pop_sync_readArbitation_translated_payload_kind;
  wire                logic_pop_sync_readArbitation_translated_payload_read;
  wire                logic_pop_sync_readArbitation_translated_payload_write;
  wire       [7:0]    logic_pop_sync_readArbitation_translated_payload_data;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [8:0]    logic_pop_sync_popReg;
  reg [10:0] logic_ram [0:255];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_data,{logic_push_onRam_write_payload_data_write,{logic_push_onRam_write_payload_data_read,logic_push_onRam_write_payload_data_kind}}};
  always @(posedge io_peripheralClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 9'h100) == 9'h0);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[7:0];
  assign logic_push_onRam_write_payload_data_kind = io_push_payload_kind;
  assign logic_push_onRam_write_payload_data_read = io_push_payload_read;
  assign logic_push_onRam_write_payload_data_write = io_push_payload_write;
  assign logic_push_onRam_write_payload_data_data = io_push_payload_data;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[7:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_kind = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_kind = _zz_logic_pop_sync_readPort_rsp_kind[0];
  assign logic_pop_sync_readPort_rsp_read = _zz_logic_pop_sync_readPort_rsp_kind[1];
  assign logic_pop_sync_readPort_rsp_write = _zz_logic_pop_sync_readPort_rsp_kind[2];
  assign logic_pop_sync_readPort_rsp_data = _zz_logic_pop_sync_readPort_rsp_kind[10 : 3];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_kind = logic_pop_sync_readPort_rsp_kind;
  assign logic_pop_sync_readArbitation_translated_payload_read = logic_pop_sync_readPort_rsp_read;
  assign logic_pop_sync_readArbitation_translated_payload_write = logic_pop_sync_readPort_rsp_write;
  assign logic_pop_sync_readArbitation_translated_payload_data = logic_pop_sync_readPort_rsp_data;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_kind = logic_pop_sync_readArbitation_translated_payload_kind;
  assign io_pop_payload_read = logic_pop_sync_readArbitation_translated_payload_read;
  assign io_pop_payload_write = logic_pop_sync_readArbitation_translated_payload_write;
  assign io_pop_payload_data = logic_pop_sync_readArbitation_translated_payload_data;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (9'h100 - logic_ptr_occupancy);
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      logic_ptr_push <= 9'h0;
      logic_ptr_pop <= 9'h0;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 9'h0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 9'h001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 9'h001);
      end
      if(io_flush) begin
        logic_ptr_push <= 9'h0;
        logic_ptr_pop <= 9'h0;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 9'h0;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module TopLevel (
  input  wire          io_config_kind_cpol,
  input  wire          io_config_kind_cpha,
  input  wire [11:0]   io_config_sclkToggle,
  input  wire [1:0]    io_config_mod,
  input  wire [0:0]    io_config_ss_activeHigh,
  input  wire [11:0]   io_config_ss_setup,
  input  wire [11:0]   io_config_ss_hold,
  input  wire [11:0]   io_config_ss_disable,
  input  wire          io_cmd_valid,
  output reg           io_cmd_ready,
  input  wire          io_cmd_payload_kind,
  input  wire          io_cmd_payload_read,
  input  wire          io_cmd_payload_write,
  input  wire [7:0]    io_cmd_payload_data,
  output wire          io_rsp_valid,
  output wire [7:0]    io_rsp_payload_data,
  output wire [0:0]    io_spi_sclk_write,
  output reg           io_spi_data_0_writeEnable,
  input  wire [0:0]    io_spi_data_0_read,
  output reg  [0:0]    io_spi_data_0_write,
  output reg           io_spi_data_1_writeEnable,
  input  wire [0:0]    io_spi_data_1_read,
  output reg  [0:0]    io_spi_data_1_write,
  output reg           io_spi_data_2_writeEnable,
  input  wire [0:0]    io_spi_data_2_read,
  output reg  [0:0]    io_spi_data_2_write,
  output reg           io_spi_data_3_writeEnable,
  input  wire [0:0]    io_spi_data_3_read,
  output reg  [0:0]    io_spi_data_3_write,
  output wire [0:0]    io_spi_ss,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  reg        [0:0]    _zz_outputPhy_dataWrite_3;
  wire       [2:0]    _zz_outputPhy_dataWrite_4;
  reg        [1:0]    _zz_outputPhy_dataWrite_5;
  wire       [1:0]    _zz_outputPhy_dataWrite_6;
  wire       [2:0]    _zz_outputPhy_dataWrite_7;
  reg        [3:0]    _zz_outputPhy_dataWrite_8;
  wire       [0:0]    _zz_outputPhy_dataWrite_9;
  wire       [2:0]    _zz_outputPhy_dataWrite_10;
  wire       [3:0]    _zz_inputPhy_dataRead;
  wire       [3:0]    _zz_inputPhy_dataRead_1;
  wire       [3:0]    _zz_inputPhy_dataRead_2;
  wire       [3:0]    _zz_inputPhy_dataRead_3;
  wire       [3:0]    _zz_inputPhy_dataRead_4;
  wire       [3:0]    _zz_inputPhy_dataRead_5;
  wire       [3:0]    _zz_inputPhy_dataRead_6;
  wire       [8:0]    _zz_inputPhy_bufferNext;
  wire       [10:0]   _zz_inputPhy_bufferNext_1;
  reg        [11:0]   timer_counter;
  reg                 timer_reset;
  wire                timer_ss_setupHit;
  wire                timer_ss_holdHit;
  wire                timer_ss_disableHit;
  wire                timer_sclkToggleHit;
  reg                 fsm_state;
  reg        [2:0]    fsm_counter;
  reg        [2:0]    _zz_fsm_counterPlus;
  wire       [2:0]    fsm_counterPlus;
  reg                 fsm_fastRate;
  reg                 fsm_isDdr;
  reg        [2:0]    fsm_counterMax;
  reg                 fsm_lateSampling;
  reg                 fsm_readFill;
  reg                 fsm_readDone;
  reg        [0:0]    fsm_ss;
  wire                when_SpiXdrMasterCtrl_l741;
  wire                when_SpiXdrMasterCtrl_l744;
  wire                when_SpiXdrMasterCtrl_l751;
  wire                when_SpiXdrMasterCtrl_l753;
  wire                when_SpiXdrMasterCtrl_l760;
  wire                when_SpiXdrMasterCtrl_l766;
  wire                when_SpiXdrMasterCtrl_l783;
  reg        [0:0]    outputPhy_sclkWrite;
  wire       [0:0]    _zz_io_spi_sclk_write;
  wire                when_SpiXdrMasterCtrl_l798;
  reg        [3:0]    outputPhy_dataWrite;
  reg        [2:0]    outputPhy_widthSel;
  reg        [2:0]    outputPhy_offset;
  wire       [7:0]    _zz_outputPhy_dataWrite;
  wire       [7:0]    _zz_outputPhy_dataWrite_1;
  wire       [7:0]    _zz_outputPhy_dataWrite_2;
  wire                when_SpiXdrMasterCtrl_l841;
  wire                when_SpiXdrMasterCtrl_l841_1;
  reg        [1:0]    io_config_mod_delay_1;
  reg        [1:0]    inputPhy_mod;
  reg                 fsm_readFill_delay_1;
  reg                 inputPhy_readFill;
  reg                 fsm_readDone_delay_1;
  reg                 inputPhy_readDone;
  reg        [6:0]    inputPhy_buffer;
  reg        [7:0]    inputPhy_bufferNext;
  reg        [2:0]    inputPhy_widthSel;
  wire       [3:0]    inputPhy_dataWrite;
  reg        [3:0]    inputPhy_dataRead;
  reg                 fsm_state_delay_1;
  reg                 fsm_state_delay_2;
  wire                when_SpiXdrMasterCtrl_l863;
  reg        [3:0]    inputPhy_dataReadBuffer;

  assign _zz_outputPhy_dataWrite_4 = (outputPhy_offset - fsm_counter);
  assign _zz_outputPhy_dataWrite_6 = (_zz_outputPhy_dataWrite_7 >>> 1'd1);
  assign _zz_outputPhy_dataWrite_7 = (outputPhy_offset - fsm_counter);
  assign _zz_outputPhy_dataWrite_9 = (_zz_outputPhy_dataWrite_10 >>> 2'd2);
  assign _zz_outputPhy_dataWrite_10 = (outputPhy_offset - fsm_counter);
  assign _zz_inputPhy_dataRead = {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
  assign _zz_inputPhy_dataRead_1 = {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
  assign _zz_inputPhy_dataRead_2 = {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
  assign _zz_inputPhy_dataRead_3 = {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
  assign _zz_inputPhy_dataRead_4 = {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
  assign _zz_inputPhy_dataRead_5 = {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
  assign _zz_inputPhy_dataRead_6 = {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
  assign _zz_inputPhy_bufferNext = {inputPhy_buffer,inputPhy_dataRead[1 : 0]};
  assign _zz_inputPhy_bufferNext_1 = {inputPhy_buffer,inputPhy_dataRead[3 : 0]};
  always @(*) begin
    case(_zz_outputPhy_dataWrite_4)
      3'b000 : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[0 : 0];
      3'b001 : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[1 : 1];
      3'b010 : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[2 : 2];
      3'b011 : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[3 : 3];
      3'b100 : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[4 : 4];
      3'b101 : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[5 : 5];
      3'b110 : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[6 : 6];
      default : _zz_outputPhy_dataWrite_3 = _zz_outputPhy_dataWrite[7 : 7];
    endcase
  end

  always @(*) begin
    case(_zz_outputPhy_dataWrite_6)
      2'b00 : _zz_outputPhy_dataWrite_5 = _zz_outputPhy_dataWrite_1[1 : 0];
      2'b01 : _zz_outputPhy_dataWrite_5 = _zz_outputPhy_dataWrite_1[3 : 2];
      2'b10 : _zz_outputPhy_dataWrite_5 = _zz_outputPhy_dataWrite_1[5 : 4];
      default : _zz_outputPhy_dataWrite_5 = _zz_outputPhy_dataWrite_1[7 : 6];
    endcase
  end

  always @(*) begin
    case(_zz_outputPhy_dataWrite_9)
      1'b0 : _zz_outputPhy_dataWrite_8 = _zz_outputPhy_dataWrite_2[3 : 0];
      default : _zz_outputPhy_dataWrite_8 = _zz_outputPhy_dataWrite_2[7 : 4];
    endcase
  end

  always @(*) begin
    timer_reset = 1'b0;
    if(io_cmd_valid) begin
      if(when_SpiXdrMasterCtrl_l741) begin
        timer_reset = timer_sclkToggleHit;
      end else begin
        if(!when_SpiXdrMasterCtrl_l760) begin
          if(when_SpiXdrMasterCtrl_l766) begin
            if(timer_ss_holdHit) begin
              timer_reset = 1'b1;
            end
          end
        end
      end
    end
    if(when_SpiXdrMasterCtrl_l783) begin
      timer_reset = 1'b1;
    end
  end

  assign timer_ss_setupHit = (timer_counter == io_config_ss_setup);
  assign timer_ss_holdHit = (timer_counter == io_config_ss_hold);
  assign timer_ss_disableHit = (timer_counter == io_config_ss_disable);
  assign timer_sclkToggleHit = (timer_counter == io_config_sclkToggle);
  always @(*) begin
    _zz_fsm_counterPlus = 3'bxxx;
    case(io_config_mod)
      2'b00 : begin
        _zz_fsm_counterPlus = 3'b001;
      end
      2'b01 : begin
        _zz_fsm_counterPlus = 3'b010;
      end
      2'b10 : begin
        _zz_fsm_counterPlus = 3'b100;
      end
      default : begin
      end
    endcase
  end

  assign fsm_counterPlus = (fsm_counter + _zz_fsm_counterPlus);
  always @(*) begin
    fsm_fastRate = 1'bx;
    case(io_config_mod)
      2'b00 : begin
        fsm_fastRate = 1'b0;
      end
      2'b01 : begin
        fsm_fastRate = 1'b0;
      end
      2'b10 : begin
        fsm_fastRate = 1'b0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_isDdr = 1'bx;
    case(io_config_mod)
      2'b00 : begin
        fsm_isDdr = 1'b0;
      end
      2'b01 : begin
        fsm_isDdr = 1'b0;
      end
      2'b10 : begin
        fsm_isDdr = 1'b0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_counterMax = 3'bxxx;
    case(io_config_mod)
      2'b00 : begin
        fsm_counterMax = 3'b111;
      end
      2'b01 : begin
        fsm_counterMax = 3'b110;
      end
      2'b10 : begin
        fsm_counterMax = 3'b100;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_lateSampling = 1'bx;
    case(io_config_mod)
      2'b00 : begin
        fsm_lateSampling = 1'b1;
      end
      2'b01 : begin
        fsm_lateSampling = 1'b1;
      end
      2'b10 : begin
        fsm_lateSampling = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_readFill = 1'b0;
    if(io_cmd_valid) begin
      if(when_SpiXdrMasterCtrl_l741) begin
        if(when_SpiXdrMasterCtrl_l744) begin
          fsm_readFill = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    fsm_readDone = 1'b0;
    if(io_cmd_valid) begin
      if(when_SpiXdrMasterCtrl_l741) begin
        if(when_SpiXdrMasterCtrl_l744) begin
          fsm_readDone = (io_cmd_payload_read && (fsm_counter == fsm_counterMax));
        end
      end
    end
  end

  assign io_spi_ss = (~ (fsm_ss ^ io_config_ss_activeHigh));
  always @(*) begin
    io_cmd_ready = 1'b0;
    if(io_cmd_valid) begin
      if(when_SpiXdrMasterCtrl_l741) begin
        if(when_SpiXdrMasterCtrl_l751) begin
          if(when_SpiXdrMasterCtrl_l753) begin
            io_cmd_ready = 1'b1;
          end
        end
      end else begin
        if(when_SpiXdrMasterCtrl_l760) begin
          if(timer_ss_setupHit) begin
            io_cmd_ready = 1'b1;
          end
        end else begin
          if(!when_SpiXdrMasterCtrl_l766) begin
            if(timer_ss_disableHit) begin
              io_cmd_ready = 1'b1;
            end
          end
        end
      end
    end
  end

  assign when_SpiXdrMasterCtrl_l741 = (! io_cmd_payload_kind);
  assign when_SpiXdrMasterCtrl_l744 = ((timer_sclkToggleHit && (((! fsm_state) ^ fsm_lateSampling) || fsm_isDdr)) || fsm_fastRate);
  assign when_SpiXdrMasterCtrl_l751 = ((timer_sclkToggleHit && (fsm_state || fsm_isDdr)) || fsm_fastRate);
  assign when_SpiXdrMasterCtrl_l753 = (fsm_counter == fsm_counterMax);
  assign when_SpiXdrMasterCtrl_l760 = io_cmd_payload_data[7];
  assign when_SpiXdrMasterCtrl_l766 = (! fsm_state);
  assign when_SpiXdrMasterCtrl_l783 = ((! io_cmd_valid) || io_cmd_ready);
  always @(*) begin
    outputPhy_sclkWrite = 1'b0;
    if(when_SpiXdrMasterCtrl_l798) begin
      case(io_config_mod)
        2'b00 : begin
          outputPhy_sclkWrite = ((fsm_state ^ io_config_kind_cpha) ? 1'b1 : 1'b0);
        end
        2'b01 : begin
          outputPhy_sclkWrite = ((fsm_state ^ io_config_kind_cpha) ? 1'b1 : 1'b0);
        end
        2'b10 : begin
          outputPhy_sclkWrite = ((fsm_state ^ io_config_kind_cpha) ? 1'b1 : 1'b0);
        end
        default : begin
        end
      endcase
    end
  end

  assign _zz_io_spi_sclk_write[0] = io_config_kind_cpol;
  assign io_spi_sclk_write = (outputPhy_sclkWrite ^ _zz_io_spi_sclk_write);
  assign when_SpiXdrMasterCtrl_l798 = (io_cmd_valid && (! io_cmd_payload_kind));
  always @(*) begin
    outputPhy_widthSel = 3'bxxx;
    case(io_config_mod)
      2'b00 : begin
        outputPhy_widthSel = 3'b000;
      end
      2'b01 : begin
        outputPhy_widthSel = 3'b001;
      end
      2'b10 : begin
        outputPhy_widthSel = 3'b010;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputPhy_offset = 3'bxxx;
    case(io_config_mod)
      2'b00 : begin
        outputPhy_offset = 3'b111;
      end
      2'b01 : begin
        outputPhy_offset = 3'b111;
      end
      2'b10 : begin
        outputPhy_offset = 3'b111;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    outputPhy_dataWrite = 4'bxxxx;
    case(outputPhy_widthSel)
      3'b000 : begin
        outputPhy_dataWrite[0 : 0] = _zz_outputPhy_dataWrite_3;
      end
      3'b001 : begin
        outputPhy_dataWrite[1 : 0] = _zz_outputPhy_dataWrite_5;
      end
      3'b010 : begin
        outputPhy_dataWrite[3 : 0] = _zz_outputPhy_dataWrite_8;
      end
      default : begin
      end
    endcase
  end

  assign _zz_outputPhy_dataWrite = io_cmd_payload_data;
  assign _zz_outputPhy_dataWrite_1 = io_cmd_payload_data;
  assign _zz_outputPhy_dataWrite_2 = io_cmd_payload_data;
  always @(*) begin
    io_spi_data_0_writeEnable = 1'b0;
    case(io_config_mod)
      2'b00 : begin
        io_spi_data_0_writeEnable = 1'b1;
      end
      2'b01 : begin
        if(when_SpiXdrMasterCtrl_l841) begin
          io_spi_data_0_writeEnable = 1'b1;
        end
      end
      2'b10 : begin
        if(when_SpiXdrMasterCtrl_l841_1) begin
          io_spi_data_0_writeEnable = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_spi_data_1_writeEnable = 1'b0;
    case(io_config_mod)
      2'b01 : begin
        if(when_SpiXdrMasterCtrl_l841) begin
          io_spi_data_1_writeEnable = 1'b1;
        end
      end
      2'b10 : begin
        if(when_SpiXdrMasterCtrl_l841_1) begin
          io_spi_data_1_writeEnable = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_spi_data_2_writeEnable = 1'b0;
    case(io_config_mod)
      2'b10 : begin
        if(when_SpiXdrMasterCtrl_l841_1) begin
          io_spi_data_2_writeEnable = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_spi_data_3_writeEnable = 1'b0;
    case(io_config_mod)
      2'b10 : begin
        if(when_SpiXdrMasterCtrl_l841_1) begin
          io_spi_data_3_writeEnable = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_spi_data_0_write = 1'bx;
    case(io_config_mod)
      2'b00 : begin
        io_spi_data_0_write[0] = (outputPhy_dataWrite[0] || (! (io_cmd_valid && io_cmd_payload_write)));
      end
      2'b01 : begin
        io_spi_data_0_write[0] = outputPhy_dataWrite[0];
      end
      2'b10 : begin
        io_spi_data_0_write[0] = outputPhy_dataWrite[0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_spi_data_1_write = 1'bx;
    case(io_config_mod)
      2'b01 : begin
        io_spi_data_1_write[0] = outputPhy_dataWrite[1];
      end
      2'b10 : begin
        io_spi_data_1_write[0] = outputPhy_dataWrite[1];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_spi_data_2_write = 1'bx;
    case(io_config_mod)
      2'b10 : begin
        io_spi_data_2_write[0] = outputPhy_dataWrite[2];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_spi_data_3_write = 1'bx;
    case(io_config_mod)
      2'b10 : begin
        io_spi_data_3_write[0] = outputPhy_dataWrite[3];
      end
      default : begin
      end
    endcase
  end

  assign when_SpiXdrMasterCtrl_l841 = (io_cmd_valid && io_cmd_payload_write);
  assign when_SpiXdrMasterCtrl_l841_1 = (io_cmd_valid && io_cmd_payload_write);
  always @(*) begin
    inputPhy_bufferNext = 8'bxxxxxxxx;
    case(inputPhy_widthSel)
      3'b000 : begin
        inputPhy_bufferNext = {inputPhy_buffer,inputPhy_dataRead[0 : 0]};
      end
      3'b001 : begin
        inputPhy_bufferNext = _zz_inputPhy_bufferNext[7:0];
      end
      3'b010 : begin
        inputPhy_bufferNext = _zz_inputPhy_bufferNext_1[7:0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    inputPhy_widthSel = 3'bxxx;
    case(inputPhy_mod)
      2'b00 : begin
        inputPhy_widthSel = 3'b000;
      end
      2'b01 : begin
        inputPhy_widthSel = 3'b001;
      end
      2'b10 : begin
        inputPhy_widthSel = 3'b010;
      end
      default : begin
      end
    endcase
  end

  assign when_SpiXdrMasterCtrl_l863 = (! fsm_state_delay_2);
  always @(*) begin
    inputPhy_dataRead = 4'bxxxx;
    case(inputPhy_mod)
      2'b00 : begin
        inputPhy_dataRead[0] = _zz_inputPhy_dataRead[1];
      end
      2'b01 : begin
        inputPhy_dataRead[0] = _zz_inputPhy_dataRead_1[0];
        inputPhy_dataRead[1] = _zz_inputPhy_dataRead_2[1];
      end
      2'b10 : begin
        inputPhy_dataRead[0] = _zz_inputPhy_dataRead_3[0];
        inputPhy_dataRead[1] = _zz_inputPhy_dataRead_4[1];
        inputPhy_dataRead[2] = _zz_inputPhy_dataRead_5[2];
        inputPhy_dataRead[3] = _zz_inputPhy_dataRead_6[3];
      end
      default : begin
      end
    endcase
  end

  assign io_rsp_valid = inputPhy_readDone;
  assign io_rsp_payload_data = inputPhy_bufferNext;
  always @(posedge io_peripheralClk) begin
    timer_counter <= (timer_counter + 12'h001);
    if(timer_reset) begin
      timer_counter <= 12'h0;
    end
    io_config_mod_delay_1 <= io_config_mod;
    inputPhy_mod <= io_config_mod_delay_1;
    fsm_state_delay_1 <= fsm_state;
    fsm_state_delay_2 <= fsm_state_delay_1;
    if(when_SpiXdrMasterCtrl_l863) begin
      inputPhy_dataReadBuffer <= {io_spi_data_3_read[0],{io_spi_data_2_read[0],{io_spi_data_1_read[0],io_spi_data_0_read[0]}}};
    end
    case(inputPhy_widthSel)
      3'b000 : begin
        if(inputPhy_readFill) begin
          inputPhy_buffer <= inputPhy_bufferNext[6:0];
        end
      end
      3'b001 : begin
        if(inputPhy_readFill) begin
          inputPhy_buffer <= inputPhy_bufferNext[6:0];
        end
      end
      3'b010 : begin
        if(inputPhy_readFill) begin
          inputPhy_buffer <= inputPhy_bufferNext[6:0];
        end
      end
      default : begin
      end
    endcase
  end

  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      fsm_state <= 1'b0;
      fsm_counter <= 3'b000;
      fsm_ss <= 1'b0;
      fsm_readFill_delay_1 <= 1'b0;
      inputPhy_readFill <= 1'b0;
      fsm_readDone_delay_1 <= 1'b0;
      inputPhy_readDone <= 1'b0;
    end else begin
      if(io_cmd_valid) begin
        if(when_SpiXdrMasterCtrl_l741) begin
          if(timer_sclkToggleHit) begin
            fsm_state <= (! fsm_state);
          end
          if(when_SpiXdrMasterCtrl_l751) begin
            fsm_counter <= fsm_counterPlus;
            if(when_SpiXdrMasterCtrl_l753) begin
              fsm_state <= 1'b0;
            end
          end
        end else begin
          if(when_SpiXdrMasterCtrl_l760) begin
            fsm_ss[0] <= 1'b1;
          end else begin
            if(when_SpiXdrMasterCtrl_l766) begin
              if(timer_ss_holdHit) begin
                fsm_state <= 1'b1;
              end
            end else begin
              fsm_ss[0] <= 1'b0;
            end
          end
        end
      end
      if(when_SpiXdrMasterCtrl_l783) begin
        fsm_state <= 1'b0;
        fsm_counter <= 3'b000;
      end
      fsm_readFill_delay_1 <= fsm_readFill;
      inputPhy_readFill <= fsm_readFill_delay_1;
      fsm_readDone_delay_1 <= fsm_readDone;
      inputPhy_readDone <= fsm_readDone_delay_1;
    end
  end


endmodule

//StreamFifo_10 replaced by StreamFifo_9

module StreamFifo_9 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [7:0]    io_push_payload,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [7:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [7:0]    io_occupancy,
  output wire [7:0]    io_availability,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  reg        [7:0]    logic_ram_spinal_port1;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [7:0]    logic_ptr_push;
  reg        [7:0]    logic_ptr_pop;
  wire       [7:0]    logic_ptr_occupancy;
  wire       [7:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [6:0]    logic_push_onRam_write_payload_address;
  wire       [7:0]    logic_push_onRam_write_payload_data;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [6:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [6:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [6:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [6:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [7:0]    logic_pop_sync_readPort_rsp;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [7:0]    logic_pop_sync_readArbitation_translated_payload;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [7:0]    logic_pop_sync_popReg;
  reg [7:0] logic_ram [0:127];

  always @(posedge io_peripheralClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= logic_push_onRam_write_payload_data;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 8'h80) == 8'h0);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[6:0];
  assign logic_push_onRam_write_payload_data = io_push_payload;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[6:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign logic_pop_sync_readPort_rsp = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload = logic_pop_sync_readPort_rsp;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload = logic_pop_sync_readArbitation_translated_payload;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (8'h80 - logic_ptr_occupancy);
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      logic_ptr_push <= 8'h0;
      logic_ptr_pop <= 8'h0;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 8'h0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 8'h01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 8'h01);
      end
      if(io_flush) begin
        logic_ptr_push <= 8'h0;
        logic_ptr_pop <= 8'h0;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 8'h0;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module UartCtrl (
  input  wire [2:0]    io_config_frame_dataLength,
  input  wire [0:0]    io_config_frame_stop,
  input  wire [1:0]    io_config_frame_parity,
  input  wire [19:0]   io_config_clockDivider,
  input  wire          io_write_valid,
  output reg           io_write_ready,
  input  wire [7:0]    io_write_payload,
  output wire          io_read_valid,
  input  wire          io_read_ready,
  output wire [7:0]    io_read_payload,
  output wire          io_uart_txd,
  input  wire          io_uart_rxd,
  output wire          io_readError,
  input  wire          io_writeBreak,
  output wire          io_readBreak,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;

  wire                tx_io_write_ready;
  wire                tx_io_txd;
  wire                rx_io_read_valid;
  wire       [7:0]    rx_io_read_payload;
  wire                rx_io_rts;
  wire                rx_io_error;
  wire                rx_io_break;
  reg        [19:0]   clockDivider_counter;
  wire                clockDivider_tick;
  reg                 clockDivider_tickReg;
  reg                 io_write_thrown_valid;
  wire                io_write_thrown_ready;
  wire       [7:0]    io_write_thrown_payload;
  `ifndef SYNTHESIS
  reg [23:0] io_config_frame_stop_string;
  reg [31:0] io_config_frame_parity_string;
  `endif


  UartCtrlTx tx (
    .io_configFrame_dataLength      (io_config_frame_dataLength[2:0]), //i
    .io_configFrame_stop            (io_config_frame_stop           ), //i
    .io_configFrame_parity          (io_config_frame_parity[1:0]    ), //i
    .io_samplingTick                (clockDivider_tickReg           ), //i
    .io_write_valid                 (io_write_thrown_valid          ), //i
    .io_write_ready                 (tx_io_write_ready              ), //o
    .io_write_payload               (io_write_thrown_payload[7:0]   ), //i
    .io_cts                         (1'b0                           ), //i
    .io_txd                         (tx_io_txd                      ), //o
    .io_break                       (io_writeBreak                  ), //i
    .io_peripheralClk               (io_peripheralClk               ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset )  //i
  );
  UartCtrlRx rx (
    .io_configFrame_dataLength      (io_config_frame_dataLength[2:0]), //i
    .io_configFrame_stop            (io_config_frame_stop           ), //i
    .io_configFrame_parity          (io_config_frame_parity[1:0]    ), //i
    .io_samplingTick                (clockDivider_tickReg           ), //i
    .io_read_valid                  (rx_io_read_valid               ), //o
    .io_read_ready                  (io_read_ready                  ), //i
    .io_read_payload                (rx_io_read_payload[7:0]        ), //o
    .io_rxd                         (io_uart_rxd                    ), //i
    .io_rts                         (rx_io_rts                      ), //o
    .io_error                       (rx_io_error                    ), //o
    .io_break                       (rx_io_break                    ), //o
    .io_peripheralClk               (io_peripheralClk               ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_config_frame_stop)
      UartStopType_ONE : io_config_frame_stop_string = "ONE";
      UartStopType_TWO : io_config_frame_stop_string = "TWO";
      default : io_config_frame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_config_frame_parity)
      UartParityType_NONE : io_config_frame_parity_string = "NONE";
      UartParityType_EVEN : io_config_frame_parity_string = "EVEN";
      UartParityType_ODD : io_config_frame_parity_string = "ODD ";
      default : io_config_frame_parity_string = "????";
    endcase
  end
  `endif

  assign clockDivider_tick = (clockDivider_counter == 20'h0);
  always @(*) begin
    io_write_thrown_valid = io_write_valid;
    if(rx_io_break) begin
      io_write_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    io_write_ready = io_write_thrown_ready;
    if(rx_io_break) begin
      io_write_ready = 1'b1;
    end
  end

  assign io_write_thrown_payload = io_write_payload;
  assign io_write_thrown_ready = tx_io_write_ready;
  assign io_read_valid = rx_io_read_valid;
  assign io_read_payload = rx_io_read_payload;
  assign io_uart_txd = tx_io_txd;
  assign io_readError = rx_io_error;
  assign io_readBreak = rx_io_break;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      clockDivider_counter <= 20'h0;
      clockDivider_tickReg <= 1'b0;
    end else begin
      clockDivider_tickReg <= clockDivider_tick;
      clockDivider_counter <= (clockDivider_counter - 20'h00001);
      if(clockDivider_tick) begin
        clockDivider_counter <= io_config_clockDivider;
      end
    end
  end


endmodule

module StreamCCByToggle_1 (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire          io_input_payload_last,
  input  wire [0:0]    io_input_payload_fragment_opcode,
  input  wire [31:0]   io_input_payload_fragment_data,
  input  wire [48:0]   io_input_payload_fragment_context,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire [31:0]   io_output_payload_fragment_data,
  output wire [48:0]   io_output_payload_fragment_context,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset,
  input  wire          io_systemClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1
);

  wire                outHitSignal_buffercc_io_dataOut;
  wire                pushArea_target_buffercc_io_dataOut;
  wire                outHitSignal;
  wire                pushArea_hit;
  wire                pushArea_accept;
  reg                 pushArea_target;
  reg                 pushArea_data_last;
  reg        [0:0]    pushArea_data_fragment_opcode;
  reg        [31:0]   pushArea_data_fragment_data;
  reg        [48:0]   pushArea_data_fragment_context;
  wire                io_input_fire;
  wire                popArea_stream_valid;
  reg                 popArea_stream_ready;
  wire                popArea_stream_payload_last;
  wire       [0:0]    popArea_stream_payload_fragment_opcode;
  wire       [31:0]   popArea_stream_payload_fragment_data;
  wire       [48:0]   popArea_stream_payload_fragment_context;
  wire                popArea_target;
  wire                popArea_stream_fire;
  reg                 popArea_hit;
  wire                popArea_stream_m2sPipe_valid;
  wire                popArea_stream_m2sPipe_ready;
  wire                popArea_stream_m2sPipe_payload_last;
  wire       [0:0]    popArea_stream_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   popArea_stream_m2sPipe_payload_fragment_data;
  wire       [48:0]   popArea_stream_m2sPipe_payload_fragment_context;
  reg                 popArea_stream_rValid;
  (* async_reg = "true" *) reg                 popArea_stream_rData_last;
  (* async_reg = "true" *) reg        [0:0]    popArea_stream_rData_fragment_opcode;
  (* async_reg = "true" *) reg        [31:0]   popArea_stream_rData_fragment_data;
  (* async_reg = "true" *) reg        [48:0]   popArea_stream_rData_fragment_context;
  wire                when_Stream_l375;

  (* keep_hierarchy = "TRUE" *) BufferCC_45 outHitSignal_buffercc (
    .io_dataIn                      (outHitSignal                    ), //i
    .io_dataOut                     (outHitSignal_buffercc_io_dataOut), //o
    .io_peripheralClk               (io_peripheralClk                ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset  )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_44 pushArea_target_buffercc (
    .io_dataIn                                                                           (pushArea_target                                                                    ), //i
    .io_dataOut                                                                          (pushArea_target_buffercc_io_dataOut                                                ), //o
    .io_systemClk                                                                        (io_systemClk                                                                       ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1)  //i
  );
  assign pushArea_hit = outHitSignal_buffercc_io_dataOut;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign pushArea_accept = io_input_fire;
  assign io_input_ready = (pushArea_hit == pushArea_target);
  assign popArea_target = pushArea_target_buffercc_io_dataOut;
  assign popArea_stream_fire = (popArea_stream_valid && popArea_stream_ready);
  assign outHitSignal = popArea_hit;
  assign popArea_stream_valid = (popArea_target != popArea_hit);
  assign popArea_stream_payload_last = pushArea_data_last;
  assign popArea_stream_payload_fragment_opcode = pushArea_data_fragment_opcode;
  assign popArea_stream_payload_fragment_data = pushArea_data_fragment_data;
  assign popArea_stream_payload_fragment_context = pushArea_data_fragment_context;
  always @(*) begin
    popArea_stream_ready = popArea_stream_m2sPipe_ready;
    if(when_Stream_l375) begin
      popArea_stream_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popArea_stream_m2sPipe_valid);
  assign popArea_stream_m2sPipe_valid = popArea_stream_rValid;
  assign popArea_stream_m2sPipe_payload_last = popArea_stream_rData_last;
  assign popArea_stream_m2sPipe_payload_fragment_opcode = popArea_stream_rData_fragment_opcode;
  assign popArea_stream_m2sPipe_payload_fragment_data = popArea_stream_rData_fragment_data;
  assign popArea_stream_m2sPipe_payload_fragment_context = popArea_stream_rData_fragment_context;
  assign io_output_valid = popArea_stream_m2sPipe_valid;
  assign popArea_stream_m2sPipe_ready = io_output_ready;
  assign io_output_payload_last = popArea_stream_m2sPipe_payload_last;
  assign io_output_payload_fragment_opcode = popArea_stream_m2sPipe_payload_fragment_opcode;
  assign io_output_payload_fragment_data = popArea_stream_m2sPipe_payload_fragment_data;
  assign io_output_payload_fragment_context = popArea_stream_m2sPipe_payload_fragment_context;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      pushArea_target <= 1'b0;
    end else begin
      if(pushArea_accept) begin
        pushArea_target <= (! pushArea_target);
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(pushArea_accept) begin
      pushArea_data_last <= io_input_payload_last;
      pushArea_data_fragment_opcode <= io_input_payload_fragment_opcode;
      pushArea_data_fragment_data <= io_input_payload_fragment_data;
      pushArea_data_fragment_context <= io_input_payload_fragment_context;
    end
  end

  always @(posedge io_systemClk) begin
    if(system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1) begin
      popArea_hit <= 1'b0;
      popArea_stream_rValid <= 1'b0;
    end else begin
      if(popArea_stream_fire) begin
        popArea_hit <= popArea_target;
      end
      if(popArea_stream_ready) begin
        popArea_stream_rValid <= popArea_stream_valid;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(popArea_stream_fire) begin
      popArea_stream_rData_last <= popArea_stream_payload_last;
      popArea_stream_rData_fragment_opcode <= popArea_stream_payload_fragment_opcode;
      popArea_stream_rData_fragment_data <= popArea_stream_payload_fragment_data;
      popArea_stream_rData_fragment_context <= popArea_stream_payload_fragment_context;
    end
  end


endmodule

module StreamCCByToggle (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire          io_input_payload_last,
  input  wire [0:0]    io_input_payload_fragment_opcode,
  input  wire [31:0]   io_input_payload_fragment_address,
  input  wire [1:0]    io_input_payload_fragment_length,
  input  wire [31:0]   io_input_payload_fragment_data,
  input  wire [3:0]    io_input_payload_fragment_mask,
  input  wire [48:0]   io_input_payload_fragment_context,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire [31:0]   io_output_payload_fragment_address,
  output wire [1:0]    io_output_payload_fragment_length,
  output wire [31:0]   io_output_payload_fragment_data,
  output wire [3:0]    io_output_payload_fragment_mask,
  output wire [48:0]   io_output_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset,
  input  wire          io_peripheralClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1
);

  wire                outHitSignal_buffercc_io_dataOut;
  wire                pushArea_target_buffercc_io_dataOut;
  wire                outHitSignal;
  wire                pushArea_hit;
  wire                pushArea_accept;
  reg                 pushArea_target;
  reg                 pushArea_data_last;
  reg        [0:0]    pushArea_data_fragment_opcode;
  reg        [31:0]   pushArea_data_fragment_address;
  reg        [1:0]    pushArea_data_fragment_length;
  reg        [31:0]   pushArea_data_fragment_data;
  reg        [3:0]    pushArea_data_fragment_mask;
  reg        [48:0]   pushArea_data_fragment_context;
  wire                io_input_fire;
  wire                popArea_stream_valid;
  reg                 popArea_stream_ready;
  wire                popArea_stream_payload_last;
  wire       [0:0]    popArea_stream_payload_fragment_opcode;
  wire       [31:0]   popArea_stream_payload_fragment_address;
  wire       [1:0]    popArea_stream_payload_fragment_length;
  wire       [31:0]   popArea_stream_payload_fragment_data;
  wire       [3:0]    popArea_stream_payload_fragment_mask;
  wire       [48:0]   popArea_stream_payload_fragment_context;
  wire                popArea_target;
  wire                popArea_stream_fire;
  reg                 popArea_hit;
  wire                popArea_stream_m2sPipe_valid;
  wire                popArea_stream_m2sPipe_ready;
  wire                popArea_stream_m2sPipe_payload_last;
  wire       [0:0]    popArea_stream_m2sPipe_payload_fragment_opcode;
  wire       [31:0]   popArea_stream_m2sPipe_payload_fragment_address;
  wire       [1:0]    popArea_stream_m2sPipe_payload_fragment_length;
  wire       [31:0]   popArea_stream_m2sPipe_payload_fragment_data;
  wire       [3:0]    popArea_stream_m2sPipe_payload_fragment_mask;
  wire       [48:0]   popArea_stream_m2sPipe_payload_fragment_context;
  reg                 popArea_stream_rValid;
  (* async_reg = "true" *) reg                 popArea_stream_rData_last;
  (* async_reg = "true" *) reg        [0:0]    popArea_stream_rData_fragment_opcode;
  (* async_reg = "true" *) reg        [31:0]   popArea_stream_rData_fragment_address;
  (* async_reg = "true" *) reg        [1:0]    popArea_stream_rData_fragment_length;
  (* async_reg = "true" *) reg        [31:0]   popArea_stream_rData_fragment_data;
  (* async_reg = "true" *) reg        [3:0]    popArea_stream_rData_fragment_mask;
  (* async_reg = "true" *) reg        [48:0]   popArea_stream_rData_fragment_context;
  wire                when_Stream_l375;

  (* keep_hierarchy = "TRUE" *) BufferCC_41 outHitSignal_buffercc (
    .io_dataIn                  (outHitSignal                    ), //i
    .io_dataOut                 (outHitSignal_buffercc_io_dataOut), //o
    .io_systemClk               (io_systemClk                    ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset      )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_42 pushArea_target_buffercc (
    .io_dataIn                                                                       (pushArea_target                                                                ), //i
    .io_dataOut                                                                      (pushArea_target_buffercc_io_dataOut                                            ), //o
    .io_peripheralClk                                                                (io_peripheralClk                                                               ), //i
    .system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1 (system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1)  //i
  );
  assign pushArea_hit = outHitSignal_buffercc_io_dataOut;
  assign io_input_fire = (io_input_valid && io_input_ready);
  assign pushArea_accept = io_input_fire;
  assign io_input_ready = (pushArea_hit == pushArea_target);
  assign popArea_target = pushArea_target_buffercc_io_dataOut;
  assign popArea_stream_fire = (popArea_stream_valid && popArea_stream_ready);
  assign outHitSignal = popArea_hit;
  assign popArea_stream_valid = (popArea_target != popArea_hit);
  assign popArea_stream_payload_last = pushArea_data_last;
  assign popArea_stream_payload_fragment_opcode = pushArea_data_fragment_opcode;
  assign popArea_stream_payload_fragment_address = pushArea_data_fragment_address;
  assign popArea_stream_payload_fragment_length = pushArea_data_fragment_length;
  assign popArea_stream_payload_fragment_data = pushArea_data_fragment_data;
  assign popArea_stream_payload_fragment_mask = pushArea_data_fragment_mask;
  assign popArea_stream_payload_fragment_context = pushArea_data_fragment_context;
  always @(*) begin
    popArea_stream_ready = popArea_stream_m2sPipe_ready;
    if(when_Stream_l375) begin
      popArea_stream_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popArea_stream_m2sPipe_valid);
  assign popArea_stream_m2sPipe_valid = popArea_stream_rValid;
  assign popArea_stream_m2sPipe_payload_last = popArea_stream_rData_last;
  assign popArea_stream_m2sPipe_payload_fragment_opcode = popArea_stream_rData_fragment_opcode;
  assign popArea_stream_m2sPipe_payload_fragment_address = popArea_stream_rData_fragment_address;
  assign popArea_stream_m2sPipe_payload_fragment_length = popArea_stream_rData_fragment_length;
  assign popArea_stream_m2sPipe_payload_fragment_data = popArea_stream_rData_fragment_data;
  assign popArea_stream_m2sPipe_payload_fragment_mask = popArea_stream_rData_fragment_mask;
  assign popArea_stream_m2sPipe_payload_fragment_context = popArea_stream_rData_fragment_context;
  assign io_output_valid = popArea_stream_m2sPipe_valid;
  assign popArea_stream_m2sPipe_ready = io_output_ready;
  assign io_output_payload_last = popArea_stream_m2sPipe_payload_last;
  assign io_output_payload_fragment_opcode = popArea_stream_m2sPipe_payload_fragment_opcode;
  assign io_output_payload_fragment_address = popArea_stream_m2sPipe_payload_fragment_address;
  assign io_output_payload_fragment_length = popArea_stream_m2sPipe_payload_fragment_length;
  assign io_output_payload_fragment_data = popArea_stream_m2sPipe_payload_fragment_data;
  assign io_output_payload_fragment_mask = popArea_stream_m2sPipe_payload_fragment_mask;
  assign io_output_payload_fragment_context = popArea_stream_m2sPipe_payload_fragment_context;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      pushArea_target <= 1'b0;
    end else begin
      if(pushArea_accept) begin
        pushArea_target <= (! pushArea_target);
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(pushArea_accept) begin
      pushArea_data_last <= io_input_payload_last;
      pushArea_data_fragment_opcode <= io_input_payload_fragment_opcode;
      pushArea_data_fragment_address <= io_input_payload_fragment_address;
      pushArea_data_fragment_length <= io_input_payload_fragment_length;
      pushArea_data_fragment_data <= io_input_payload_fragment_data;
      pushArea_data_fragment_mask <= io_input_payload_fragment_mask;
      pushArea_data_fragment_context <= io_input_payload_fragment_context;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1) begin
      popArea_hit <= 1'b0;
      popArea_stream_rValid <= 1'b0;
    end else begin
      if(popArea_stream_fire) begin
        popArea_hit <= popArea_target;
      end
      if(popArea_stream_ready) begin
        popArea_stream_rValid <= popArea_stream_valid;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(popArea_stream_fire) begin
      popArea_stream_rData_last <= popArea_stream_payload_last;
      popArea_stream_rData_fragment_opcode <= popArea_stream_payload_fragment_opcode;
      popArea_stream_rData_fragment_address <= popArea_stream_payload_fragment_address;
      popArea_stream_rData_fragment_length <= popArea_stream_payload_fragment_length;
      popArea_stream_rData_fragment_data <= popArea_stream_payload_fragment_data;
      popArea_stream_rData_fragment_mask <= popArea_stream_payload_fragment_mask;
      popArea_stream_rData_fragment_context <= popArea_stream_payload_fragment_context;
    end
  end


endmodule

module StreamFifoCC_13 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire          io_push_payload_last,
  input  wire [1:0]    io_push_payload_fragment_source,
  input  wire [0:0]    io_push_payload_fragment_opcode,
  input  wire [31:0]   io_push_payload_fragment_data,
  input  wire [44:0]   io_push_payload_fragment_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire          io_pop_payload_last,
  output wire [1:0]    io_pop_payload_fragment_source,
  output wire [0:0]    io_pop_payload_fragment_opcode,
  output wire [31:0]   io_pop_payload_fragment_data,
  output wire [44:0]   io_pop_payload_fragment_context,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset,
  input  wire          io_systemClk,
  output wire          system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1
);

  reg        [80:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [80:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire                popCC_readPort_rsp_last;
  wire       [1:0]    popCC_readPort_rsp_fragment_source;
  wire       [0:0]    popCC_readPort_rsp_fragment_opcode;
  wire       [31:0]   popCC_readPort_rsp_fragment_data;
  wire       [44:0]   popCC_readPort_rsp_fragment_context;
  wire       [80:0]   _zz_popCC_readPort_rsp_last;
  wire       [79:0]   _zz_popCC_readPort_rsp_fragment_source;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire                popCC_readArbitation_translated_payload_last;
  wire       [1:0]    popCC_readArbitation_translated_payload_fragment_source;
  wire       [0:0]    popCC_readArbitation_translated_payload_fragment_opcode;
  wire       [31:0]   popCC_readArbitation_translated_payload_fragment_data;
  wire       [44:0]   popCC_readArbitation_translated_payload_fragment_context;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [80:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {{io_push_payload_fragment_context,{io_push_payload_fragment_data,{io_push_payload_fragment_opcode,io_push_payload_fragment_source}}},io_push_payload_last};
  always @(posedge io_peripheralClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_systemClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_38 popToPushGray_buffercc (
    .io_dataIn                      (popToPushGray[4:0]                    ), //i
    .io_dataOut                     (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_peripheralClk               (io_peripheralClk                      ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset        )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_39 system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn                      (system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut                     (system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_systemClk                   (io_systemClk                                                                                                    ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset                                                                                  )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_40 pushToPopGray_buffercc (
    .io_dataIn                                                                         (pushToPopGray[4:0]                                                               ), //i
    .io_dataOut                                                                        (pushToPopGray_buffercc_io_dataOut[4:0]                                           ), //o
    .io_systemClk                                                                      (io_systemClk                                                                     ), //i
    .system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized (system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized = system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_last = ram_spinal_port1;
  assign _zz_popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_last[80 : 1];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_last[0];
  assign popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_fragment_source[1 : 0];
  assign popCC_readPort_rsp_fragment_opcode = _zz_popCC_readPort_rsp_fragment_source[2 : 2];
  assign popCC_readPort_rsp_fragment_data = _zz_popCC_readPort_rsp_fragment_source[34 : 3];
  assign popCC_readPort_rsp_fragment_context = _zz_popCC_readPort_rsp_fragment_source[79 : 35];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign popCC_readArbitation_translated_payload_fragment_source = popCC_readPort_rsp_fragment_source;
  assign popCC_readArbitation_translated_payload_fragment_opcode = popCC_readPort_rsp_fragment_opcode;
  assign popCC_readArbitation_translated_payload_fragment_data = popCC_readPort_rsp_fragment_data;
  assign popCC_readArbitation_translated_payload_fragment_context = popCC_readPort_rsp_fragment_context;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign io_pop_payload_fragment_source = popCC_readArbitation_translated_payload_fragment_source;
  assign io_pop_payload_fragment_opcode = popCC_readArbitation_translated_payload_fragment_opcode;
  assign io_pop_payload_fragment_data = popCC_readArbitation_translated_payload_fragment_data;
  assign io_pop_payload_fragment_context = popCC_readArbitation_translated_payload_fragment_context;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1 = system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_12 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire          io_push_payload_last,
  input  wire [1:0]    io_push_payload_fragment_source,
  input  wire [0:0]    io_push_payload_fragment_opcode,
  input  wire [31:0]   io_push_payload_fragment_address,
  input  wire [5:0]    io_push_payload_fragment_length,
  input  wire [31:0]   io_push_payload_fragment_data,
  input  wire [3:0]    io_push_payload_fragment_mask,
  input  wire [44:0]   io_push_payload_fragment_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire          io_pop_payload_last,
  output wire [1:0]    io_pop_payload_fragment_source,
  output wire [0:0]    io_pop_payload_fragment_opcode,
  output wire [31:0]   io_pop_payload_fragment_address,
  output wire [5:0]    io_pop_payload_fragment_length,
  output wire [31:0]   io_pop_payload_fragment_data,
  output wire [3:0]    io_pop_payload_fragment_mask,
  output wire [44:0]   io_pop_payload_fragment_context,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset,
  input  wire          io_peripheralClk,
  output wire          system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1
);

  reg        [122:0]  ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [122:0]  _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire                popCC_readPort_rsp_last;
  wire       [1:0]    popCC_readPort_rsp_fragment_source;
  wire       [0:0]    popCC_readPort_rsp_fragment_opcode;
  wire       [31:0]   popCC_readPort_rsp_fragment_address;
  wire       [5:0]    popCC_readPort_rsp_fragment_length;
  wire       [31:0]   popCC_readPort_rsp_fragment_data;
  wire       [3:0]    popCC_readPort_rsp_fragment_mask;
  wire       [44:0]   popCC_readPort_rsp_fragment_context;
  wire       [122:0]  _zz_popCC_readPort_rsp_last;
  wire       [121:0]  _zz_popCC_readPort_rsp_fragment_source;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire                popCC_readArbitation_translated_payload_last;
  wire       [1:0]    popCC_readArbitation_translated_payload_fragment_source;
  wire       [0:0]    popCC_readArbitation_translated_payload_fragment_opcode;
  wire       [31:0]   popCC_readArbitation_translated_payload_fragment_address;
  wire       [5:0]    popCC_readArbitation_translated_payload_fragment_length;
  wire       [31:0]   popCC_readArbitation_translated_payload_fragment_data;
  wire       [3:0]    popCC_readArbitation_translated_payload_fragment_mask;
  wire       [44:0]   popCC_readArbitation_translated_payload_fragment_context;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [122:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {{io_push_payload_fragment_context,{io_push_payload_fragment_mask,{io_push_payload_fragment_data,{io_push_payload_fragment_length,{io_push_payload_fragment_address,{io_push_payload_fragment_opcode,io_push_payload_fragment_source}}}}}},io_push_payload_last};
  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_35 popToPushGray_buffercc (
    .io_dataIn                  (popToPushGray[4:0]                    ), //i
    .io_dataOut                 (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_systemClk               (io_systemClk                          ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset            )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_36 system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn                  (system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut                 (system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_peripheralClk           (io_peripheralClk                                                                                            ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                                                                                  )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_37 pushToPopGray_buffercc (
    .io_dataIn                                                                     (pushToPopGray[4:0]                                                           ), //i
    .io_dataOut                                                                    (pushToPopGray_buffercc_io_dataOut[4:0]                                       ), //o
    .io_peripheralClk                                                              (io_peripheralClk                                                             ), //i
    .system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized (system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized = system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_last = ram_spinal_port1;
  assign _zz_popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_last[122 : 1];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_last[0];
  assign popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_fragment_source[1 : 0];
  assign popCC_readPort_rsp_fragment_opcode = _zz_popCC_readPort_rsp_fragment_source[2 : 2];
  assign popCC_readPort_rsp_fragment_address = _zz_popCC_readPort_rsp_fragment_source[34 : 3];
  assign popCC_readPort_rsp_fragment_length = _zz_popCC_readPort_rsp_fragment_source[40 : 35];
  assign popCC_readPort_rsp_fragment_data = _zz_popCC_readPort_rsp_fragment_source[72 : 41];
  assign popCC_readPort_rsp_fragment_mask = _zz_popCC_readPort_rsp_fragment_source[76 : 73];
  assign popCC_readPort_rsp_fragment_context = _zz_popCC_readPort_rsp_fragment_source[121 : 77];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign popCC_readArbitation_translated_payload_fragment_source = popCC_readPort_rsp_fragment_source;
  assign popCC_readArbitation_translated_payload_fragment_opcode = popCC_readPort_rsp_fragment_opcode;
  assign popCC_readArbitation_translated_payload_fragment_address = popCC_readPort_rsp_fragment_address;
  assign popCC_readArbitation_translated_payload_fragment_length = popCC_readPort_rsp_fragment_length;
  assign popCC_readArbitation_translated_payload_fragment_data = popCC_readPort_rsp_fragment_data;
  assign popCC_readArbitation_translated_payload_fragment_mask = popCC_readPort_rsp_fragment_mask;
  assign popCC_readArbitation_translated_payload_fragment_context = popCC_readPort_rsp_fragment_context;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign io_pop_payload_fragment_source = popCC_readArbitation_translated_payload_fragment_source;
  assign io_pop_payload_fragment_opcode = popCC_readArbitation_translated_payload_fragment_opcode;
  assign io_pop_payload_fragment_address = popCC_readArbitation_translated_payload_fragment_address;
  assign io_pop_payload_fragment_length = popCC_readArbitation_translated_payload_fragment_length;
  assign io_pop_payload_fragment_data = popCC_readArbitation_translated_payload_fragment_data;
  assign io_pop_payload_fragment_mask = popCC_readArbitation_translated_payload_fragment_mask;
  assign io_pop_payload_fragment_context = popCC_readArbitation_translated_payload_fragment_context;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1 = system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamArbiter_9 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire          io_inputs_0_payload_last,
  input  wire [1:0]    io_inputs_0_payload_fragment_source,
  input  wire [0:0]    io_inputs_0_payload_fragment_opcode,
  input  wire [63:0]   io_inputs_0_payload_fragment_data,
  input  wire [43:0]   io_inputs_0_payload_fragment_context,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire          io_inputs_1_payload_last,
  input  wire [1:0]    io_inputs_1_payload_fragment_source,
  input  wire [0:0]    io_inputs_1_payload_fragment_opcode,
  input  wire [63:0]   io_inputs_1_payload_fragment_data,
  input  wire [43:0]   io_inputs_1_payload_fragment_context,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire          io_inputs_2_payload_last,
  input  wire [1:0]    io_inputs_2_payload_fragment_source,
  input  wire [0:0]    io_inputs_2_payload_fragment_opcode,
  input  wire [63:0]   io_inputs_2_payload_fragment_data,
  input  wire [43:0]   io_inputs_2_payload_fragment_context,
  input  wire          io_inputs_3_valid,
  output wire          io_inputs_3_ready,
  input  wire          io_inputs_3_payload_last,
  input  wire [1:0]    io_inputs_3_payload_fragment_source,
  input  wire [0:0]    io_inputs_3_payload_fragment_opcode,
  input  wire [63:0]   io_inputs_3_payload_fragment_data,
  input  wire [43:0]   io_inputs_3_payload_fragment_context,
  input  wire          io_inputs_4_valid,
  output wire          io_inputs_4_ready,
  input  wire          io_inputs_4_payload_last,
  input  wire [1:0]    io_inputs_4_payload_fragment_source,
  input  wire [0:0]    io_inputs_4_payload_fragment_opcode,
  input  wire [63:0]   io_inputs_4_payload_fragment_data,
  input  wire [43:0]   io_inputs_4_payload_fragment_context,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [1:0]    io_output_payload_fragment_source,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire [63:0]   io_output_payload_fragment_data,
  output wire [43:0]   io_output_payload_fragment_context,
  output wire [2:0]    io_chosen,
  output wire [4:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [9:0]    _zz__zz_maskProposal_0_2;
  wire       [9:0]    _zz__zz_maskProposal_0_2_1;
  wire       [4:0]    _zz__zz_maskProposal_0_2_2;
  reg                 _zz_io_output_payload_last_3;
  reg        [1:0]    _zz_io_output_payload_fragment_source;
  reg        [0:0]    _zz_io_output_payload_fragment_opcode;
  reg        [63:0]   _zz_io_output_payload_fragment_data;
  reg        [43:0]   _zz_io_output_payload_fragment_context;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  wire                maskProposal_3;
  wire                maskProposal_4;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  reg                 maskLocked_3;
  reg                 maskLocked_4;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire                maskRouted_3;
  wire                maskRouted_4;
  wire       [4:0]    _zz_maskProposal_0;
  wire       [9:0]    _zz_maskProposal_0_1;
  wire       [9:0]    _zz_maskProposal_0_2;
  wire       [4:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                when_Stream_l683;
  wire                _zz_io_output_payload_last;
  wire                _zz_io_output_payload_last_1;
  wire       [2:0]    _zz_io_output_payload_last_2;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  wire                _zz_io_chosen_2;
  wire                _zz_io_chosen_3;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_3,{maskLocked_2,{maskLocked_1,{maskLocked_0,maskLocked_4}}}};
  assign _zz__zz_maskProposal_0_2_1 = {5'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(_zz_io_output_payload_last_2)
      3'b000 : begin
        _zz_io_output_payload_last_3 = io_inputs_0_payload_last;
        _zz_io_output_payload_fragment_source = io_inputs_0_payload_fragment_source;
        _zz_io_output_payload_fragment_opcode = io_inputs_0_payload_fragment_opcode;
        _zz_io_output_payload_fragment_data = io_inputs_0_payload_fragment_data;
        _zz_io_output_payload_fragment_context = io_inputs_0_payload_fragment_context;
      end
      3'b001 : begin
        _zz_io_output_payload_last_3 = io_inputs_1_payload_last;
        _zz_io_output_payload_fragment_source = io_inputs_1_payload_fragment_source;
        _zz_io_output_payload_fragment_opcode = io_inputs_1_payload_fragment_opcode;
        _zz_io_output_payload_fragment_data = io_inputs_1_payload_fragment_data;
        _zz_io_output_payload_fragment_context = io_inputs_1_payload_fragment_context;
      end
      3'b010 : begin
        _zz_io_output_payload_last_3 = io_inputs_2_payload_last;
        _zz_io_output_payload_fragment_source = io_inputs_2_payload_fragment_source;
        _zz_io_output_payload_fragment_opcode = io_inputs_2_payload_fragment_opcode;
        _zz_io_output_payload_fragment_data = io_inputs_2_payload_fragment_data;
        _zz_io_output_payload_fragment_context = io_inputs_2_payload_fragment_context;
      end
      3'b011 : begin
        _zz_io_output_payload_last_3 = io_inputs_3_payload_last;
        _zz_io_output_payload_fragment_source = io_inputs_3_payload_fragment_source;
        _zz_io_output_payload_fragment_opcode = io_inputs_3_payload_fragment_opcode;
        _zz_io_output_payload_fragment_data = io_inputs_3_payload_fragment_data;
        _zz_io_output_payload_fragment_context = io_inputs_3_payload_fragment_context;
      end
      default : begin
        _zz_io_output_payload_last_3 = io_inputs_4_payload_last;
        _zz_io_output_payload_fragment_source = io_inputs_4_payload_fragment_source;
        _zz_io_output_payload_fragment_opcode = io_inputs_4_payload_fragment_opcode;
        _zz_io_output_payload_fragment_data = io_inputs_4_payload_fragment_data;
        _zz_io_output_payload_fragment_context = io_inputs_4_payload_fragment_context;
      end
    endcase
  end

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign maskRouted_3 = (locked ? maskLocked_3 : maskProposal_3);
  assign maskRouted_4 = (locked ? maskLocked_4 : maskProposal_4);
  assign _zz_maskProposal_0 = {io_inputs_4_valid,{io_inputs_3_valid,{io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}}}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[9 : 5] | _zz_maskProposal_0_2[4 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign maskProposal_3 = _zz_maskProposal_0_3[3];
  assign maskProposal_4 = _zz_maskProposal_0_3[4];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l683 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = (((((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2)) || (io_inputs_3_valid && maskRouted_3)) || (io_inputs_4_valid && maskRouted_4));
  assign _zz_io_output_payload_last = (maskRouted_1 || maskRouted_3);
  assign _zz_io_output_payload_last_1 = (maskRouted_2 || maskRouted_3);
  assign _zz_io_output_payload_last_2 = {maskRouted_4,{_zz_io_output_payload_last_1,_zz_io_output_payload_last}};
  assign io_output_payload_last = _zz_io_output_payload_last_3;
  assign io_output_payload_fragment_source = _zz_io_output_payload_fragment_source;
  assign io_output_payload_fragment_opcode = _zz_io_output_payload_fragment_opcode;
  assign io_output_payload_fragment_data = _zz_io_output_payload_fragment_data;
  assign io_output_payload_fragment_context = _zz_io_output_payload_fragment_context;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_inputs_3_ready = (maskRouted_3 && io_output_ready);
  assign io_inputs_4_ready = (maskRouted_4 && io_output_ready);
  assign io_chosenOH = {maskRouted_4,{maskRouted_3,{maskRouted_2,{maskRouted_1,maskRouted_0}}}};
  assign _zz_io_chosen = io_chosenOH[3];
  assign _zz_io_chosen_1 = io_chosenOH[4];
  assign _zz_io_chosen_2 = (io_chosenOH[1] || _zz_io_chosen);
  assign _zz_io_chosen_3 = (io_chosenOH[2] || _zz_io_chosen);
  assign io_chosen = {_zz_io_chosen_1,{_zz_io_chosen_3,_zz_io_chosen_2}};
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b0;
      maskLocked_3 <= 1'b0;
      maskLocked_4 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
        maskLocked_3 <= maskRouted_3;
        maskLocked_4 <= maskRouted_4;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l683) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module BmbErrorSlave (
  input  wire          io_input_cmd_valid,
  output reg           io_input_cmd_ready,
  input  wire          io_input_cmd_payload_last,
  input  wire [1:0]    io_input_cmd_payload_fragment_source,
  input  wire [0:0]    io_input_cmd_payload_fragment_opcode,
  input  wire [31:0]   io_input_cmd_payload_fragment_address,
  input  wire [5:0]    io_input_cmd_payload_fragment_length,
  input  wire [63:0]   io_input_cmd_payload_fragment_data,
  input  wire [7:0]    io_input_cmd_payload_fragment_mask,
  input  wire [43:0]   io_input_cmd_payload_fragment_context,
  output reg           io_input_rsp_valid,
  input  wire          io_input_rsp_ready,
  output wire          io_input_rsp_payload_last,
  output wire [1:0]    io_input_rsp_payload_fragment_source,
  output wire [0:0]    io_input_rsp_payload_fragment_opcode,
  output wire [63:0]   io_input_rsp_payload_fragment_data,
  output wire [43:0]   io_input_rsp_payload_fragment_context,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg                 busy;
  reg        [2:0]    beats;
  reg        [1:0]    source;
  reg        [43:0]   context_1;
  reg        [0:0]    opcode;
  wire                when_BmbDecoder_l122;

  assign io_input_rsp_payload_fragment_opcode = 1'b1;
  assign io_input_rsp_payload_fragment_source = source;
  assign io_input_rsp_payload_fragment_context = context_1;
  assign io_input_rsp_payload_fragment_data = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  assign io_input_rsp_payload_last = ((beats == 3'b000) || (opcode == 1'b1));
  assign when_BmbDecoder_l122 = (! busy);
  always @(*) begin
    if(when_BmbDecoder_l122) begin
      io_input_cmd_ready = 1'b1;
    end else begin
      io_input_cmd_ready = 1'b0;
    end
  end

  always @(*) begin
    if(when_BmbDecoder_l122) begin
      io_input_rsp_valid = 1'b0;
    end else begin
      io_input_rsp_valid = 1'b1;
    end
  end

  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      busy <= 1'b0;
    end else begin
      if(when_BmbDecoder_l122) begin
        busy <= (io_input_cmd_valid && io_input_cmd_payload_last);
      end else begin
        if(io_input_rsp_ready) begin
          if(io_input_rsp_payload_last) begin
            busy <= 1'b0;
          end
        end
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(when_BmbDecoder_l122) begin
      beats <= io_input_cmd_payload_fragment_length[5 : 3];
      source <= io_input_cmd_payload_fragment_source;
      context_1 <= io_input_cmd_payload_fragment_context;
      opcode <= io_input_cmd_payload_fragment_opcode;
    end else begin
      if(io_input_rsp_ready) begin
        beats <= (beats - 3'b001);
      end
    end
  end


endmodule

//StreamFifo_8 replaced by StreamFifo_7

module StreamFifo_7 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [1:0]    io_push_payload_source,
  input  wire [44:0]   io_push_payload_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [1:0]    io_pop_payload_source,
  output wire [44:0]   io_pop_payload_context,
  input  wire          io_flush,
  output wire [3:0]    io_occupancy,
  output wire [3:0]    io_availability,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  reg        [46:0]   logic_ram_spinal_port1;
  wire       [46:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [3:0]    logic_ptr_push;
  reg        [3:0]    logic_ptr_pop;
  wire       [3:0]    logic_ptr_occupancy;
  wire       [3:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [2:0]    logic_push_onRam_write_payload_address;
  wire       [1:0]    logic_push_onRam_write_payload_data_source;
  wire       [44:0]   logic_push_onRam_write_payload_data_context;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [2:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [2:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [2:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [2:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [1:0]    logic_pop_sync_readPort_rsp_source;
  wire       [44:0]   logic_pop_sync_readPort_rsp_context;
  wire       [46:0]   _zz_logic_pop_sync_readPort_rsp_source;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [1:0]    logic_pop_sync_readArbitation_translated_payload_source;
  wire       [44:0]   logic_pop_sync_readArbitation_translated_payload_context;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [3:0]    logic_pop_sync_popReg;
  reg [46:0] logic_ram [0:7];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_context,logic_push_onRam_write_payload_data_source};
  always @(posedge io_peripheralClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 4'b1000) == 4'b0000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[2:0];
  assign logic_push_onRam_write_payload_data_source = io_push_payload_source;
  assign logic_push_onRam_write_payload_data_context = io_push_payload_context;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[2:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_source = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_source = _zz_logic_pop_sync_readPort_rsp_source[1 : 0];
  assign logic_pop_sync_readPort_rsp_context = _zz_logic_pop_sync_readPort_rsp_source[46 : 2];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_source = logic_pop_sync_readPort_rsp_source;
  assign logic_pop_sync_readArbitation_translated_payload_context = logic_pop_sync_readPort_rsp_context;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_source = logic_pop_sync_readArbitation_translated_payload_source;
  assign io_pop_payload_context = logic_pop_sync_readArbitation_translated_payload_context;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (4'b1000 - logic_ptr_occupancy);
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      logic_ptr_push <= 4'b0000;
      logic_ptr_pop <= 4'b0000;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 4'b0000;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 4'b0001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 4'b0001);
      end
      if(io_flush) begin
        logic_ptr_push <= 4'b0000;
        logic_ptr_pop <= 4'b0000;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 4'b0000;
      end
    end
  end

  always @(posedge io_peripheralClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module StreamFifo_6 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [7:0]    io_push_payload_len,
  output reg           io_pop_valid,
  input  wire          io_pop_ready,
  output reg  [7:0]    io_pop_payload_len,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_ddrAReset_reset
);

  wire       [7:0]    logic_ram_spinal_port1;
  wire       [7:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  reg                 logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [7:0]    logic_push_onRam_write_payload_data_len;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [7:0]    logic_pop_async_readed_len;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [7:0]    logic_pop_addressGen_translated_payload_len;
  (* ram_style = "distributed" *) reg [7:0] logic_ram [0:3];

  assign _zz_logic_ram_port = logic_push_onRam_write_payload_data_len;
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  assign logic_ram_spinal_port1 = logic_ram[logic_pop_addressGen_payload];
  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 3'b100) == 3'b000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  always @(*) begin
    logic_ptr_doPush = io_push_fire;
    if(logic_ptr_empty) begin
      if(io_pop_ready) begin
        logic_ptr_doPush = 1'b0;
      end
    end
  end

  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[1:0];
  assign logic_push_onRam_write_payload_data_len = io_push_payload_len;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[1:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign logic_pop_async_readed_len = logic_ram_spinal_port1[7 : 0];
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload_len = logic_pop_async_readed_len;
  always @(*) begin
    io_pop_valid = logic_pop_addressGen_translated_valid;
    if(logic_ptr_empty) begin
      io_pop_valid = io_push_valid;
    end
  end

  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  always @(*) begin
    io_pop_payload_len = logic_pop_addressGen_translated_payload_len;
    if(logic_ptr_empty) begin
      io_pop_payload_len = io_push_payload_len;
    end
  end

  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b100 - logic_ptr_occupancy);
  always @(posedge io_memoryClk or posedge system_ddr_ddrLogic_ddrAReset_reset) begin
    if(system_ddr_ddrLogic_ddrAReset_reset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
    end
  end


endmodule

module Axi4WriteOnlyUpsizer_1 (
  input  wire          io_input_aw_valid,
  output reg           io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [3:0]    io_input_aw_payload_region,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire [0:0]    io_input_aw_payload_lock,
  input  wire [3:0]    io_input_aw_payload_cache,
  input  wire [3:0]    io_input_aw_payload_qos,
  input  wire [2:0]    io_input_aw_payload_prot,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [63:0]   io_input_w_payload_data,
  input  wire [7:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output wire [3:0]    io_input_b_payload_id,
  output wire [1:0]    io_input_b_payload_resp,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [3:0]    io_output_aw_payload_id,
  output wire [3:0]    io_output_aw_payload_region,
  output reg  [7:0]    io_output_aw_payload_len,
  output reg  [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire [0:0]    io_output_aw_payload_lock,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [3:0]    io_output_aw_payload_qos,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [127:0]  io_output_w_payload_data,
  output wire [15:0]   io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [3:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire       [14:0]   _zz_cmdLogic_byteCount;
  wire       [11:0]   _zz_cmdLogic_incrLen;
  wire       [11:0]   _zz_cmdLogic_incrLen_1;
  wire       [3:0]    _zz_cmdLogic_incrLen_2;
  wire       [4:0]    _zz_dataLogic_byteCounterNext;
  wire       [7:0]    _zz_dataLogic_byteCounterNext_1;
  reg        [15:0]   _zz_dataLogic_byteActivity;
  wire       [1:0]    _zz_dataLogic_byteActivity_1;
  wire                cmdLogic_outputFork_valid;
  wire                cmdLogic_outputFork_ready;
  wire       [31:0]   cmdLogic_outputFork_payload_addr;
  wire       [3:0]    cmdLogic_outputFork_payload_id;
  wire       [3:0]    cmdLogic_outputFork_payload_region;
  wire       [7:0]    cmdLogic_outputFork_payload_len;
  wire       [2:0]    cmdLogic_outputFork_payload_size;
  wire       [1:0]    cmdLogic_outputFork_payload_burst;
  wire       [0:0]    cmdLogic_outputFork_payload_lock;
  wire       [3:0]    cmdLogic_outputFork_payload_cache;
  wire       [3:0]    cmdLogic_outputFork_payload_qos;
  wire       [2:0]    cmdLogic_outputFork_payload_prot;
  wire                cmdLogic_dataFork_valid;
  wire                cmdLogic_dataFork_ready;
  wire       [31:0]   cmdLogic_dataFork_payload_addr;
  wire       [3:0]    cmdLogic_dataFork_payload_id;
  wire       [3:0]    cmdLogic_dataFork_payload_region;
  wire       [7:0]    cmdLogic_dataFork_payload_len;
  wire       [2:0]    cmdLogic_dataFork_payload_size;
  wire       [1:0]    cmdLogic_dataFork_payload_burst;
  wire       [0:0]    cmdLogic_dataFork_payload_lock;
  wire       [3:0]    cmdLogic_dataFork_payload_cache;
  wire       [3:0]    cmdLogic_dataFork_payload_qos;
  wire       [2:0]    cmdLogic_dataFork_payload_prot;
  reg                 io_input_aw_fork2_logic_linkEnable_0;
  reg                 io_input_aw_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdLogic_outputFork_fire;
  wire                cmdLogic_dataFork_fire;
  wire       [10:0]   cmdLogic_byteCount;
  wire       [7:0]    cmdLogic_incrLen;
  wire                when_Axi4Upsizer_l21;
  wire                when_Axi4Upsizer_l24;
  reg        [3:0]    dataLogic_byteCounter;
  reg        [2:0]    dataLogic_size;
  reg                 dataLogic_outputValid;
  reg                 dataLogic_outputLast;
  reg                 dataLogic_busy;
  reg                 dataLogic_incrementByteCounter;
  reg                 dataLogic_alwaysFire;
  wire       [4:0]    dataLogic_byteCounterNext;
  reg        [127:0]  dataLogic_dataBuffer;
  reg        [15:0]   dataLogic_maskBuffer;
  wire       [15:0]   dataLogic_byteActivity;
  wire                io_output_w_fire;
  wire                io_output_w_isStall;
  wire                io_input_w_fire;
  wire                when_Axi4Upsizer_l59;
  wire                when_Axi4Upsizer_l59_1;
  wire                when_Axi4Upsizer_l59_2;
  wire                when_Axi4Upsizer_l59_3;
  wire                when_Axi4Upsizer_l59_4;
  wire                when_Axi4Upsizer_l59_5;
  wire                when_Axi4Upsizer_l59_6;
  wire                when_Axi4Upsizer_l59_7;
  wire                when_Axi4Upsizer_l59_8;
  wire                when_Axi4Upsizer_l59_9;
  wire                when_Axi4Upsizer_l59_10;
  wire                when_Axi4Upsizer_l59_11;
  wire                when_Axi4Upsizer_l59_12;
  wire                when_Axi4Upsizer_l59_13;
  wire                when_Axi4Upsizer_l59_14;
  wire                when_Axi4Upsizer_l59_15;
  wire                when_Axi4Upsizer_l68;
  wire                when_Axi4Upsizer_l68_1;
  wire                when_Axi4Upsizer_l68_2;
  wire                when_Axi4Upsizer_l68_3;

  assign _zz_cmdLogic_byteCount = ({7'd0,io_input_aw_payload_len} <<< io_input_aw_payload_size);
  assign _zz_cmdLogic_incrLen = ({1'b0,cmdLogic_byteCount} + _zz_cmdLogic_incrLen_1);
  assign _zz_cmdLogic_incrLen_2 = io_input_aw_payload_addr[3 : 0];
  assign _zz_cmdLogic_incrLen_1 = {8'd0, _zz_cmdLogic_incrLen_2};
  assign _zz_dataLogic_byteCounterNext_1 = ({7'd0,1'b1} <<< dataLogic_size);
  assign _zz_dataLogic_byteCounterNext = _zz_dataLogic_byteCounterNext_1[4:0];
  assign _zz_dataLogic_byteActivity_1 = dataLogic_size[1:0];
  always @(*) begin
    case(_zz_dataLogic_byteActivity_1)
      2'b00 : _zz_dataLogic_byteActivity = 16'h0001;
      2'b01 : _zz_dataLogic_byteActivity = 16'h0003;
      2'b10 : _zz_dataLogic_byteActivity = 16'h000f;
      default : _zz_dataLogic_byteActivity = 16'h00ff;
    endcase
  end

  always @(*) begin
    io_input_aw_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_input_aw_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_input_aw_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdLogic_outputFork_ready) && io_input_aw_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdLogic_dataFork_ready) && io_input_aw_fork2_logic_linkEnable_1);
  assign cmdLogic_outputFork_valid = (io_input_aw_valid && io_input_aw_fork2_logic_linkEnable_0);
  assign cmdLogic_outputFork_payload_addr = io_input_aw_payload_addr;
  assign cmdLogic_outputFork_payload_id = io_input_aw_payload_id;
  assign cmdLogic_outputFork_payload_region = io_input_aw_payload_region;
  assign cmdLogic_outputFork_payload_len = io_input_aw_payload_len;
  assign cmdLogic_outputFork_payload_size = io_input_aw_payload_size;
  assign cmdLogic_outputFork_payload_burst = io_input_aw_payload_burst;
  assign cmdLogic_outputFork_payload_lock = io_input_aw_payload_lock;
  assign cmdLogic_outputFork_payload_cache = io_input_aw_payload_cache;
  assign cmdLogic_outputFork_payload_qos = io_input_aw_payload_qos;
  assign cmdLogic_outputFork_payload_prot = io_input_aw_payload_prot;
  assign cmdLogic_outputFork_fire = (cmdLogic_outputFork_valid && cmdLogic_outputFork_ready);
  assign cmdLogic_dataFork_valid = (io_input_aw_valid && io_input_aw_fork2_logic_linkEnable_1);
  assign cmdLogic_dataFork_payload_addr = io_input_aw_payload_addr;
  assign cmdLogic_dataFork_payload_id = io_input_aw_payload_id;
  assign cmdLogic_dataFork_payload_region = io_input_aw_payload_region;
  assign cmdLogic_dataFork_payload_len = io_input_aw_payload_len;
  assign cmdLogic_dataFork_payload_size = io_input_aw_payload_size;
  assign cmdLogic_dataFork_payload_burst = io_input_aw_payload_burst;
  assign cmdLogic_dataFork_payload_lock = io_input_aw_payload_lock;
  assign cmdLogic_dataFork_payload_cache = io_input_aw_payload_cache;
  assign cmdLogic_dataFork_payload_qos = io_input_aw_payload_qos;
  assign cmdLogic_dataFork_payload_prot = io_input_aw_payload_prot;
  assign cmdLogic_dataFork_fire = (cmdLogic_dataFork_valid && cmdLogic_dataFork_ready);
  assign io_output_aw_valid = cmdLogic_outputFork_valid;
  assign cmdLogic_outputFork_ready = io_output_aw_ready;
  assign io_output_aw_payload_addr = cmdLogic_outputFork_payload_addr;
  assign io_output_aw_payload_id = cmdLogic_outputFork_payload_id;
  assign io_output_aw_payload_region = cmdLogic_outputFork_payload_region;
  always @(*) begin
    io_output_aw_payload_len = cmdLogic_outputFork_payload_len;
    if(when_Axi4Upsizer_l21) begin
      io_output_aw_payload_len = cmdLogic_incrLen;
    end
  end

  always @(*) begin
    io_output_aw_payload_size = cmdLogic_outputFork_payload_size;
    if(when_Axi4Upsizer_l21) begin
      io_output_aw_payload_size = 3'b100;
      if(when_Axi4Upsizer_l24) begin
        io_output_aw_payload_size = io_input_aw_payload_size;
      end
    end
  end

  assign io_output_aw_payload_burst = cmdLogic_outputFork_payload_burst;
  assign io_output_aw_payload_lock = cmdLogic_outputFork_payload_lock;
  assign io_output_aw_payload_cache = cmdLogic_outputFork_payload_cache;
  assign io_output_aw_payload_qos = cmdLogic_outputFork_payload_qos;
  assign io_output_aw_payload_prot = cmdLogic_outputFork_payload_prot;
  assign cmdLogic_byteCount = _zz_cmdLogic_byteCount[10:0];
  assign cmdLogic_incrLen = _zz_cmdLogic_incrLen[11 : 4];
  assign when_Axi4Upsizer_l21 = (io_output_aw_payload_burst == 2'b01);
  assign when_Axi4Upsizer_l24 = (io_input_aw_payload_len == 8'h0);
  assign dataLogic_byteCounterNext = ({1'b0,dataLogic_byteCounter} + _zz_dataLogic_byteCounterNext);
  assign dataLogic_byteActivity = (_zz_dataLogic_byteActivity <<< dataLogic_byteCounter);
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign io_output_w_valid = dataLogic_outputValid;
  assign io_output_w_isStall = (io_output_w_valid && (! io_output_w_ready));
  assign io_input_w_ready = (dataLogic_busy && (! io_output_w_isStall));
  assign io_output_w_payload_data = dataLogic_dataBuffer;
  assign io_output_w_payload_strb = dataLogic_maskBuffer;
  assign io_output_w_payload_last = dataLogic_outputLast;
  assign io_input_w_fire = (io_input_w_valid && io_input_w_ready);
  assign when_Axi4Upsizer_l59 = dataLogic_byteActivity[0];
  assign when_Axi4Upsizer_l59_1 = dataLogic_byteActivity[1];
  assign when_Axi4Upsizer_l59_2 = dataLogic_byteActivity[2];
  assign when_Axi4Upsizer_l59_3 = dataLogic_byteActivity[3];
  assign when_Axi4Upsizer_l59_4 = dataLogic_byteActivity[4];
  assign when_Axi4Upsizer_l59_5 = dataLogic_byteActivity[5];
  assign when_Axi4Upsizer_l59_6 = dataLogic_byteActivity[6];
  assign when_Axi4Upsizer_l59_7 = dataLogic_byteActivity[7];
  assign when_Axi4Upsizer_l59_8 = dataLogic_byteActivity[8];
  assign when_Axi4Upsizer_l59_9 = dataLogic_byteActivity[9];
  assign when_Axi4Upsizer_l59_10 = dataLogic_byteActivity[10];
  assign when_Axi4Upsizer_l59_11 = dataLogic_byteActivity[11];
  assign when_Axi4Upsizer_l59_12 = dataLogic_byteActivity[12];
  assign when_Axi4Upsizer_l59_13 = dataLogic_byteActivity[13];
  assign when_Axi4Upsizer_l59_14 = dataLogic_byteActivity[14];
  assign when_Axi4Upsizer_l59_15 = dataLogic_byteActivity[15];
  assign when_Axi4Upsizer_l68 = (3'b000 < cmdLogic_dataFork_payload_size);
  assign when_Axi4Upsizer_l68_1 = (3'b001 < cmdLogic_dataFork_payload_size);
  assign when_Axi4Upsizer_l68_2 = (3'b010 < cmdLogic_dataFork_payload_size);
  assign when_Axi4Upsizer_l68_3 = (3'b011 < cmdLogic_dataFork_payload_size);
  assign cmdLogic_dataFork_ready = (! dataLogic_busy);
  assign io_input_b_valid = io_output_b_valid;
  assign io_output_b_ready = io_input_b_ready;
  assign io_input_b_payload_id = io_output_b_payload_id;
  assign io_input_b_payload_resp = io_output_b_payload_resp;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      io_input_aw_fork2_logic_linkEnable_0 <= 1'b1;
      io_input_aw_fork2_logic_linkEnable_1 <= 1'b1;
      dataLogic_outputValid <= 1'b0;
      dataLogic_busy <= 1'b0;
      dataLogic_maskBuffer <= 16'h0;
    end else begin
      if(cmdLogic_outputFork_fire) begin
        io_input_aw_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdLogic_dataFork_fire) begin
        io_input_aw_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_aw_ready) begin
        io_input_aw_fork2_logic_linkEnable_0 <= 1'b1;
        io_input_aw_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(io_output_w_ready) begin
        dataLogic_outputValid <= 1'b0;
      end
      if(io_output_w_fire) begin
        dataLogic_maskBuffer <= 16'h0;
      end
      if(io_input_w_fire) begin
        dataLogic_outputValid <= ((dataLogic_byteCounterNext[4] || io_input_w_payload_last) || dataLogic_alwaysFire);
        if(io_input_w_payload_last) begin
          dataLogic_busy <= 1'b0;
        end
        if(when_Axi4Upsizer_l59) begin
          dataLogic_maskBuffer[0] <= io_input_w_payload_strb[0];
        end
        if(when_Axi4Upsizer_l59_1) begin
          dataLogic_maskBuffer[1] <= io_input_w_payload_strb[1];
        end
        if(when_Axi4Upsizer_l59_2) begin
          dataLogic_maskBuffer[2] <= io_input_w_payload_strb[2];
        end
        if(when_Axi4Upsizer_l59_3) begin
          dataLogic_maskBuffer[3] <= io_input_w_payload_strb[3];
        end
        if(when_Axi4Upsizer_l59_4) begin
          dataLogic_maskBuffer[4] <= io_input_w_payload_strb[4];
        end
        if(when_Axi4Upsizer_l59_5) begin
          dataLogic_maskBuffer[5] <= io_input_w_payload_strb[5];
        end
        if(when_Axi4Upsizer_l59_6) begin
          dataLogic_maskBuffer[6] <= io_input_w_payload_strb[6];
        end
        if(when_Axi4Upsizer_l59_7) begin
          dataLogic_maskBuffer[7] <= io_input_w_payload_strb[7];
        end
        if(when_Axi4Upsizer_l59_8) begin
          dataLogic_maskBuffer[8] <= io_input_w_payload_strb[0];
        end
        if(when_Axi4Upsizer_l59_9) begin
          dataLogic_maskBuffer[9] <= io_input_w_payload_strb[1];
        end
        if(when_Axi4Upsizer_l59_10) begin
          dataLogic_maskBuffer[10] <= io_input_w_payload_strb[2];
        end
        if(when_Axi4Upsizer_l59_11) begin
          dataLogic_maskBuffer[11] <= io_input_w_payload_strb[3];
        end
        if(when_Axi4Upsizer_l59_12) begin
          dataLogic_maskBuffer[12] <= io_input_w_payload_strb[4];
        end
        if(when_Axi4Upsizer_l59_13) begin
          dataLogic_maskBuffer[13] <= io_input_w_payload_strb[5];
        end
        if(when_Axi4Upsizer_l59_14) begin
          dataLogic_maskBuffer[14] <= io_input_w_payload_strb[6];
        end
        if(when_Axi4Upsizer_l59_15) begin
          dataLogic_maskBuffer[15] <= io_input_w_payload_strb[7];
        end
      end
      if(cmdLogic_dataFork_fire) begin
        dataLogic_busy <= 1'b1;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(io_input_w_fire) begin
      if(dataLogic_incrementByteCounter) begin
        dataLogic_byteCounter <= dataLogic_byteCounterNext[3:0];
      end
      dataLogic_outputLast <= io_input_w_payload_last;
      if(when_Axi4Upsizer_l59) begin
        dataLogic_dataBuffer[7 : 0] <= io_input_w_payload_data[7 : 0];
      end
      if(when_Axi4Upsizer_l59_1) begin
        dataLogic_dataBuffer[15 : 8] <= io_input_w_payload_data[15 : 8];
      end
      if(when_Axi4Upsizer_l59_2) begin
        dataLogic_dataBuffer[23 : 16] <= io_input_w_payload_data[23 : 16];
      end
      if(when_Axi4Upsizer_l59_3) begin
        dataLogic_dataBuffer[31 : 24] <= io_input_w_payload_data[31 : 24];
      end
      if(when_Axi4Upsizer_l59_4) begin
        dataLogic_dataBuffer[39 : 32] <= io_input_w_payload_data[39 : 32];
      end
      if(when_Axi4Upsizer_l59_5) begin
        dataLogic_dataBuffer[47 : 40] <= io_input_w_payload_data[47 : 40];
      end
      if(when_Axi4Upsizer_l59_6) begin
        dataLogic_dataBuffer[55 : 48] <= io_input_w_payload_data[55 : 48];
      end
      if(when_Axi4Upsizer_l59_7) begin
        dataLogic_dataBuffer[63 : 56] <= io_input_w_payload_data[63 : 56];
      end
      if(when_Axi4Upsizer_l59_8) begin
        dataLogic_dataBuffer[71 : 64] <= io_input_w_payload_data[7 : 0];
      end
      if(when_Axi4Upsizer_l59_9) begin
        dataLogic_dataBuffer[79 : 72] <= io_input_w_payload_data[15 : 8];
      end
      if(when_Axi4Upsizer_l59_10) begin
        dataLogic_dataBuffer[87 : 80] <= io_input_w_payload_data[23 : 16];
      end
      if(when_Axi4Upsizer_l59_11) begin
        dataLogic_dataBuffer[95 : 88] <= io_input_w_payload_data[31 : 24];
      end
      if(when_Axi4Upsizer_l59_12) begin
        dataLogic_dataBuffer[103 : 96] <= io_input_w_payload_data[39 : 32];
      end
      if(when_Axi4Upsizer_l59_13) begin
        dataLogic_dataBuffer[111 : 104] <= io_input_w_payload_data[47 : 40];
      end
      if(when_Axi4Upsizer_l59_14) begin
        dataLogic_dataBuffer[119 : 112] <= io_input_w_payload_data[55 : 48];
      end
      if(when_Axi4Upsizer_l59_15) begin
        dataLogic_dataBuffer[127 : 120] <= io_input_w_payload_data[63 : 56];
      end
    end
    if(cmdLogic_dataFork_fire) begin
      dataLogic_byteCounter <= cmdLogic_dataFork_payload_addr[3:0];
      if(when_Axi4Upsizer_l68) begin
        dataLogic_byteCounter[0] <= 1'b0;
      end
      if(when_Axi4Upsizer_l68_1) begin
        dataLogic_byteCounter[1] <= 1'b0;
      end
      if(when_Axi4Upsizer_l68_2) begin
        dataLogic_byteCounter[2] <= 1'b0;
      end
      if(when_Axi4Upsizer_l68_3) begin
        dataLogic_byteCounter[3] <= 1'b0;
      end
      dataLogic_size <= cmdLogic_dataFork_payload_size;
      dataLogic_alwaysFire <= (! (cmdLogic_dataFork_payload_burst == 2'b01));
      dataLogic_incrementByteCounter <= (! (cmdLogic_dataFork_payload_burst == 2'b00));
    end
  end


endmodule

module Axi4ReadOnlyUpsizer_1 (
  input  wire          io_input_ar_valid,
  output reg           io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [3:0]    io_input_ar_payload_region,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  input  wire [0:0]    io_input_ar_payload_lock,
  input  wire [3:0]    io_input_ar_payload_cache,
  input  wire [3:0]    io_input_ar_payload_qos,
  input  wire [2:0]    io_input_ar_payload_prot,
  output wire          io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [63:0]   io_input_r_payload_data,
  output wire [3:0]    io_input_r_payload_id,
  output wire [1:0]    io_input_r_payload_resp,
  output wire          io_input_r_payload_last,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [3:0]    io_output_ar_payload_id,
  output wire [3:0]    io_output_ar_payload_region,
  output wire [7:0]    io_output_ar_payload_len,
  output reg  [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  output wire [0:0]    io_output_ar_payload_lock,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [3:0]    io_output_ar_payload_qos,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [127:0]  io_output_r_payload_data,
  input  wire [3:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                dataLogic_cmdPush_fifo_io_pop_ready;
  wire                dataLogic_cmdPush_fifo_io_push_ready;
  wire                dataLogic_cmdPush_fifo_io_pop_valid;
  wire       [3:0]    dataLogic_cmdPush_fifo_io_pop_payload_startAt;
  wire       [3:0]    dataLogic_cmdPush_fifo_io_pop_payload_endAt;
  wire       [2:0]    dataLogic_cmdPush_fifo_io_pop_payload_size;
  wire       [3:0]    dataLogic_cmdPush_fifo_io_pop_payload_id;
  wire       [2:0]    dataLogic_cmdPush_fifo_io_occupancy;
  wire       [2:0]    dataLogic_cmdPush_fifo_io_availability;
  wire       [14:0]   _zz_cmdLogic_byteCount;
  wire       [11:0]   _zz_cmdLogic_incrLen;
  wire       [11:0]   _zz_cmdLogic_incrLen_1;
  wire       [3:0]    _zz_cmdLogic_incrLen_2;
  wire       [31:0]   _zz_dataLogic_cmdPush_payload_endAt;
  wire       [31:0]   _zz_dataLogic_cmdPush_payload_endAt_1;
  wire       [14:0]   _zz_dataLogic_cmdPush_payload_endAt_2;
  wire       [4:0]    _zz_dataLogic_byteCounterNext;
  wire       [7:0]    _zz_dataLogic_byteCounterNext_1;
  reg        [63:0]   _zz_io_input_r_payload_data;
  wire       [0:0]    _zz_io_input_r_payload_data_1;
  wire                cmdLogic_outputFork_valid;
  wire                cmdLogic_outputFork_ready;
  wire       [31:0]   cmdLogic_outputFork_payload_addr;
  wire       [3:0]    cmdLogic_outputFork_payload_id;
  wire       [3:0]    cmdLogic_outputFork_payload_region;
  wire       [7:0]    cmdLogic_outputFork_payload_len;
  wire       [2:0]    cmdLogic_outputFork_payload_size;
  wire       [1:0]    cmdLogic_outputFork_payload_burst;
  wire       [0:0]    cmdLogic_outputFork_payload_lock;
  wire       [3:0]    cmdLogic_outputFork_payload_cache;
  wire       [3:0]    cmdLogic_outputFork_payload_qos;
  wire       [2:0]    cmdLogic_outputFork_payload_prot;
  wire                cmdLogic_dataFork_valid;
  wire                cmdLogic_dataFork_ready;
  wire       [31:0]   cmdLogic_dataFork_payload_addr;
  wire       [3:0]    cmdLogic_dataFork_payload_id;
  wire       [3:0]    cmdLogic_dataFork_payload_region;
  wire       [7:0]    cmdLogic_dataFork_payload_len;
  wire       [2:0]    cmdLogic_dataFork_payload_size;
  wire       [1:0]    cmdLogic_dataFork_payload_burst;
  wire       [0:0]    cmdLogic_dataFork_payload_lock;
  wire       [3:0]    cmdLogic_dataFork_payload_cache;
  wire       [3:0]    cmdLogic_dataFork_payload_qos;
  wire       [2:0]    cmdLogic_dataFork_payload_prot;
  reg                 io_input_ar_fork2_logic_linkEnable_0;
  reg                 io_input_ar_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdLogic_outputFork_fire;
  wire                cmdLogic_dataFork_fire;
  wire       [10:0]   cmdLogic_byteCount;
  wire       [7:0]    cmdLogic_incrLen;
  wire                when_Axi4Upsizer_l108;
  wire                dataLogic_cmdPush_valid;
  wire                dataLogic_cmdPush_ready;
  wire       [3:0]    dataLogic_cmdPush_payload_startAt;
  wire       [3:0]    dataLogic_cmdPush_payload_endAt;
  wire       [2:0]    dataLogic_cmdPush_payload_size;
  wire       [3:0]    dataLogic_cmdPush_payload_id;
  reg        [2:0]    dataLogic_size;
  reg                 dataLogic_busy;
  reg        [3:0]    dataLogic_id;
  reg        [3:0]    dataLogic_byteCounter;
  reg        [3:0]    dataLogic_byteCounterLast;
  wire       [4:0]    dataLogic_byteCounterNext;
  wire                dataLogic_cmdPush_fifo_io_pop_fire;
  wire                io_input_r_fire;

  assign _zz_cmdLogic_byteCount = ({7'd0,io_input_ar_payload_len} <<< io_input_ar_payload_size);
  assign _zz_cmdLogic_incrLen = ({1'b0,cmdLogic_byteCount} + _zz_cmdLogic_incrLen_1);
  assign _zz_cmdLogic_incrLen_2 = io_input_ar_payload_addr[3 : 0];
  assign _zz_cmdLogic_incrLen_1 = {8'd0, _zz_cmdLogic_incrLen_2};
  assign _zz_dataLogic_cmdPush_payload_endAt = (cmdLogic_dataFork_payload_addr + _zz_dataLogic_cmdPush_payload_endAt_1);
  assign _zz_dataLogic_cmdPush_payload_endAt_2 = ({7'd0,cmdLogic_dataFork_payload_len} <<< cmdLogic_dataFork_payload_size);
  assign _zz_dataLogic_cmdPush_payload_endAt_1 = {17'd0, _zz_dataLogic_cmdPush_payload_endAt_2};
  assign _zz_dataLogic_byteCounterNext_1 = ({7'd0,1'b1} <<< dataLogic_size);
  assign _zz_dataLogic_byteCounterNext = _zz_dataLogic_byteCounterNext_1[4:0];
  assign _zz_io_input_r_payload_data_1 = (dataLogic_byteCounter >>> 2'd3);
  StreamFifo_4 dataLogic_cmdPush_fifo (
    .io_push_valid           (dataLogic_cmdPush_valid                           ), //i
    .io_push_ready           (dataLogic_cmdPush_fifo_io_push_ready              ), //o
    .io_push_payload_startAt (dataLogic_cmdPush_payload_startAt[3:0]            ), //i
    .io_push_payload_endAt   (dataLogic_cmdPush_payload_endAt[3:0]              ), //i
    .io_push_payload_size    (dataLogic_cmdPush_payload_size[2:0]               ), //i
    .io_push_payload_id      (dataLogic_cmdPush_payload_id[3:0]                 ), //i
    .io_pop_valid            (dataLogic_cmdPush_fifo_io_pop_valid               ), //o
    .io_pop_ready            (dataLogic_cmdPush_fifo_io_pop_ready               ), //i
    .io_pop_payload_startAt  (dataLogic_cmdPush_fifo_io_pop_payload_startAt[3:0]), //o
    .io_pop_payload_endAt    (dataLogic_cmdPush_fifo_io_pop_payload_endAt[3:0]  ), //o
    .io_pop_payload_size     (dataLogic_cmdPush_fifo_io_pop_payload_size[2:0]   ), //o
    .io_pop_payload_id       (dataLogic_cmdPush_fifo_io_pop_payload_id[3:0]     ), //o
    .io_flush                (1'b0                                              ), //i
    .io_occupancy            (dataLogic_cmdPush_fifo_io_occupancy[2:0]          ), //o
    .io_availability         (dataLogic_cmdPush_fifo_io_availability[2:0]       ), //o
    .io_memoryClk            (io_memoryClk                                      ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                           )  //i
  );
  always @(*) begin
    case(_zz_io_input_r_payload_data_1)
      1'b0 : _zz_io_input_r_payload_data = io_output_r_payload_data[63 : 0];
      default : _zz_io_input_r_payload_data = io_output_r_payload_data[127 : 64];
    endcase
  end

  always @(*) begin
    io_input_ar_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_input_ar_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_input_ar_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdLogic_outputFork_ready) && io_input_ar_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdLogic_dataFork_ready) && io_input_ar_fork2_logic_linkEnable_1);
  assign cmdLogic_outputFork_valid = (io_input_ar_valid && io_input_ar_fork2_logic_linkEnable_0);
  assign cmdLogic_outputFork_payload_addr = io_input_ar_payload_addr;
  assign cmdLogic_outputFork_payload_id = io_input_ar_payload_id;
  assign cmdLogic_outputFork_payload_region = io_input_ar_payload_region;
  assign cmdLogic_outputFork_payload_len = io_input_ar_payload_len;
  assign cmdLogic_outputFork_payload_size = io_input_ar_payload_size;
  assign cmdLogic_outputFork_payload_burst = io_input_ar_payload_burst;
  assign cmdLogic_outputFork_payload_lock = io_input_ar_payload_lock;
  assign cmdLogic_outputFork_payload_cache = io_input_ar_payload_cache;
  assign cmdLogic_outputFork_payload_qos = io_input_ar_payload_qos;
  assign cmdLogic_outputFork_payload_prot = io_input_ar_payload_prot;
  assign cmdLogic_outputFork_fire = (cmdLogic_outputFork_valid && cmdLogic_outputFork_ready);
  assign cmdLogic_dataFork_valid = (io_input_ar_valid && io_input_ar_fork2_logic_linkEnable_1);
  assign cmdLogic_dataFork_payload_addr = io_input_ar_payload_addr;
  assign cmdLogic_dataFork_payload_id = io_input_ar_payload_id;
  assign cmdLogic_dataFork_payload_region = io_input_ar_payload_region;
  assign cmdLogic_dataFork_payload_len = io_input_ar_payload_len;
  assign cmdLogic_dataFork_payload_size = io_input_ar_payload_size;
  assign cmdLogic_dataFork_payload_burst = io_input_ar_payload_burst;
  assign cmdLogic_dataFork_payload_lock = io_input_ar_payload_lock;
  assign cmdLogic_dataFork_payload_cache = io_input_ar_payload_cache;
  assign cmdLogic_dataFork_payload_qos = io_input_ar_payload_qos;
  assign cmdLogic_dataFork_payload_prot = io_input_ar_payload_prot;
  assign cmdLogic_dataFork_fire = (cmdLogic_dataFork_valid && cmdLogic_dataFork_ready);
  assign io_output_ar_valid = cmdLogic_outputFork_valid;
  assign cmdLogic_outputFork_ready = io_output_ar_ready;
  assign io_output_ar_payload_addr = cmdLogic_outputFork_payload_addr;
  assign io_output_ar_payload_region = cmdLogic_outputFork_payload_region;
  assign io_output_ar_payload_burst = cmdLogic_outputFork_payload_burst;
  assign io_output_ar_payload_lock = cmdLogic_outputFork_payload_lock;
  assign io_output_ar_payload_cache = cmdLogic_outputFork_payload_cache;
  assign io_output_ar_payload_qos = cmdLogic_outputFork_payload_qos;
  assign io_output_ar_payload_prot = cmdLogic_outputFork_payload_prot;
  assign cmdLogic_byteCount = _zz_cmdLogic_byteCount[10:0];
  assign cmdLogic_incrLen = _zz_cmdLogic_incrLen[11 : 4];
  always @(*) begin
    io_output_ar_payload_size = 3'b100;
    if(when_Axi4Upsizer_l108) begin
      io_output_ar_payload_size = io_input_ar_payload_size;
    end
  end

  assign io_output_ar_payload_len = cmdLogic_incrLen;
  assign io_output_ar_payload_id = 4'b0000;
  assign when_Axi4Upsizer_l108 = (io_input_ar_payload_len == 8'h0);
  assign dataLogic_cmdPush_valid = cmdLogic_dataFork_valid;
  assign cmdLogic_dataFork_ready = dataLogic_cmdPush_ready;
  assign dataLogic_cmdPush_payload_startAt = cmdLogic_dataFork_payload_addr[3:0];
  assign dataLogic_cmdPush_payload_endAt = _zz_dataLogic_cmdPush_payload_endAt[3:0];
  assign dataLogic_cmdPush_payload_size = cmdLogic_dataFork_payload_size;
  assign dataLogic_cmdPush_payload_id = cmdLogic_dataFork_payload_id;
  assign dataLogic_cmdPush_ready = dataLogic_cmdPush_fifo_io_push_ready;
  assign dataLogic_byteCounterNext = ({1'b0,dataLogic_byteCounter} + _zz_dataLogic_byteCounterNext);
  assign dataLogic_cmdPush_fifo_io_pop_fire = (dataLogic_cmdPush_fifo_io_pop_valid && dataLogic_cmdPush_fifo_io_pop_ready);
  assign dataLogic_cmdPush_fifo_io_pop_ready = (! dataLogic_busy);
  assign io_input_r_fire = (io_input_r_valid && io_input_r_ready);
  assign io_input_r_valid = (io_output_r_valid && dataLogic_busy);
  assign io_input_r_payload_last = (io_output_r_payload_last && (dataLogic_byteCounter == dataLogic_byteCounterLast));
  assign io_input_r_payload_resp = io_output_r_payload_resp;
  assign io_input_r_payload_data = _zz_io_input_r_payload_data;
  assign io_input_r_payload_id = dataLogic_id;
  assign io_output_r_ready = ((dataLogic_busy && io_input_r_ready) && (io_input_r_payload_last || dataLogic_byteCounterNext[4]));
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      io_input_ar_fork2_logic_linkEnable_0 <= 1'b1;
      io_input_ar_fork2_logic_linkEnable_1 <= 1'b1;
      dataLogic_busy <= 1'b0;
    end else begin
      if(cmdLogic_outputFork_fire) begin
        io_input_ar_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdLogic_dataFork_fire) begin
        io_input_ar_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_ar_ready) begin
        io_input_ar_fork2_logic_linkEnable_0 <= 1'b1;
        io_input_ar_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(dataLogic_cmdPush_fifo_io_pop_fire) begin
        dataLogic_busy <= 1'b1;
      end
      if(io_input_r_fire) begin
        if(io_input_r_payload_last) begin
          dataLogic_busy <= 1'b0;
        end
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(dataLogic_cmdPush_fifo_io_pop_fire) begin
      dataLogic_byteCounter <= dataLogic_cmdPush_fifo_io_pop_payload_startAt;
      dataLogic_byteCounterLast <= dataLogic_cmdPush_fifo_io_pop_payload_endAt;
      dataLogic_size <= dataLogic_cmdPush_fifo_io_pop_payload_size;
      dataLogic_id <= dataLogic_cmdPush_fifo_io_pop_payload_id;
    end
    if(io_input_r_fire) begin
      dataLogic_byteCounter <= dataLogic_byteCounterNext[3:0];
    end
  end


endmodule

module StreamFifoCC_11 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [3:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [3:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset,
  input  wire          io_ddrMasters_0_clk,
  input  wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1
);

  reg        [5:0]    ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [5:0]    _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [1:0]    popCC_readPort_rsp_resp;
  wire       [5:0]    _zz_popCC_readPort_rsp_id;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [1:0]    popCC_readArbitation_translated_payload_resp;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [5:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_resp,io_push_payload_id};
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_14 popToPushGray_buffercc (
    .io_dataIn               (popToPushGray[4:0]                    ), //i
    .io_dataOut              (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_memoryClk            (io_memoryClk                          ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_34 pushToPopGray_buffercc (
    .io_dataIn                                                                                 (pushToPopGray[4:0]                                                                       ), //i
    .io_dataOut                                                                                (pushToPopGray_buffercc_io_dataOut[4:0]                                                   ), //o
    .io_ddrMasters_0_clk                                                                       (io_ddrMasters_0_clk                                                                      ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_id = ram_spinal_port1;
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_id[3 : 0];
  assign popCC_readPort_rsp_resp = _zz_popCC_readPort_rsp_id[5 : 4];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_resp = popCC_readPort_rsp_resp;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = popCC_readArbitation_translated_payload_resp;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_10 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [63:0]   io_push_payload_data,
  input  wire [7:0]    io_push_payload_strb,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [63:0]   io_pop_payload_data,
  output wire [7:0]    io_pop_payload_strb,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_ddrMasters_0_clk,
  input  wire          io_ddrMasters_0_reset,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1
);

  reg        [72:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [72:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [63:0]   popCC_readPort_rsp_data;
  wire       [7:0]    popCC_readPort_rsp_strb;
  wire                popCC_readPort_rsp_last;
  wire       [72:0]   _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [63:0]   popCC_readArbitation_translated_payload_data;
  wire       [7:0]    popCC_readArbitation_translated_payload_strb;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [72:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_strb,io_push_payload_data}};
  always @(posedge io_ddrMasters_0_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_23 popToPushGray_buffercc (
    .io_dataIn             (popToPushGray[4:0]                    ), //i
    .io_dataOut            (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_ddrMasters_0_clk   (io_ddrMasters_0_clk                   ), //i
    .io_ddrMasters_0_reset (io_ddrMasters_0_reset                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_30 pushToPopGray_buffercc (
    .io_dataIn                                                                               (pushToPopGray[4:0]                                                                     ), //i
    .io_dataOut                                                                              (pushToPopGray_buffercc_io_dataOut[4:0]                                                 ), //o
    .io_memoryClk                                                                            (io_memoryClk                                                                           ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1 (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[63 : 0];
  assign popCC_readPort_rsp_strb = _zz_popCC_readPort_rsp_data[71 : 64];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[72];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_strb = popCC_readPort_rsp_strb;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_strb = popCC_readArbitation_translated_payload_strb;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_ddrMasters_0_clk) begin
    if(io_ddrMasters_0_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_9 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_addr,
  input  wire [3:0]    io_push_payload_id,
  input  wire [3:0]    io_push_payload_region,
  input  wire [7:0]    io_push_payload_len,
  input  wire [2:0]    io_push_payload_size,
  input  wire [1:0]    io_push_payload_burst,
  input  wire [0:0]    io_push_payload_lock,
  input  wire [3:0]    io_push_payload_cache,
  input  wire [3:0]    io_push_payload_qos,
  input  wire [2:0]    io_push_payload_prot,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_addr,
  output wire [3:0]    io_pop_payload_id,
  output wire [3:0]    io_pop_payload_region,
  output wire [7:0]    io_pop_payload_len,
  output wire [2:0]    io_pop_payload_size,
  output wire [1:0]    io_pop_payload_burst,
  output wire [0:0]    io_pop_payload_lock,
  output wire [3:0]    io_pop_payload_cache,
  output wire [3:0]    io_pop_payload_qos,
  output wire [2:0]    io_pop_payload_prot,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_ddrMasters_0_clk,
  input  wire          io_ddrMasters_0_reset,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1
);

  reg        [64:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [64:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [31:0]   popCC_readPort_rsp_addr;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [3:0]    popCC_readPort_rsp_region;
  wire       [7:0]    popCC_readPort_rsp_len;
  wire       [2:0]    popCC_readPort_rsp_size;
  wire       [1:0]    popCC_readPort_rsp_burst;
  wire       [0:0]    popCC_readPort_rsp_lock;
  wire       [3:0]    popCC_readPort_rsp_cache;
  wire       [3:0]    popCC_readPort_rsp_qos;
  wire       [2:0]    popCC_readPort_rsp_prot;
  wire       [64:0]   _zz_popCC_readPort_rsp_addr;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [31:0]   popCC_readArbitation_translated_payload_addr;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [3:0]    popCC_readArbitation_translated_payload_region;
  wire       [7:0]    popCC_readArbitation_translated_payload_len;
  wire       [2:0]    popCC_readArbitation_translated_payload_size;
  wire       [1:0]    popCC_readArbitation_translated_payload_burst;
  wire       [0:0]    popCC_readArbitation_translated_payload_lock;
  wire       [3:0]    popCC_readArbitation_translated_payload_cache;
  wire       [3:0]    popCC_readArbitation_translated_payload_qos;
  wire       [2:0]    popCC_readArbitation_translated_payload_prot;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [64:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_prot,{io_push_payload_qos,{io_push_payload_cache,{io_push_payload_lock,{io_push_payload_burst,{io_push_payload_size,{io_push_payload_len,{io_push_payload_region,{io_push_payload_id,io_push_payload_addr}}}}}}}}};
  always @(posedge io_ddrMasters_0_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_23 popToPushGray_buffercc (
    .io_dataIn             (popToPushGray[4:0]                    ), //i
    .io_dataOut            (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_ddrMasters_0_clk   (io_ddrMasters_0_clk                   ), //i
    .io_ddrMasters_0_reset (io_ddrMasters_0_reset                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_30 pushToPopGray_buffercc (
    .io_dataIn                                                                               (pushToPopGray[4:0]                                                                     ), //i
    .io_dataOut                                                                              (pushToPopGray_buffercc_io_dataOut[4:0]                                                 ), //o
    .io_memoryClk                                                                            (io_memoryClk                                                                           ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1 (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_addr = ram_spinal_port1;
  assign popCC_readPort_rsp_addr = _zz_popCC_readPort_rsp_addr[31 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_addr[35 : 32];
  assign popCC_readPort_rsp_region = _zz_popCC_readPort_rsp_addr[39 : 36];
  assign popCC_readPort_rsp_len = _zz_popCC_readPort_rsp_addr[47 : 40];
  assign popCC_readPort_rsp_size = _zz_popCC_readPort_rsp_addr[50 : 48];
  assign popCC_readPort_rsp_burst = _zz_popCC_readPort_rsp_addr[52 : 51];
  assign popCC_readPort_rsp_lock = _zz_popCC_readPort_rsp_addr[53 : 53];
  assign popCC_readPort_rsp_cache = _zz_popCC_readPort_rsp_addr[57 : 54];
  assign popCC_readPort_rsp_qos = _zz_popCC_readPort_rsp_addr[61 : 58];
  assign popCC_readPort_rsp_prot = _zz_popCC_readPort_rsp_addr[64 : 62];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_addr = popCC_readPort_rsp_addr;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_region = popCC_readPort_rsp_region;
  assign popCC_readArbitation_translated_payload_len = popCC_readPort_rsp_len;
  assign popCC_readArbitation_translated_payload_size = popCC_readPort_rsp_size;
  assign popCC_readArbitation_translated_payload_burst = popCC_readPort_rsp_burst;
  assign popCC_readArbitation_translated_payload_lock = popCC_readPort_rsp_lock;
  assign popCC_readArbitation_translated_payload_cache = popCC_readPort_rsp_cache;
  assign popCC_readArbitation_translated_payload_qos = popCC_readPort_rsp_qos;
  assign popCC_readArbitation_translated_payload_prot = popCC_readPort_rsp_prot;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_addr = popCC_readArbitation_translated_payload_addr;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_region = popCC_readArbitation_translated_payload_region;
  assign io_pop_payload_len = popCC_readArbitation_translated_payload_len;
  assign io_pop_payload_size = popCC_readArbitation_translated_payload_size;
  assign io_pop_payload_burst = popCC_readArbitation_translated_payload_burst;
  assign io_pop_payload_lock = popCC_readArbitation_translated_payload_lock;
  assign io_pop_payload_cache = popCC_readArbitation_translated_payload_cache;
  assign io_pop_payload_qos = popCC_readArbitation_translated_payload_qos;
  assign io_pop_payload_prot = popCC_readArbitation_translated_payload_prot;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_ddrMasters_0_clk) begin
    if(io_ddrMasters_0_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_8 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [63:0]   io_push_payload_data,
  input  wire [3:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [63:0]   io_pop_payload_data,
  output wire [3:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset,
  input  wire          io_ddrMasters_0_clk,
  output wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1
);

  reg        [70:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [70:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [63:0]   popCC_readPort_rsp_data;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [1:0]    popCC_readPort_rsp_resp;
  wire                popCC_readPort_rsp_last;
  wire       [70:0]   _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [63:0]   popCC_readArbitation_translated_payload_data;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [1:0]    popCC_readArbitation_translated_payload_resp;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [70:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_resp,{io_push_payload_id,io_push_payload_data}}};
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_14 popToPushGray_buffercc (
    .io_dataIn               (popToPushGray[4:0]                    ), //i
    .io_dataOut              (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_memoryClk            (io_memoryClk                          ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_27 system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn               (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut              (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_ddrMasters_0_clk     (io_ddrMasters_0_clk                                                                                                   ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                                                                                               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_28 pushToPopGray_buffercc (
    .io_dataIn                                                                               (pushToPopGray[4:0]                                                                     ), //i
    .io_dataOut                                                                              (pushToPopGray_buffercc_io_dataOut[4:0]                                                 ), //o
    .io_ddrMasters_0_clk                                                                     (io_ddrMasters_0_clk                                                                    ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized = system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[63 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_data[67 : 64];
  assign popCC_readPort_rsp_resp = _zz_popCC_readPort_rsp_data[69 : 68];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[70];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_resp = popCC_readPort_rsp_resp;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = popCC_readArbitation_translated_payload_resp;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 = system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_ddrMasters_0_clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_7 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_addr,
  input  wire [3:0]    io_push_payload_id,
  input  wire [3:0]    io_push_payload_region,
  input  wire [7:0]    io_push_payload_len,
  input  wire [2:0]    io_push_payload_size,
  input  wire [1:0]    io_push_payload_burst,
  input  wire [0:0]    io_push_payload_lock,
  input  wire [3:0]    io_push_payload_cache,
  input  wire [3:0]    io_push_payload_qos,
  input  wire [2:0]    io_push_payload_prot,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_addr,
  output wire [3:0]    io_pop_payload_id,
  output wire [3:0]    io_pop_payload_region,
  output wire [7:0]    io_pop_payload_len,
  output wire [2:0]    io_pop_payload_size,
  output wire [1:0]    io_pop_payload_burst,
  output wire [0:0]    io_pop_payload_lock,
  output wire [3:0]    io_pop_payload_cache,
  output wire [3:0]    io_pop_payload_qos,
  output wire [2:0]    io_pop_payload_prot,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_ddrMasters_0_clk,
  input  wire          io_ddrMasters_0_reset,
  input  wire          io_memoryClk,
  output wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1
);

  reg        [64:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [64:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_asyncAssertSyncDeassert;
  wire                system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [31:0]   popCC_readPort_rsp_addr;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [3:0]    popCC_readPort_rsp_region;
  wire       [7:0]    popCC_readPort_rsp_len;
  wire       [2:0]    popCC_readPort_rsp_size;
  wire       [1:0]    popCC_readPort_rsp_burst;
  wire       [0:0]    popCC_readPort_rsp_lock;
  wire       [3:0]    popCC_readPort_rsp_cache;
  wire       [3:0]    popCC_readPort_rsp_qos;
  wire       [2:0]    popCC_readPort_rsp_prot;
  wire       [64:0]   _zz_popCC_readPort_rsp_addr;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [31:0]   popCC_readArbitation_translated_payload_addr;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [3:0]    popCC_readArbitation_translated_payload_region;
  wire       [7:0]    popCC_readArbitation_translated_payload_len;
  wire       [2:0]    popCC_readArbitation_translated_payload_size;
  wire       [1:0]    popCC_readArbitation_translated_payload_burst;
  wire       [0:0]    popCC_readArbitation_translated_payload_lock;
  wire       [3:0]    popCC_readArbitation_translated_payload_cache;
  wire       [3:0]    popCC_readArbitation_translated_payload_qos;
  wire       [2:0]    popCC_readArbitation_translated_payload_prot;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [64:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_prot,{io_push_payload_qos,{io_push_payload_cache,{io_push_payload_lock,{io_push_payload_burst,{io_push_payload_size,{io_push_payload_len,{io_push_payload_region,{io_push_payload_id,io_push_payload_addr}}}}}}}}};
  always @(posedge io_ddrMasters_0_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_23 popToPushGray_buffercc (
    .io_dataIn             (popToPushGray[4:0]                    ), //i
    .io_dataOut            (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_ddrMasters_0_clk   (io_ddrMasters_0_clk                   ), //i
    .io_ddrMasters_0_reset (io_ddrMasters_0_reset                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_24 system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn             (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut            (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_memoryClk          (io_memoryClk                                                                                                        ), //i
    .io_ddrMasters_0_reset (io_ddrMasters_0_reset                                                                                               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_25 pushToPopGray_buffercc (
    .io_dataIn                                                                             (pushToPopGray[4:0]                                                                   ), //i
    .io_dataOut                                                                            (pushToPopGray_buffercc_io_dataOut[4:0]                                               ), //o
    .io_memoryClk                                                                          (io_memoryClk                                                                         ), //i
    .system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized (system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized = system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_addr = ram_spinal_port1;
  assign popCC_readPort_rsp_addr = _zz_popCC_readPort_rsp_addr[31 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_addr[35 : 32];
  assign popCC_readPort_rsp_region = _zz_popCC_readPort_rsp_addr[39 : 36];
  assign popCC_readPort_rsp_len = _zz_popCC_readPort_rsp_addr[47 : 40];
  assign popCC_readPort_rsp_size = _zz_popCC_readPort_rsp_addr[50 : 48];
  assign popCC_readPort_rsp_burst = _zz_popCC_readPort_rsp_addr[52 : 51];
  assign popCC_readPort_rsp_lock = _zz_popCC_readPort_rsp_addr[53 : 53];
  assign popCC_readPort_rsp_cache = _zz_popCC_readPort_rsp_addr[57 : 54];
  assign popCC_readPort_rsp_qos = _zz_popCC_readPort_rsp_addr[61 : 58];
  assign popCC_readPort_rsp_prot = _zz_popCC_readPort_rsp_addr[64 : 62];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_addr = popCC_readPort_rsp_addr;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_region = popCC_readPort_rsp_region;
  assign popCC_readArbitation_translated_payload_len = popCC_readPort_rsp_len;
  assign popCC_readArbitation_translated_payload_size = popCC_readPort_rsp_size;
  assign popCC_readArbitation_translated_payload_burst = popCC_readPort_rsp_burst;
  assign popCC_readArbitation_translated_payload_lock = popCC_readPort_rsp_lock;
  assign popCC_readArbitation_translated_payload_cache = popCC_readPort_rsp_cache;
  assign popCC_readArbitation_translated_payload_qos = popCC_readPort_rsp_qos;
  assign popCC_readArbitation_translated_payload_prot = popCC_readPort_rsp_prot;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_addr = popCC_readArbitation_translated_payload_addr;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_region = popCC_readArbitation_translated_payload_region;
  assign io_pop_payload_len = popCC_readArbitation_translated_payload_len;
  assign io_pop_payload_size = popCC_readArbitation_translated_payload_size;
  assign io_pop_payload_burst = popCC_readArbitation_translated_payload_burst;
  assign io_pop_payload_lock = popCC_readArbitation_translated_payload_lock;
  assign io_pop_payload_cache = popCC_readArbitation_translated_payload_cache;
  assign io_pop_payload_qos = popCC_readArbitation_translated_payload_qos;
  assign io_pop_payload_prot = popCC_readArbitation_translated_payload_prot;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1 = system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized;
  always @(posedge io_ddrMasters_0_clk) begin
    if(io_ddrMasters_0_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module Axi4WriteOnlyUpsizer (
  input  wire          io_input_aw_valid,
  output reg           io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [3:0]    io_input_aw_payload_region,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire [0:0]    io_input_aw_payload_lock,
  input  wire [3:0]    io_input_aw_payload_cache,
  input  wire [3:0]    io_input_aw_payload_qos,
  input  wire [2:0]    io_input_aw_payload_prot,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [31:0]   io_input_w_payload_data,
  input  wire [3:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output wire [3:0]    io_input_b_payload_id,
  output wire [1:0]    io_input_b_payload_resp,
  output wire          io_output_aw_valid,
  input  wire          io_output_aw_ready,
  output wire [31:0]   io_output_aw_payload_addr,
  output wire [3:0]    io_output_aw_payload_id,
  output wire [3:0]    io_output_aw_payload_region,
  output reg  [7:0]    io_output_aw_payload_len,
  output reg  [2:0]    io_output_aw_payload_size,
  output wire [1:0]    io_output_aw_payload_burst,
  output wire [0:0]    io_output_aw_payload_lock,
  output wire [3:0]    io_output_aw_payload_cache,
  output wire [3:0]    io_output_aw_payload_qos,
  output wire [2:0]    io_output_aw_payload_prot,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [127:0]  io_output_w_payload_data,
  output wire [15:0]   io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [3:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire       [14:0]   _zz_cmdLogic_byteCount;
  wire       [10:0]   _zz_cmdLogic_incrLen;
  wire       [10:0]   _zz_cmdLogic_incrLen_1;
  wire       [3:0]    _zz_cmdLogic_incrLen_2;
  wire       [4:0]    _zz_dataLogic_byteCounterNext;
  wire       [7:0]    _zz_dataLogic_byteCounterNext_1;
  reg        [15:0]   _zz_dataLogic_byteActivity;
  wire       [1:0]    _zz_dataLogic_byteActivity_1;
  wire                cmdLogic_outputFork_valid;
  wire                cmdLogic_outputFork_ready;
  wire       [31:0]   cmdLogic_outputFork_payload_addr;
  wire       [3:0]    cmdLogic_outputFork_payload_id;
  wire       [3:0]    cmdLogic_outputFork_payload_region;
  wire       [7:0]    cmdLogic_outputFork_payload_len;
  wire       [2:0]    cmdLogic_outputFork_payload_size;
  wire       [1:0]    cmdLogic_outputFork_payload_burst;
  wire       [0:0]    cmdLogic_outputFork_payload_lock;
  wire       [3:0]    cmdLogic_outputFork_payload_cache;
  wire       [3:0]    cmdLogic_outputFork_payload_qos;
  wire       [2:0]    cmdLogic_outputFork_payload_prot;
  wire                cmdLogic_dataFork_valid;
  wire                cmdLogic_dataFork_ready;
  wire       [31:0]   cmdLogic_dataFork_payload_addr;
  wire       [3:0]    cmdLogic_dataFork_payload_id;
  wire       [3:0]    cmdLogic_dataFork_payload_region;
  wire       [7:0]    cmdLogic_dataFork_payload_len;
  wire       [2:0]    cmdLogic_dataFork_payload_size;
  wire       [1:0]    cmdLogic_dataFork_payload_burst;
  wire       [0:0]    cmdLogic_dataFork_payload_lock;
  wire       [3:0]    cmdLogic_dataFork_payload_cache;
  wire       [3:0]    cmdLogic_dataFork_payload_qos;
  wire       [2:0]    cmdLogic_dataFork_payload_prot;
  reg                 io_input_aw_fork2_logic_linkEnable_0;
  reg                 io_input_aw_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdLogic_outputFork_fire;
  wire                cmdLogic_dataFork_fire;
  wire       [9:0]    cmdLogic_byteCount;
  wire       [6:0]    cmdLogic_incrLen;
  wire                when_Axi4Upsizer_l21;
  wire                when_Axi4Upsizer_l24;
  reg        [3:0]    dataLogic_byteCounter;
  reg        [2:0]    dataLogic_size;
  reg                 dataLogic_outputValid;
  reg                 dataLogic_outputLast;
  reg                 dataLogic_busy;
  reg                 dataLogic_incrementByteCounter;
  reg                 dataLogic_alwaysFire;
  wire       [4:0]    dataLogic_byteCounterNext;
  reg        [127:0]  dataLogic_dataBuffer;
  reg        [15:0]   dataLogic_maskBuffer;
  wire       [15:0]   dataLogic_byteActivity;
  wire                io_output_w_fire;
  wire                io_output_w_isStall;
  wire                io_input_w_fire;
  wire                when_Axi4Upsizer_l59;
  wire                when_Axi4Upsizer_l59_1;
  wire                when_Axi4Upsizer_l59_2;
  wire                when_Axi4Upsizer_l59_3;
  wire                when_Axi4Upsizer_l59_4;
  wire                when_Axi4Upsizer_l59_5;
  wire                when_Axi4Upsizer_l59_6;
  wire                when_Axi4Upsizer_l59_7;
  wire                when_Axi4Upsizer_l59_8;
  wire                when_Axi4Upsizer_l59_9;
  wire                when_Axi4Upsizer_l59_10;
  wire                when_Axi4Upsizer_l59_11;
  wire                when_Axi4Upsizer_l59_12;
  wire                when_Axi4Upsizer_l59_13;
  wire                when_Axi4Upsizer_l59_14;
  wire                when_Axi4Upsizer_l59_15;
  wire                when_Axi4Upsizer_l68;
  wire                when_Axi4Upsizer_l68_1;
  wire                when_Axi4Upsizer_l68_2;
  wire                when_Axi4Upsizer_l68_3;

  assign _zz_cmdLogic_byteCount = ({7'd0,io_input_aw_payload_len} <<< io_input_aw_payload_size);
  assign _zz_cmdLogic_incrLen = ({1'b0,cmdLogic_byteCount} + _zz_cmdLogic_incrLen_1);
  assign _zz_cmdLogic_incrLen_2 = io_input_aw_payload_addr[3 : 0];
  assign _zz_cmdLogic_incrLen_1 = {7'd0, _zz_cmdLogic_incrLen_2};
  assign _zz_dataLogic_byteCounterNext_1 = ({7'd0,1'b1} <<< dataLogic_size);
  assign _zz_dataLogic_byteCounterNext = _zz_dataLogic_byteCounterNext_1[4:0];
  assign _zz_dataLogic_byteActivity_1 = dataLogic_size[1:0];
  always @(*) begin
    case(_zz_dataLogic_byteActivity_1)
      2'b00 : _zz_dataLogic_byteActivity = 16'h0001;
      2'b01 : _zz_dataLogic_byteActivity = 16'h0003;
      2'b10 : _zz_dataLogic_byteActivity = 16'h000f;
      default : _zz_dataLogic_byteActivity = 16'h00ff;
    endcase
  end

  always @(*) begin
    io_input_aw_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_input_aw_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_input_aw_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdLogic_outputFork_ready) && io_input_aw_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdLogic_dataFork_ready) && io_input_aw_fork2_logic_linkEnable_1);
  assign cmdLogic_outputFork_valid = (io_input_aw_valid && io_input_aw_fork2_logic_linkEnable_0);
  assign cmdLogic_outputFork_payload_addr = io_input_aw_payload_addr;
  assign cmdLogic_outputFork_payload_id = io_input_aw_payload_id;
  assign cmdLogic_outputFork_payload_region = io_input_aw_payload_region;
  assign cmdLogic_outputFork_payload_len = io_input_aw_payload_len;
  assign cmdLogic_outputFork_payload_size = io_input_aw_payload_size;
  assign cmdLogic_outputFork_payload_burst = io_input_aw_payload_burst;
  assign cmdLogic_outputFork_payload_lock = io_input_aw_payload_lock;
  assign cmdLogic_outputFork_payload_cache = io_input_aw_payload_cache;
  assign cmdLogic_outputFork_payload_qos = io_input_aw_payload_qos;
  assign cmdLogic_outputFork_payload_prot = io_input_aw_payload_prot;
  assign cmdLogic_outputFork_fire = (cmdLogic_outputFork_valid && cmdLogic_outputFork_ready);
  assign cmdLogic_dataFork_valid = (io_input_aw_valid && io_input_aw_fork2_logic_linkEnable_1);
  assign cmdLogic_dataFork_payload_addr = io_input_aw_payload_addr;
  assign cmdLogic_dataFork_payload_id = io_input_aw_payload_id;
  assign cmdLogic_dataFork_payload_region = io_input_aw_payload_region;
  assign cmdLogic_dataFork_payload_len = io_input_aw_payload_len;
  assign cmdLogic_dataFork_payload_size = io_input_aw_payload_size;
  assign cmdLogic_dataFork_payload_burst = io_input_aw_payload_burst;
  assign cmdLogic_dataFork_payload_lock = io_input_aw_payload_lock;
  assign cmdLogic_dataFork_payload_cache = io_input_aw_payload_cache;
  assign cmdLogic_dataFork_payload_qos = io_input_aw_payload_qos;
  assign cmdLogic_dataFork_payload_prot = io_input_aw_payload_prot;
  assign cmdLogic_dataFork_fire = (cmdLogic_dataFork_valid && cmdLogic_dataFork_ready);
  assign io_output_aw_valid = cmdLogic_outputFork_valid;
  assign cmdLogic_outputFork_ready = io_output_aw_ready;
  assign io_output_aw_payload_addr = cmdLogic_outputFork_payload_addr;
  assign io_output_aw_payload_id = cmdLogic_outputFork_payload_id;
  assign io_output_aw_payload_region = cmdLogic_outputFork_payload_region;
  always @(*) begin
    io_output_aw_payload_len = cmdLogic_outputFork_payload_len;
    if(when_Axi4Upsizer_l21) begin
      io_output_aw_payload_len = {1'd0, cmdLogic_incrLen};
    end
  end

  always @(*) begin
    io_output_aw_payload_size = cmdLogic_outputFork_payload_size;
    if(when_Axi4Upsizer_l21) begin
      io_output_aw_payload_size = 3'b100;
      if(when_Axi4Upsizer_l24) begin
        io_output_aw_payload_size = io_input_aw_payload_size;
      end
    end
  end

  assign io_output_aw_payload_burst = cmdLogic_outputFork_payload_burst;
  assign io_output_aw_payload_lock = cmdLogic_outputFork_payload_lock;
  assign io_output_aw_payload_cache = cmdLogic_outputFork_payload_cache;
  assign io_output_aw_payload_qos = cmdLogic_outputFork_payload_qos;
  assign io_output_aw_payload_prot = cmdLogic_outputFork_payload_prot;
  assign cmdLogic_byteCount = _zz_cmdLogic_byteCount[9:0];
  assign cmdLogic_incrLen = _zz_cmdLogic_incrLen[10 : 4];
  assign when_Axi4Upsizer_l21 = (io_output_aw_payload_burst == 2'b01);
  assign when_Axi4Upsizer_l24 = (io_input_aw_payload_len == 8'h0);
  assign dataLogic_byteCounterNext = ({1'b0,dataLogic_byteCounter} + _zz_dataLogic_byteCounterNext);
  assign dataLogic_byteActivity = (_zz_dataLogic_byteActivity <<< dataLogic_byteCounter);
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign io_output_w_valid = dataLogic_outputValid;
  assign io_output_w_isStall = (io_output_w_valid && (! io_output_w_ready));
  assign io_input_w_ready = (dataLogic_busy && (! io_output_w_isStall));
  assign io_output_w_payload_data = dataLogic_dataBuffer;
  assign io_output_w_payload_strb = dataLogic_maskBuffer;
  assign io_output_w_payload_last = dataLogic_outputLast;
  assign io_input_w_fire = (io_input_w_valid && io_input_w_ready);
  assign when_Axi4Upsizer_l59 = dataLogic_byteActivity[0];
  assign when_Axi4Upsizer_l59_1 = dataLogic_byteActivity[1];
  assign when_Axi4Upsizer_l59_2 = dataLogic_byteActivity[2];
  assign when_Axi4Upsizer_l59_3 = dataLogic_byteActivity[3];
  assign when_Axi4Upsizer_l59_4 = dataLogic_byteActivity[4];
  assign when_Axi4Upsizer_l59_5 = dataLogic_byteActivity[5];
  assign when_Axi4Upsizer_l59_6 = dataLogic_byteActivity[6];
  assign when_Axi4Upsizer_l59_7 = dataLogic_byteActivity[7];
  assign when_Axi4Upsizer_l59_8 = dataLogic_byteActivity[8];
  assign when_Axi4Upsizer_l59_9 = dataLogic_byteActivity[9];
  assign when_Axi4Upsizer_l59_10 = dataLogic_byteActivity[10];
  assign when_Axi4Upsizer_l59_11 = dataLogic_byteActivity[11];
  assign when_Axi4Upsizer_l59_12 = dataLogic_byteActivity[12];
  assign when_Axi4Upsizer_l59_13 = dataLogic_byteActivity[13];
  assign when_Axi4Upsizer_l59_14 = dataLogic_byteActivity[14];
  assign when_Axi4Upsizer_l59_15 = dataLogic_byteActivity[15];
  assign when_Axi4Upsizer_l68 = (3'b000 < cmdLogic_dataFork_payload_size);
  assign when_Axi4Upsizer_l68_1 = (3'b001 < cmdLogic_dataFork_payload_size);
  assign when_Axi4Upsizer_l68_2 = (3'b010 < cmdLogic_dataFork_payload_size);
  assign when_Axi4Upsizer_l68_3 = (3'b011 < cmdLogic_dataFork_payload_size);
  assign cmdLogic_dataFork_ready = (! dataLogic_busy);
  assign io_input_b_valid = io_output_b_valid;
  assign io_output_b_ready = io_input_b_ready;
  assign io_input_b_payload_id = io_output_b_payload_id;
  assign io_input_b_payload_resp = io_output_b_payload_resp;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      io_input_aw_fork2_logic_linkEnable_0 <= 1'b1;
      io_input_aw_fork2_logic_linkEnable_1 <= 1'b1;
      dataLogic_outputValid <= 1'b0;
      dataLogic_busy <= 1'b0;
      dataLogic_maskBuffer <= 16'h0;
    end else begin
      if(cmdLogic_outputFork_fire) begin
        io_input_aw_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdLogic_dataFork_fire) begin
        io_input_aw_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_aw_ready) begin
        io_input_aw_fork2_logic_linkEnable_0 <= 1'b1;
        io_input_aw_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(io_output_w_ready) begin
        dataLogic_outputValid <= 1'b0;
      end
      if(io_output_w_fire) begin
        dataLogic_maskBuffer <= 16'h0;
      end
      if(io_input_w_fire) begin
        dataLogic_outputValid <= ((dataLogic_byteCounterNext[4] || io_input_w_payload_last) || dataLogic_alwaysFire);
        if(io_input_w_payload_last) begin
          dataLogic_busy <= 1'b0;
        end
        if(when_Axi4Upsizer_l59) begin
          dataLogic_maskBuffer[0] <= io_input_w_payload_strb[0];
        end
        if(when_Axi4Upsizer_l59_1) begin
          dataLogic_maskBuffer[1] <= io_input_w_payload_strb[1];
        end
        if(when_Axi4Upsizer_l59_2) begin
          dataLogic_maskBuffer[2] <= io_input_w_payload_strb[2];
        end
        if(when_Axi4Upsizer_l59_3) begin
          dataLogic_maskBuffer[3] <= io_input_w_payload_strb[3];
        end
        if(when_Axi4Upsizer_l59_4) begin
          dataLogic_maskBuffer[4] <= io_input_w_payload_strb[0];
        end
        if(when_Axi4Upsizer_l59_5) begin
          dataLogic_maskBuffer[5] <= io_input_w_payload_strb[1];
        end
        if(when_Axi4Upsizer_l59_6) begin
          dataLogic_maskBuffer[6] <= io_input_w_payload_strb[2];
        end
        if(when_Axi4Upsizer_l59_7) begin
          dataLogic_maskBuffer[7] <= io_input_w_payload_strb[3];
        end
        if(when_Axi4Upsizer_l59_8) begin
          dataLogic_maskBuffer[8] <= io_input_w_payload_strb[0];
        end
        if(when_Axi4Upsizer_l59_9) begin
          dataLogic_maskBuffer[9] <= io_input_w_payload_strb[1];
        end
        if(when_Axi4Upsizer_l59_10) begin
          dataLogic_maskBuffer[10] <= io_input_w_payload_strb[2];
        end
        if(when_Axi4Upsizer_l59_11) begin
          dataLogic_maskBuffer[11] <= io_input_w_payload_strb[3];
        end
        if(when_Axi4Upsizer_l59_12) begin
          dataLogic_maskBuffer[12] <= io_input_w_payload_strb[0];
        end
        if(when_Axi4Upsizer_l59_13) begin
          dataLogic_maskBuffer[13] <= io_input_w_payload_strb[1];
        end
        if(when_Axi4Upsizer_l59_14) begin
          dataLogic_maskBuffer[14] <= io_input_w_payload_strb[2];
        end
        if(when_Axi4Upsizer_l59_15) begin
          dataLogic_maskBuffer[15] <= io_input_w_payload_strb[3];
        end
      end
      if(cmdLogic_dataFork_fire) begin
        dataLogic_busy <= 1'b1;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(io_input_w_fire) begin
      if(dataLogic_incrementByteCounter) begin
        dataLogic_byteCounter <= dataLogic_byteCounterNext[3:0];
      end
      dataLogic_outputLast <= io_input_w_payload_last;
      if(when_Axi4Upsizer_l59) begin
        dataLogic_dataBuffer[7 : 0] <= io_input_w_payload_data[7 : 0];
      end
      if(when_Axi4Upsizer_l59_1) begin
        dataLogic_dataBuffer[15 : 8] <= io_input_w_payload_data[15 : 8];
      end
      if(when_Axi4Upsizer_l59_2) begin
        dataLogic_dataBuffer[23 : 16] <= io_input_w_payload_data[23 : 16];
      end
      if(when_Axi4Upsizer_l59_3) begin
        dataLogic_dataBuffer[31 : 24] <= io_input_w_payload_data[31 : 24];
      end
      if(when_Axi4Upsizer_l59_4) begin
        dataLogic_dataBuffer[39 : 32] <= io_input_w_payload_data[7 : 0];
      end
      if(when_Axi4Upsizer_l59_5) begin
        dataLogic_dataBuffer[47 : 40] <= io_input_w_payload_data[15 : 8];
      end
      if(when_Axi4Upsizer_l59_6) begin
        dataLogic_dataBuffer[55 : 48] <= io_input_w_payload_data[23 : 16];
      end
      if(when_Axi4Upsizer_l59_7) begin
        dataLogic_dataBuffer[63 : 56] <= io_input_w_payload_data[31 : 24];
      end
      if(when_Axi4Upsizer_l59_8) begin
        dataLogic_dataBuffer[71 : 64] <= io_input_w_payload_data[7 : 0];
      end
      if(when_Axi4Upsizer_l59_9) begin
        dataLogic_dataBuffer[79 : 72] <= io_input_w_payload_data[15 : 8];
      end
      if(when_Axi4Upsizer_l59_10) begin
        dataLogic_dataBuffer[87 : 80] <= io_input_w_payload_data[23 : 16];
      end
      if(when_Axi4Upsizer_l59_11) begin
        dataLogic_dataBuffer[95 : 88] <= io_input_w_payload_data[31 : 24];
      end
      if(when_Axi4Upsizer_l59_12) begin
        dataLogic_dataBuffer[103 : 96] <= io_input_w_payload_data[7 : 0];
      end
      if(when_Axi4Upsizer_l59_13) begin
        dataLogic_dataBuffer[111 : 104] <= io_input_w_payload_data[15 : 8];
      end
      if(when_Axi4Upsizer_l59_14) begin
        dataLogic_dataBuffer[119 : 112] <= io_input_w_payload_data[23 : 16];
      end
      if(when_Axi4Upsizer_l59_15) begin
        dataLogic_dataBuffer[127 : 120] <= io_input_w_payload_data[31 : 24];
      end
    end
    if(cmdLogic_dataFork_fire) begin
      dataLogic_byteCounter <= cmdLogic_dataFork_payload_addr[3:0];
      if(when_Axi4Upsizer_l68) begin
        dataLogic_byteCounter[0] <= 1'b0;
      end
      if(when_Axi4Upsizer_l68_1) begin
        dataLogic_byteCounter[1] <= 1'b0;
      end
      if(when_Axi4Upsizer_l68_2) begin
        dataLogic_byteCounter[2] <= 1'b0;
      end
      if(when_Axi4Upsizer_l68_3) begin
        dataLogic_byteCounter[3] <= 1'b0;
      end
      dataLogic_size <= cmdLogic_dataFork_payload_size;
      dataLogic_alwaysFire <= (! (cmdLogic_dataFork_payload_burst == 2'b01));
      dataLogic_incrementByteCounter <= (! (cmdLogic_dataFork_payload_burst == 2'b00));
    end
  end


endmodule

module Axi4ReadOnlyUpsizer (
  input  wire          io_input_ar_valid,
  output reg           io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [3:0]    io_input_ar_payload_region,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  input  wire [0:0]    io_input_ar_payload_lock,
  input  wire [3:0]    io_input_ar_payload_cache,
  input  wire [3:0]    io_input_ar_payload_qos,
  input  wire [2:0]    io_input_ar_payload_prot,
  output wire          io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [31:0]   io_input_r_payload_data,
  output wire [3:0]    io_input_r_payload_id,
  output wire [1:0]    io_input_r_payload_resp,
  output wire          io_input_r_payload_last,
  output wire          io_output_ar_valid,
  input  wire          io_output_ar_ready,
  output wire [31:0]   io_output_ar_payload_addr,
  output wire [3:0]    io_output_ar_payload_id,
  output wire [3:0]    io_output_ar_payload_region,
  output wire [7:0]    io_output_ar_payload_len,
  output reg  [2:0]    io_output_ar_payload_size,
  output wire [1:0]    io_output_ar_payload_burst,
  output wire [0:0]    io_output_ar_payload_lock,
  output wire [3:0]    io_output_ar_payload_cache,
  output wire [3:0]    io_output_ar_payload_qos,
  output wire [2:0]    io_output_ar_payload_prot,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [127:0]  io_output_r_payload_data,
  input  wire [3:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                dataLogic_cmdPush_fifo_io_pop_ready;
  wire                dataLogic_cmdPush_fifo_io_push_ready;
  wire                dataLogic_cmdPush_fifo_io_pop_valid;
  wire       [3:0]    dataLogic_cmdPush_fifo_io_pop_payload_startAt;
  wire       [3:0]    dataLogic_cmdPush_fifo_io_pop_payload_endAt;
  wire       [2:0]    dataLogic_cmdPush_fifo_io_pop_payload_size;
  wire       [3:0]    dataLogic_cmdPush_fifo_io_pop_payload_id;
  wire       [2:0]    dataLogic_cmdPush_fifo_io_occupancy;
  wire       [2:0]    dataLogic_cmdPush_fifo_io_availability;
  wire       [14:0]   _zz_cmdLogic_byteCount;
  wire       [10:0]   _zz_cmdLogic_incrLen;
  wire       [10:0]   _zz_cmdLogic_incrLen_1;
  wire       [3:0]    _zz_cmdLogic_incrLen_2;
  wire       [31:0]   _zz_dataLogic_cmdPush_payload_endAt;
  wire       [31:0]   _zz_dataLogic_cmdPush_payload_endAt_1;
  wire       [14:0]   _zz_dataLogic_cmdPush_payload_endAt_2;
  wire       [4:0]    _zz_dataLogic_byteCounterNext;
  wire       [7:0]    _zz_dataLogic_byteCounterNext_1;
  reg        [31:0]   _zz_io_input_r_payload_data;
  wire       [1:0]    _zz_io_input_r_payload_data_1;
  wire                cmdLogic_outputFork_valid;
  wire                cmdLogic_outputFork_ready;
  wire       [31:0]   cmdLogic_outputFork_payload_addr;
  wire       [3:0]    cmdLogic_outputFork_payload_id;
  wire       [3:0]    cmdLogic_outputFork_payload_region;
  wire       [7:0]    cmdLogic_outputFork_payload_len;
  wire       [2:0]    cmdLogic_outputFork_payload_size;
  wire       [1:0]    cmdLogic_outputFork_payload_burst;
  wire       [0:0]    cmdLogic_outputFork_payload_lock;
  wire       [3:0]    cmdLogic_outputFork_payload_cache;
  wire       [3:0]    cmdLogic_outputFork_payload_qos;
  wire       [2:0]    cmdLogic_outputFork_payload_prot;
  wire                cmdLogic_dataFork_valid;
  wire                cmdLogic_dataFork_ready;
  wire       [31:0]   cmdLogic_dataFork_payload_addr;
  wire       [3:0]    cmdLogic_dataFork_payload_id;
  wire       [3:0]    cmdLogic_dataFork_payload_region;
  wire       [7:0]    cmdLogic_dataFork_payload_len;
  wire       [2:0]    cmdLogic_dataFork_payload_size;
  wire       [1:0]    cmdLogic_dataFork_payload_burst;
  wire       [0:0]    cmdLogic_dataFork_payload_lock;
  wire       [3:0]    cmdLogic_dataFork_payload_cache;
  wire       [3:0]    cmdLogic_dataFork_payload_qos;
  wire       [2:0]    cmdLogic_dataFork_payload_prot;
  reg                 io_input_ar_fork2_logic_linkEnable_0;
  reg                 io_input_ar_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdLogic_outputFork_fire;
  wire                cmdLogic_dataFork_fire;
  wire       [9:0]    cmdLogic_byteCount;
  wire       [6:0]    cmdLogic_incrLen;
  wire                when_Axi4Upsizer_l108;
  wire                dataLogic_cmdPush_valid;
  wire                dataLogic_cmdPush_ready;
  wire       [3:0]    dataLogic_cmdPush_payload_startAt;
  wire       [3:0]    dataLogic_cmdPush_payload_endAt;
  wire       [2:0]    dataLogic_cmdPush_payload_size;
  wire       [3:0]    dataLogic_cmdPush_payload_id;
  reg        [2:0]    dataLogic_size;
  reg                 dataLogic_busy;
  reg        [3:0]    dataLogic_id;
  reg        [3:0]    dataLogic_byteCounter;
  reg        [3:0]    dataLogic_byteCounterLast;
  wire       [4:0]    dataLogic_byteCounterNext;
  wire                dataLogic_cmdPush_fifo_io_pop_fire;
  wire                io_input_r_fire;

  assign _zz_cmdLogic_byteCount = ({7'd0,io_input_ar_payload_len} <<< io_input_ar_payload_size);
  assign _zz_cmdLogic_incrLen = ({1'b0,cmdLogic_byteCount} + _zz_cmdLogic_incrLen_1);
  assign _zz_cmdLogic_incrLen_2 = io_input_ar_payload_addr[3 : 0];
  assign _zz_cmdLogic_incrLen_1 = {7'd0, _zz_cmdLogic_incrLen_2};
  assign _zz_dataLogic_cmdPush_payload_endAt = (cmdLogic_dataFork_payload_addr + _zz_dataLogic_cmdPush_payload_endAt_1);
  assign _zz_dataLogic_cmdPush_payload_endAt_2 = ({7'd0,cmdLogic_dataFork_payload_len} <<< cmdLogic_dataFork_payload_size);
  assign _zz_dataLogic_cmdPush_payload_endAt_1 = {17'd0, _zz_dataLogic_cmdPush_payload_endAt_2};
  assign _zz_dataLogic_byteCounterNext_1 = ({7'd0,1'b1} <<< dataLogic_size);
  assign _zz_dataLogic_byteCounterNext = _zz_dataLogic_byteCounterNext_1[4:0];
  assign _zz_io_input_r_payload_data_1 = (dataLogic_byteCounter >>> 2'd2);
  StreamFifo_4 dataLogic_cmdPush_fifo (
    .io_push_valid           (dataLogic_cmdPush_valid                           ), //i
    .io_push_ready           (dataLogic_cmdPush_fifo_io_push_ready              ), //o
    .io_push_payload_startAt (dataLogic_cmdPush_payload_startAt[3:0]            ), //i
    .io_push_payload_endAt   (dataLogic_cmdPush_payload_endAt[3:0]              ), //i
    .io_push_payload_size    (dataLogic_cmdPush_payload_size[2:0]               ), //i
    .io_push_payload_id      (dataLogic_cmdPush_payload_id[3:0]                 ), //i
    .io_pop_valid            (dataLogic_cmdPush_fifo_io_pop_valid               ), //o
    .io_pop_ready            (dataLogic_cmdPush_fifo_io_pop_ready               ), //i
    .io_pop_payload_startAt  (dataLogic_cmdPush_fifo_io_pop_payload_startAt[3:0]), //o
    .io_pop_payload_endAt    (dataLogic_cmdPush_fifo_io_pop_payload_endAt[3:0]  ), //o
    .io_pop_payload_size     (dataLogic_cmdPush_fifo_io_pop_payload_size[2:0]   ), //o
    .io_pop_payload_id       (dataLogic_cmdPush_fifo_io_pop_payload_id[3:0]     ), //o
    .io_flush                (1'b0                                              ), //i
    .io_occupancy            (dataLogic_cmdPush_fifo_io_occupancy[2:0]          ), //o
    .io_availability         (dataLogic_cmdPush_fifo_io_availability[2:0]       ), //o
    .io_memoryClk            (io_memoryClk                                      ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                           )  //i
  );
  always @(*) begin
    case(_zz_io_input_r_payload_data_1)
      2'b00 : _zz_io_input_r_payload_data = io_output_r_payload_data[31 : 0];
      2'b01 : _zz_io_input_r_payload_data = io_output_r_payload_data[63 : 32];
      2'b10 : _zz_io_input_r_payload_data = io_output_r_payload_data[95 : 64];
      default : _zz_io_input_r_payload_data = io_output_r_payload_data[127 : 96];
    endcase
  end

  always @(*) begin
    io_input_ar_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_input_ar_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_input_ar_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdLogic_outputFork_ready) && io_input_ar_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdLogic_dataFork_ready) && io_input_ar_fork2_logic_linkEnable_1);
  assign cmdLogic_outputFork_valid = (io_input_ar_valid && io_input_ar_fork2_logic_linkEnable_0);
  assign cmdLogic_outputFork_payload_addr = io_input_ar_payload_addr;
  assign cmdLogic_outputFork_payload_id = io_input_ar_payload_id;
  assign cmdLogic_outputFork_payload_region = io_input_ar_payload_region;
  assign cmdLogic_outputFork_payload_len = io_input_ar_payload_len;
  assign cmdLogic_outputFork_payload_size = io_input_ar_payload_size;
  assign cmdLogic_outputFork_payload_burst = io_input_ar_payload_burst;
  assign cmdLogic_outputFork_payload_lock = io_input_ar_payload_lock;
  assign cmdLogic_outputFork_payload_cache = io_input_ar_payload_cache;
  assign cmdLogic_outputFork_payload_qos = io_input_ar_payload_qos;
  assign cmdLogic_outputFork_payload_prot = io_input_ar_payload_prot;
  assign cmdLogic_outputFork_fire = (cmdLogic_outputFork_valid && cmdLogic_outputFork_ready);
  assign cmdLogic_dataFork_valid = (io_input_ar_valid && io_input_ar_fork2_logic_linkEnable_1);
  assign cmdLogic_dataFork_payload_addr = io_input_ar_payload_addr;
  assign cmdLogic_dataFork_payload_id = io_input_ar_payload_id;
  assign cmdLogic_dataFork_payload_region = io_input_ar_payload_region;
  assign cmdLogic_dataFork_payload_len = io_input_ar_payload_len;
  assign cmdLogic_dataFork_payload_size = io_input_ar_payload_size;
  assign cmdLogic_dataFork_payload_burst = io_input_ar_payload_burst;
  assign cmdLogic_dataFork_payload_lock = io_input_ar_payload_lock;
  assign cmdLogic_dataFork_payload_cache = io_input_ar_payload_cache;
  assign cmdLogic_dataFork_payload_qos = io_input_ar_payload_qos;
  assign cmdLogic_dataFork_payload_prot = io_input_ar_payload_prot;
  assign cmdLogic_dataFork_fire = (cmdLogic_dataFork_valid && cmdLogic_dataFork_ready);
  assign io_output_ar_valid = cmdLogic_outputFork_valid;
  assign cmdLogic_outputFork_ready = io_output_ar_ready;
  assign io_output_ar_payload_addr = cmdLogic_outputFork_payload_addr;
  assign io_output_ar_payload_region = cmdLogic_outputFork_payload_region;
  assign io_output_ar_payload_burst = cmdLogic_outputFork_payload_burst;
  assign io_output_ar_payload_lock = cmdLogic_outputFork_payload_lock;
  assign io_output_ar_payload_cache = cmdLogic_outputFork_payload_cache;
  assign io_output_ar_payload_qos = cmdLogic_outputFork_payload_qos;
  assign io_output_ar_payload_prot = cmdLogic_outputFork_payload_prot;
  assign cmdLogic_byteCount = _zz_cmdLogic_byteCount[9:0];
  assign cmdLogic_incrLen = _zz_cmdLogic_incrLen[10 : 4];
  always @(*) begin
    io_output_ar_payload_size = 3'b100;
    if(when_Axi4Upsizer_l108) begin
      io_output_ar_payload_size = io_input_ar_payload_size;
    end
  end

  assign io_output_ar_payload_len = {1'd0, cmdLogic_incrLen};
  assign io_output_ar_payload_id = 4'b0000;
  assign when_Axi4Upsizer_l108 = (io_input_ar_payload_len == 8'h0);
  assign dataLogic_cmdPush_valid = cmdLogic_dataFork_valid;
  assign cmdLogic_dataFork_ready = dataLogic_cmdPush_ready;
  assign dataLogic_cmdPush_payload_startAt = cmdLogic_dataFork_payload_addr[3:0];
  assign dataLogic_cmdPush_payload_endAt = _zz_dataLogic_cmdPush_payload_endAt[3:0];
  assign dataLogic_cmdPush_payload_size = cmdLogic_dataFork_payload_size;
  assign dataLogic_cmdPush_payload_id = cmdLogic_dataFork_payload_id;
  assign dataLogic_cmdPush_ready = dataLogic_cmdPush_fifo_io_push_ready;
  assign dataLogic_byteCounterNext = ({1'b0,dataLogic_byteCounter} + _zz_dataLogic_byteCounterNext);
  assign dataLogic_cmdPush_fifo_io_pop_fire = (dataLogic_cmdPush_fifo_io_pop_valid && dataLogic_cmdPush_fifo_io_pop_ready);
  assign dataLogic_cmdPush_fifo_io_pop_ready = (! dataLogic_busy);
  assign io_input_r_fire = (io_input_r_valid && io_input_r_ready);
  assign io_input_r_valid = (io_output_r_valid && dataLogic_busy);
  assign io_input_r_payload_last = (io_output_r_payload_last && (dataLogic_byteCounter == dataLogic_byteCounterLast));
  assign io_input_r_payload_resp = io_output_r_payload_resp;
  assign io_input_r_payload_data = _zz_io_input_r_payload_data;
  assign io_input_r_payload_id = dataLogic_id;
  assign io_output_r_ready = ((dataLogic_busy && io_input_r_ready) && (io_input_r_payload_last || dataLogic_byteCounterNext[4]));
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      io_input_ar_fork2_logic_linkEnable_0 <= 1'b1;
      io_input_ar_fork2_logic_linkEnable_1 <= 1'b1;
      dataLogic_busy <= 1'b0;
    end else begin
      if(cmdLogic_outputFork_fire) begin
        io_input_ar_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdLogic_dataFork_fire) begin
        io_input_ar_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_ar_ready) begin
        io_input_ar_fork2_logic_linkEnable_0 <= 1'b1;
        io_input_ar_fork2_logic_linkEnable_1 <= 1'b1;
      end
      if(dataLogic_cmdPush_fifo_io_pop_fire) begin
        dataLogic_busy <= 1'b1;
      end
      if(io_input_r_fire) begin
        if(io_input_r_payload_last) begin
          dataLogic_busy <= 1'b0;
        end
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(dataLogic_cmdPush_fifo_io_pop_fire) begin
      dataLogic_byteCounter <= dataLogic_cmdPush_fifo_io_pop_payload_startAt;
      dataLogic_byteCounterLast <= dataLogic_cmdPush_fifo_io_pop_payload_endAt;
      dataLogic_size <= dataLogic_cmdPush_fifo_io_pop_payload_size;
      dataLogic_id <= dataLogic_cmdPush_fifo_io_pop_payload_id;
    end
    if(io_input_r_fire) begin
      dataLogic_byteCounter <= dataLogic_byteCounterNext[3:0];
    end
  end


endmodule

module StreamFifoCC_6 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [3:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [3:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset,
  input  wire          io_ddrMasters_1_clk,
  input  wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1
);

  reg        [5:0]    ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [5:0]    _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [1:0]    popCC_readPort_rsp_resp;
  wire       [5:0]    _zz_popCC_readPort_rsp_id;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [1:0]    popCC_readArbitation_translated_payload_resp;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [5:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_resp,io_push_payload_id};
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_14 popToPushGray_buffercc (
    .io_dataIn               (popToPushGray[4:0]                    ), //i
    .io_dataOut              (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_memoryClk            (io_memoryClk                          ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_22 pushToPopGray_buffercc (
    .io_dataIn                                                                                 (pushToPopGray[4:0]                                                                       ), //i
    .io_dataOut                                                                                (pushToPopGray_buffercc_io_dataOut[4:0]                                                   ), //o
    .io_ddrMasters_1_clk                                                                       (io_ddrMasters_1_clk                                                                      ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_id = ram_spinal_port1;
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_id[3 : 0];
  assign popCC_readPort_rsp_resp = _zz_popCC_readPort_rsp_id[5 : 4];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_resp = popCC_readPort_rsp_resp;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = popCC_readArbitation_translated_payload_resp;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_5 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_data,
  input  wire [3:0]    io_push_payload_strb,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_data,
  output wire [3:0]    io_pop_payload_strb,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_ddrMasters_1_clk,
  input  wire          io_ddrMasters_1_reset,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1
);

  reg        [36:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [36:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [31:0]   popCC_readPort_rsp_data;
  wire       [3:0]    popCC_readPort_rsp_strb;
  wire                popCC_readPort_rsp_last;
  wire       [36:0]   _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [31:0]   popCC_readArbitation_translated_payload_data;
  wire       [3:0]    popCC_readArbitation_translated_payload_strb;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [36:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_strb,io_push_payload_data}};
  always @(posedge io_ddrMasters_1_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_11 popToPushGray_buffercc (
    .io_dataIn             (popToPushGray[4:0]                    ), //i
    .io_dataOut            (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_ddrMasters_1_clk   (io_ddrMasters_1_clk                   ), //i
    .io_ddrMasters_1_reset (io_ddrMasters_1_reset                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_18 pushToPopGray_buffercc (
    .io_dataIn                                                                               (pushToPopGray[4:0]                                                                     ), //i
    .io_dataOut                                                                              (pushToPopGray_buffercc_io_dataOut[4:0]                                                 ), //o
    .io_memoryClk                                                                            (io_memoryClk                                                                           ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1 (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[31 : 0];
  assign popCC_readPort_rsp_strb = _zz_popCC_readPort_rsp_data[35 : 32];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[36];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_strb = popCC_readPort_rsp_strb;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_strb = popCC_readArbitation_translated_payload_strb;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_ddrMasters_1_clk) begin
    if(io_ddrMasters_1_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_4 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_addr,
  input  wire [3:0]    io_push_payload_id,
  input  wire [3:0]    io_push_payload_region,
  input  wire [7:0]    io_push_payload_len,
  input  wire [2:0]    io_push_payload_size,
  input  wire [1:0]    io_push_payload_burst,
  input  wire [0:0]    io_push_payload_lock,
  input  wire [3:0]    io_push_payload_cache,
  input  wire [3:0]    io_push_payload_qos,
  input  wire [2:0]    io_push_payload_prot,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_addr,
  output wire [3:0]    io_pop_payload_id,
  output wire [3:0]    io_pop_payload_region,
  output wire [7:0]    io_pop_payload_len,
  output wire [2:0]    io_pop_payload_size,
  output wire [1:0]    io_pop_payload_burst,
  output wire [0:0]    io_pop_payload_lock,
  output wire [3:0]    io_pop_payload_cache,
  output wire [3:0]    io_pop_payload_qos,
  output wire [2:0]    io_pop_payload_prot,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_ddrMasters_1_clk,
  input  wire          io_ddrMasters_1_reset,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1
);

  reg        [64:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [64:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [31:0]   popCC_readPort_rsp_addr;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [3:0]    popCC_readPort_rsp_region;
  wire       [7:0]    popCC_readPort_rsp_len;
  wire       [2:0]    popCC_readPort_rsp_size;
  wire       [1:0]    popCC_readPort_rsp_burst;
  wire       [0:0]    popCC_readPort_rsp_lock;
  wire       [3:0]    popCC_readPort_rsp_cache;
  wire       [3:0]    popCC_readPort_rsp_qos;
  wire       [2:0]    popCC_readPort_rsp_prot;
  wire       [64:0]   _zz_popCC_readPort_rsp_addr;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [31:0]   popCC_readArbitation_translated_payload_addr;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [3:0]    popCC_readArbitation_translated_payload_region;
  wire       [7:0]    popCC_readArbitation_translated_payload_len;
  wire       [2:0]    popCC_readArbitation_translated_payload_size;
  wire       [1:0]    popCC_readArbitation_translated_payload_burst;
  wire       [0:0]    popCC_readArbitation_translated_payload_lock;
  wire       [3:0]    popCC_readArbitation_translated_payload_cache;
  wire       [3:0]    popCC_readArbitation_translated_payload_qos;
  wire       [2:0]    popCC_readArbitation_translated_payload_prot;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [64:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_prot,{io_push_payload_qos,{io_push_payload_cache,{io_push_payload_lock,{io_push_payload_burst,{io_push_payload_size,{io_push_payload_len,{io_push_payload_region,{io_push_payload_id,io_push_payload_addr}}}}}}}}};
  always @(posedge io_ddrMasters_1_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_11 popToPushGray_buffercc (
    .io_dataIn             (popToPushGray[4:0]                    ), //i
    .io_dataOut            (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_ddrMasters_1_clk   (io_ddrMasters_1_clk                   ), //i
    .io_ddrMasters_1_reset (io_ddrMasters_1_reset                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_18 pushToPopGray_buffercc (
    .io_dataIn                                                                               (pushToPopGray[4:0]                                                                     ), //i
    .io_dataOut                                                                              (pushToPopGray_buffercc_io_dataOut[4:0]                                                 ), //o
    .io_memoryClk                                                                            (io_memoryClk                                                                           ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1 (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_addr = ram_spinal_port1;
  assign popCC_readPort_rsp_addr = _zz_popCC_readPort_rsp_addr[31 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_addr[35 : 32];
  assign popCC_readPort_rsp_region = _zz_popCC_readPort_rsp_addr[39 : 36];
  assign popCC_readPort_rsp_len = _zz_popCC_readPort_rsp_addr[47 : 40];
  assign popCC_readPort_rsp_size = _zz_popCC_readPort_rsp_addr[50 : 48];
  assign popCC_readPort_rsp_burst = _zz_popCC_readPort_rsp_addr[52 : 51];
  assign popCC_readPort_rsp_lock = _zz_popCC_readPort_rsp_addr[53 : 53];
  assign popCC_readPort_rsp_cache = _zz_popCC_readPort_rsp_addr[57 : 54];
  assign popCC_readPort_rsp_qos = _zz_popCC_readPort_rsp_addr[61 : 58];
  assign popCC_readPort_rsp_prot = _zz_popCC_readPort_rsp_addr[64 : 62];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_addr = popCC_readPort_rsp_addr;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_region = popCC_readPort_rsp_region;
  assign popCC_readArbitation_translated_payload_len = popCC_readPort_rsp_len;
  assign popCC_readArbitation_translated_payload_size = popCC_readPort_rsp_size;
  assign popCC_readArbitation_translated_payload_burst = popCC_readPort_rsp_burst;
  assign popCC_readArbitation_translated_payload_lock = popCC_readPort_rsp_lock;
  assign popCC_readArbitation_translated_payload_cache = popCC_readPort_rsp_cache;
  assign popCC_readArbitation_translated_payload_qos = popCC_readPort_rsp_qos;
  assign popCC_readArbitation_translated_payload_prot = popCC_readPort_rsp_prot;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_addr = popCC_readArbitation_translated_payload_addr;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_region = popCC_readArbitation_translated_payload_region;
  assign io_pop_payload_len = popCC_readArbitation_translated_payload_len;
  assign io_pop_payload_size = popCC_readArbitation_translated_payload_size;
  assign io_pop_payload_burst = popCC_readArbitation_translated_payload_burst;
  assign io_pop_payload_lock = popCC_readArbitation_translated_payload_lock;
  assign io_pop_payload_cache = popCC_readArbitation_translated_payload_cache;
  assign io_pop_payload_qos = popCC_readArbitation_translated_payload_qos;
  assign io_pop_payload_prot = popCC_readArbitation_translated_payload_prot;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_ddrMasters_1_clk) begin
    if(io_ddrMasters_1_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_3 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_data,
  input  wire [3:0]    io_push_payload_id,
  input  wire [1:0]    io_push_payload_resp,
  input  wire          io_push_payload_last,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_data,
  output wire [3:0]    io_pop_payload_id,
  output wire [1:0]    io_pop_payload_resp,
  output wire          io_pop_payload_last,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset,
  input  wire          io_ddrMasters_1_clk,
  output wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1
);

  reg        [38:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [38:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [31:0]   popCC_readPort_rsp_data;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [1:0]    popCC_readPort_rsp_resp;
  wire                popCC_readPort_rsp_last;
  wire       [38:0]   _zz_popCC_readPort_rsp_data;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [31:0]   popCC_readArbitation_translated_payload_data;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [1:0]    popCC_readArbitation_translated_payload_resp;
  wire                popCC_readArbitation_translated_payload_last;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [38:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_last,{io_push_payload_resp,{io_push_payload_id,io_push_payload_data}}};
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_14 popToPushGray_buffercc (
    .io_dataIn               (popToPushGray[4:0]                    ), //i
    .io_dataOut              (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_memoryClk            (io_memoryClk                          ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_15 system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn               (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut              (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_ddrMasters_1_clk     (io_ddrMasters_1_clk                                                                                                   ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                                                                                               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_16 pushToPopGray_buffercc (
    .io_dataIn                                                                               (pushToPopGray[4:0]                                                                     ), //i
    .io_dataOut                                                                              (pushToPopGray_buffercc_io_dataOut[4:0]                                                 ), //o
    .io_ddrMasters_1_clk                                                                     (io_ddrMasters_1_clk                                                                    ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized = system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_data = ram_spinal_port1;
  assign popCC_readPort_rsp_data = _zz_popCC_readPort_rsp_data[31 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_data[35 : 32];
  assign popCC_readPort_rsp_resp = _zz_popCC_readPort_rsp_data[37 : 36];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_data[38];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_data = popCC_readPort_rsp_data;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_resp = popCC_readPort_rsp_resp;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_data = popCC_readArbitation_translated_payload_data;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_resp = popCC_readArbitation_translated_payload_resp;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1 = system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_ddrMasters_1_clk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC_2 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_addr,
  input  wire [3:0]    io_push_payload_id,
  input  wire [3:0]    io_push_payload_region,
  input  wire [7:0]    io_push_payload_len,
  input  wire [2:0]    io_push_payload_size,
  input  wire [1:0]    io_push_payload_burst,
  input  wire [0:0]    io_push_payload_lock,
  input  wire [3:0]    io_push_payload_cache,
  input  wire [3:0]    io_push_payload_qos,
  input  wire [2:0]    io_push_payload_prot,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_addr,
  output wire [3:0]    io_pop_payload_id,
  output wire [3:0]    io_pop_payload_region,
  output wire [7:0]    io_pop_payload_len,
  output wire [2:0]    io_pop_payload_size,
  output wire [1:0]    io_pop_payload_burst,
  output wire [0:0]    io_pop_payload_lock,
  output wire [3:0]    io_pop_payload_cache,
  output wire [3:0]    io_pop_payload_qos,
  output wire [2:0]    io_pop_payload_prot,
  output wire [4:0]    io_pushOccupancy,
  output wire [4:0]    io_popOccupancy,
  input  wire          io_ddrMasters_1_clk,
  input  wire          io_ddrMasters_1_reset,
  input  wire          io_memoryClk,
  output wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1
);

  reg        [64:0]   ram_spinal_port1;
  wire       [4:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [4:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [4:0]    _zz_pushCC_pushPtrGray;
  wire       [3:0]    _zz_ram_port;
  wire       [64:0]   _zz_ram_port_1;
  wire       [4:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [4:0]    popToPushGray;
  wire       [4:0]    pushToPopGray;
  reg        [4:0]    pushCC_pushPtr;
  wire       [4:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [4:0]    pushCC_pushPtrGray;
  wire       [4:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_asyncAssertSyncDeassert;
  wire                system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized;
  reg        [4:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [4:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [4:0]    popCC_popPtrGray;
  wire       [4:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [3:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [3:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [3:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [3:0]    popCC_readPort_cmd_payload;
  wire       [31:0]   popCC_readPort_rsp_addr;
  wire       [3:0]    popCC_readPort_rsp_id;
  wire       [3:0]    popCC_readPort_rsp_region;
  wire       [7:0]    popCC_readPort_rsp_len;
  wire       [2:0]    popCC_readPort_rsp_size;
  wire       [1:0]    popCC_readPort_rsp_burst;
  wire       [0:0]    popCC_readPort_rsp_lock;
  wire       [3:0]    popCC_readPort_rsp_cache;
  wire       [3:0]    popCC_readPort_rsp_qos;
  wire       [2:0]    popCC_readPort_rsp_prot;
  wire       [64:0]   _zz_popCC_readPort_rsp_addr;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire       [31:0]   popCC_readArbitation_translated_payload_addr;
  wire       [3:0]    popCC_readArbitation_translated_payload_id;
  wire       [3:0]    popCC_readArbitation_translated_payload_region;
  wire       [7:0]    popCC_readArbitation_translated_payload_len;
  wire       [2:0]    popCC_readArbitation_translated_payload_size;
  wire       [1:0]    popCC_readArbitation_translated_payload_burst;
  wire       [0:0]    popCC_readArbitation_translated_payload_lock;
  wire       [3:0]    popCC_readArbitation_translated_payload_cache;
  wire       [3:0]    popCC_readArbitation_translated_payload_qos;
  wire       [2:0]    popCC_readArbitation_translated_payload_prot;
  wire                popCC_readArbitation_fire;
  reg        [4:0]    popCC_ptrToPush;
  reg        [4:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  reg [64:0] ram [0:15];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[3:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {io_push_payload_prot,{io_push_payload_qos,{io_push_payload_cache,{io_push_payload_lock,{io_push_payload_burst,{io_push_payload_size,{io_push_payload_len,{io_push_payload_region,{io_push_payload_id,io_push_payload_addr}}}}}}}}};
  always @(posedge io_ddrMasters_1_clk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_11 popToPushGray_buffercc (
    .io_dataIn             (popToPushGray[4:0]                    ), //i
    .io_dataOut            (popToPushGray_buffercc_io_dataOut[4:0]), //o
    .io_ddrMasters_1_clk   (io_ddrMasters_1_clk                   ), //i
    .io_ddrMasters_1_reset (io_ddrMasters_1_reset                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_12 system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn             (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut            (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_memoryClk          (io_memoryClk                                                                                                        ), //i
    .io_ddrMasters_1_reset (io_ddrMasters_1_reset                                                                                               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_13 pushToPopGray_buffercc (
    .io_dataIn                                                                             (pushToPopGray[4:0]                                                                   ), //i
    .io_dataOut                                                                            (pushToPopGray_buffercc_io_dataOut[4:0]                                               ), //o
    .io_memoryClk                                                                          (io_memoryClk                                                                         ), //i
    .system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized (system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 5'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[4 : 3] == (~ pushCC_popPtrGray[4 : 3])) && (pushCC_pushPtrGray[2 : 0] == pushCC_popPtrGray[2 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = pushCC_popPtrGray[4];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}});
  assign system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized = system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 5'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[3:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_addr = ram_spinal_port1;
  assign popCC_readPort_rsp_addr = _zz_popCC_readPort_rsp_addr[31 : 0];
  assign popCC_readPort_rsp_id = _zz_popCC_readPort_rsp_addr[35 : 32];
  assign popCC_readPort_rsp_region = _zz_popCC_readPort_rsp_addr[39 : 36];
  assign popCC_readPort_rsp_len = _zz_popCC_readPort_rsp_addr[47 : 40];
  assign popCC_readPort_rsp_size = _zz_popCC_readPort_rsp_addr[50 : 48];
  assign popCC_readPort_rsp_burst = _zz_popCC_readPort_rsp_addr[52 : 51];
  assign popCC_readPort_rsp_lock = _zz_popCC_readPort_rsp_addr[53 : 53];
  assign popCC_readPort_rsp_cache = _zz_popCC_readPort_rsp_addr[57 : 54];
  assign popCC_readPort_rsp_qos = _zz_popCC_readPort_rsp_addr[61 : 58];
  assign popCC_readPort_rsp_prot = _zz_popCC_readPort_rsp_addr[64 : 62];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_addr = popCC_readPort_rsp_addr;
  assign popCC_readArbitation_translated_payload_id = popCC_readPort_rsp_id;
  assign popCC_readArbitation_translated_payload_region = popCC_readPort_rsp_region;
  assign popCC_readArbitation_translated_payload_len = popCC_readPort_rsp_len;
  assign popCC_readArbitation_translated_payload_size = popCC_readPort_rsp_size;
  assign popCC_readArbitation_translated_payload_burst = popCC_readPort_rsp_burst;
  assign popCC_readArbitation_translated_payload_lock = popCC_readPort_rsp_lock;
  assign popCC_readArbitation_translated_payload_cache = popCC_readPort_rsp_cache;
  assign popCC_readArbitation_translated_payload_qos = popCC_readPort_rsp_qos;
  assign popCC_readArbitation_translated_payload_prot = popCC_readPort_rsp_prot;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_addr = popCC_readArbitation_translated_payload_addr;
  assign io_pop_payload_id = popCC_readArbitation_translated_payload_id;
  assign io_pop_payload_region = popCC_readArbitation_translated_payload_region;
  assign io_pop_payload_len = popCC_readArbitation_translated_payload_len;
  assign io_pop_payload_size = popCC_readArbitation_translated_payload_size;
  assign io_pop_payload_burst = popCC_readArbitation_translated_payload_burst;
  assign io_pop_payload_lock = popCC_readArbitation_translated_payload_lock;
  assign io_pop_payload_cache = popCC_readArbitation_translated_payload_cache;
  assign io_pop_payload_qos = popCC_readArbitation_translated_payload_qos;
  assign io_pop_payload_prot = popCC_readArbitation_translated_payload_prot;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = popCC_pushPtrGray[4];
  assign io_popOccupancy = ({_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  assign system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1 = system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized;
  always @(posedge io_ddrMasters_1_clk) begin
    if(io_ddrMasters_1_reset) begin
      pushCC_pushPtr <= 5'h0;
      pushCC_pushPtrGray <= 5'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized) begin
      popCC_popPtr <= 5'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 5'h0;
      popCC_ptrToOccupancy <= 5'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoLowLatency (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [1:0]    io_push_payload,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [1:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [1:0]    fifo_io_pop_payload;
  wire       [2:0]    fifo_io_occupancy;
  wire       [2:0]    fifo_io_availability;

  StreamFifo_3 fifo (
    .io_push_valid           (io_push_valid            ), //i
    .io_push_ready           (fifo_io_push_ready       ), //o
    .io_push_payload         (io_push_payload[1:0]     ), //i
    .io_pop_valid            (fifo_io_pop_valid        ), //o
    .io_pop_ready            (io_pop_ready             ), //i
    .io_pop_payload          (fifo_io_pop_payload[1:0] ), //o
    .io_flush                (io_flush                 ), //i
    .io_occupancy            (fifo_io_occupancy[2:0]   ), //o
    .io_availability         (fifo_io_availability[2:0]), //o
    .io_memoryClk            (io_memoryClk             ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset  )  //i
  );
  assign io_push_ready = fifo_io_push_ready;
  assign io_pop_valid = fifo_io_pop_valid;
  assign io_pop_payload = fifo_io_pop_payload;
  assign io_occupancy = fifo_io_occupancy;
  assign io_availability = fifo_io_availability;

endmodule

//StreamArbiter_8 replaced by StreamArbiter_7

module StreamArbiter_7 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [31:0]   io_inputs_0_payload_addr,
  input  wire [5:0]    io_inputs_0_payload_id,
  input  wire [3:0]    io_inputs_0_payload_region,
  input  wire [7:0]    io_inputs_0_payload_len,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire [1:0]    io_inputs_0_payload_burst,
  input  wire [0:0]    io_inputs_0_payload_lock,
  input  wire [3:0]    io_inputs_0_payload_cache,
  input  wire [3:0]    io_inputs_0_payload_qos,
  input  wire [2:0]    io_inputs_0_payload_prot,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [31:0]   io_inputs_1_payload_addr,
  input  wire [5:0]    io_inputs_1_payload_id,
  input  wire [3:0]    io_inputs_1_payload_region,
  input  wire [7:0]    io_inputs_1_payload_len,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire [1:0]    io_inputs_1_payload_burst,
  input  wire [0:0]    io_inputs_1_payload_lock,
  input  wire [3:0]    io_inputs_1_payload_cache,
  input  wire [3:0]    io_inputs_1_payload_qos,
  input  wire [2:0]    io_inputs_1_payload_prot,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [31:0]   io_inputs_2_payload_addr,
  input  wire [5:0]    io_inputs_2_payload_id,
  input  wire [3:0]    io_inputs_2_payload_region,
  input  wire [7:0]    io_inputs_2_payload_len,
  input  wire [2:0]    io_inputs_2_payload_size,
  input  wire [1:0]    io_inputs_2_payload_burst,
  input  wire [0:0]    io_inputs_2_payload_lock,
  input  wire [3:0]    io_inputs_2_payload_cache,
  input  wire [3:0]    io_inputs_2_payload_qos,
  input  wire [2:0]    io_inputs_2_payload_prot,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [31:0]   io_output_payload_addr,
  output wire [5:0]    io_output_payload_id,
  output wire [3:0]    io_output_payload_region,
  output wire [7:0]    io_output_payload_len,
  output wire [2:0]    io_output_payload_size,
  output wire [1:0]    io_output_payload_burst,
  output wire [0:0]    io_output_payload_lock,
  output wire [3:0]    io_output_payload_cache,
  output wire [3:0]    io_output_payload_qos,
  output wire [2:0]    io_output_payload_prot,
  output wire [1:0]    io_chosen,
  output wire [2:0]    io_chosenOH,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire       [5:0]    _zz__zz_maskProposal_0_2;
  wire       [5:0]    _zz__zz_maskProposal_0_2_1;
  wire       [2:0]    _zz__zz_maskProposal_0_2_2;
  reg        [31:0]   _zz_io_output_payload_addr_1;
  reg        [5:0]    _zz_io_output_payload_id;
  reg        [3:0]    _zz_io_output_payload_region;
  reg        [7:0]    _zz_io_output_payload_len;
  reg        [2:0]    _zz_io_output_payload_size;
  reg        [1:0]    _zz_io_output_payload_burst;
  reg        [0:0]    _zz_io_output_payload_lock;
  reg        [3:0]    _zz_io_output_payload_cache;
  reg        [3:0]    _zz_io_output_payload_qos;
  reg        [2:0]    _zz_io_output_payload_prot;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire       [2:0]    _zz_maskProposal_0;
  wire       [5:0]    _zz_maskProposal_0_1;
  wire       [5:0]    _zz_maskProposal_0_2;
  wire       [2:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire       [1:0]    _zz_io_output_payload_addr;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_1,{maskLocked_0,maskLocked_2}};
  assign _zz__zz_maskProposal_0_2_1 = {3'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(_zz_io_output_payload_addr)
      2'b00 : begin
        _zz_io_output_payload_addr_1 = io_inputs_0_payload_addr;
        _zz_io_output_payload_id = io_inputs_0_payload_id;
        _zz_io_output_payload_region = io_inputs_0_payload_region;
        _zz_io_output_payload_len = io_inputs_0_payload_len;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_burst = io_inputs_0_payload_burst;
        _zz_io_output_payload_lock = io_inputs_0_payload_lock;
        _zz_io_output_payload_cache = io_inputs_0_payload_cache;
        _zz_io_output_payload_qos = io_inputs_0_payload_qos;
        _zz_io_output_payload_prot = io_inputs_0_payload_prot;
      end
      2'b01 : begin
        _zz_io_output_payload_addr_1 = io_inputs_1_payload_addr;
        _zz_io_output_payload_id = io_inputs_1_payload_id;
        _zz_io_output_payload_region = io_inputs_1_payload_region;
        _zz_io_output_payload_len = io_inputs_1_payload_len;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_burst = io_inputs_1_payload_burst;
        _zz_io_output_payload_lock = io_inputs_1_payload_lock;
        _zz_io_output_payload_cache = io_inputs_1_payload_cache;
        _zz_io_output_payload_qos = io_inputs_1_payload_qos;
        _zz_io_output_payload_prot = io_inputs_1_payload_prot;
      end
      default : begin
        _zz_io_output_payload_addr_1 = io_inputs_2_payload_addr;
        _zz_io_output_payload_id = io_inputs_2_payload_id;
        _zz_io_output_payload_region = io_inputs_2_payload_region;
        _zz_io_output_payload_len = io_inputs_2_payload_len;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_burst = io_inputs_2_payload_burst;
        _zz_io_output_payload_lock = io_inputs_2_payload_lock;
        _zz_io_output_payload_cache = io_inputs_2_payload_cache;
        _zz_io_output_payload_qos = io_inputs_2_payload_qos;
        _zz_io_output_payload_prot = io_inputs_2_payload_prot;
      end
    endcase
  end

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign _zz_maskProposal_0 = {io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[5 : 3] | _zz_maskProposal_0_2[2 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = (((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2));
  assign _zz_io_output_payload_addr = {maskRouted_2,maskRouted_1};
  assign io_output_payload_addr = _zz_io_output_payload_addr_1;
  assign io_output_payload_id = _zz_io_output_payload_id;
  assign io_output_payload_region = _zz_io_output_payload_region;
  assign io_output_payload_len = _zz_io_output_payload_len;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_burst = _zz_io_output_payload_burst;
  assign io_output_payload_lock = _zz_io_output_payload_lock;
  assign io_output_payload_cache = _zz_io_output_payload_cache;
  assign io_output_payload_qos = _zz_io_output_payload_qos;
  assign io_output_payload_prot = _zz_io_output_payload_prot;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_chosenOH = {maskRouted_2,{maskRouted_1,maskRouted_0}};
  assign _zz_io_chosen = io_chosenOH[1];
  assign _zz_io_chosen_1 = io_chosenOH[2];
  assign io_chosen = {_zz_io_chosen_1,_zz_io_chosen};
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamFifoCC_1 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire          io_push_payload_last,
  input  wire [1:0]    io_push_payload_fragment_source,
  input  wire [0:0]    io_push_payload_fragment_opcode,
  input  wire [127:0]  io_push_payload_fragment_data,
  input  wire [45:0]   io_push_payload_fragment_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire          io_pop_payload_last,
  output wire [1:0]    io_pop_payload_fragment_source,
  output wire [0:0]    io_pop_payload_fragment_opcode,
  output wire [127:0]  io_pop_payload_fragment_data,
  output wire [45:0]   io_pop_payload_fragment_context,
  output wire [6:0]    io_pushOccupancy,
  output wire [6:0]    io_popOccupancy,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset,
  input  wire          io_systemClk
);

  reg        [177:0]  ram_spinal_port1;
  wire       [6:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [6:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [6:0]    _zz_pushCC_pushPtrGray;
  wire       [5:0]    _zz_ram_port;
  wire       [177:0]  _zz_ram_port_1;
  wire       [6:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [6:0]    popToPushGray;
  wire       [6:0]    pushToPopGray;
  reg        [6:0]    pushCC_pushPtr;
  wire       [6:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [6:0]    pushCC_pushPtrGray;
  wire       [6:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                _zz_io_pushOccupancy_4;
  wire                _zz_io_pushOccupancy_5;
  wire                system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_synchronized;
  reg        [6:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [6:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [6:0]    popCC_popPtrGray;
  wire       [6:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [5:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [5:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [5:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [5:0]    popCC_readPort_cmd_payload;
  wire                popCC_readPort_rsp_last;
  wire       [1:0]    popCC_readPort_rsp_fragment_source;
  wire       [0:0]    popCC_readPort_rsp_fragment_opcode;
  wire       [127:0]  popCC_readPort_rsp_fragment_data;
  wire       [45:0]   popCC_readPort_rsp_fragment_context;
  wire       [177:0]  _zz_popCC_readPort_rsp_last;
  wire       [176:0]  _zz_popCC_readPort_rsp_fragment_source;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire                popCC_readArbitation_translated_payload_last;
  wire       [1:0]    popCC_readArbitation_translated_payload_fragment_source;
  wire       [0:0]    popCC_readArbitation_translated_payload_fragment_opcode;
  wire       [127:0]  popCC_readArbitation_translated_payload_fragment_data;
  wire       [45:0]   popCC_readArbitation_translated_payload_fragment_context;
  wire                popCC_readArbitation_fire;
  reg        [6:0]    popCC_ptrToPush;
  reg        [6:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  wire                _zz_io_popOccupancy_4;
  wire                _zz_io_popOccupancy_5;
  reg [177:0] ram [0:63];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[5:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {{io_push_payload_fragment_context,{io_push_payload_fragment_data,{io_push_payload_fragment_opcode,io_push_payload_fragment_source}}},io_push_payload_last};
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_systemClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_8 popToPushGray_buffercc (
    .io_dataIn               (popToPushGray[6:0]                    ), //i
    .io_dataOut              (popToPushGray_buffercc_io_dataOut[6:0]), //o
    .io_memoryClk            (io_memoryClk                          ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset               )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_9 system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn               (system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut              (system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_systemClk            (io_systemClk                                                                                            ), //i
    .ddrCd_logic_outputReset (ddrCd_logic_outputReset                                                                                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_10 pushToPopGray_buffercc (
    .io_dataIn                                                                 (pushToPopGray[6:0]                                                       ), //i
    .io_dataOut                                                                (pushToPopGray_buffercc_io_dataOut[6:0]                                   ), //o
    .io_systemClk                                                              (io_systemClk                                                             ), //i
    .system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_synchronized (system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 7'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[6 : 5] == (~ pushCC_popPtrGray[6 : 5])) && (pushCC_pushPtrGray[4 : 0] == pushCC_popPtrGray[4 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = (pushCC_popPtrGray[4] ^ _zz_io_pushOccupancy_4);
  assign _zz_io_pushOccupancy_4 = (pushCC_popPtrGray[5] ^ _zz_io_pushOccupancy_5);
  assign _zz_io_pushOccupancy_5 = pushCC_popPtrGray[6];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_5,{_zz_io_pushOccupancy_4,{_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}}}});
  assign system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_synchronized = system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 7'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[5:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_last = ram_spinal_port1;
  assign _zz_popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_last[177 : 1];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_last[0];
  assign popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_fragment_source[1 : 0];
  assign popCC_readPort_rsp_fragment_opcode = _zz_popCC_readPort_rsp_fragment_source[2 : 2];
  assign popCC_readPort_rsp_fragment_data = _zz_popCC_readPort_rsp_fragment_source[130 : 3];
  assign popCC_readPort_rsp_fragment_context = _zz_popCC_readPort_rsp_fragment_source[176 : 131];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign popCC_readArbitation_translated_payload_fragment_source = popCC_readPort_rsp_fragment_source;
  assign popCC_readArbitation_translated_payload_fragment_opcode = popCC_readPort_rsp_fragment_opcode;
  assign popCC_readArbitation_translated_payload_fragment_data = popCC_readPort_rsp_fragment_data;
  assign popCC_readArbitation_translated_payload_fragment_context = popCC_readPort_rsp_fragment_context;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign io_pop_payload_fragment_source = popCC_readArbitation_translated_payload_fragment_source;
  assign io_pop_payload_fragment_opcode = popCC_readArbitation_translated_payload_fragment_opcode;
  assign io_pop_payload_fragment_data = popCC_readArbitation_translated_payload_fragment_data;
  assign io_pop_payload_fragment_context = popCC_readArbitation_translated_payload_fragment_context;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = (popCC_pushPtrGray[4] ^ _zz_io_popOccupancy_4);
  assign _zz_io_popOccupancy_4 = (popCC_pushPtrGray[5] ^ _zz_io_popOccupancy_5);
  assign _zz_io_popOccupancy_5 = popCC_pushPtrGray[6];
  assign io_popOccupancy = ({_zz_io_popOccupancy_5,{_zz_io_popOccupancy_4,{_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      pushCC_pushPtr <= 7'h0;
      pushCC_pushPtrGray <= 7'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_synchronized) begin
      popCC_popPtr <= 7'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 7'h0;
      popCC_ptrToOccupancy <= 7'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

module StreamFifoCC (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire          io_push_payload_last,
  input  wire [1:0]    io_push_payload_fragment_source,
  input  wire [0:0]    io_push_payload_fragment_opcode,
  input  wire [31:0]   io_push_payload_fragment_address,
  input  wire [5:0]    io_push_payload_fragment_length,
  input  wire [127:0]  io_push_payload_fragment_data,
  input  wire [15:0]   io_push_payload_fragment_mask,
  input  wire [45:0]   io_push_payload_fragment_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire          io_pop_payload_last,
  output wire [1:0]    io_pop_payload_fragment_source,
  output wire [0:0]    io_pop_payload_fragment_opcode,
  output wire [31:0]   io_pop_payload_fragment_address,
  output wire [5:0]    io_pop_payload_fragment_length,
  output wire [127:0]  io_pop_payload_fragment_data,
  output wire [15:0]   io_pop_payload_fragment_mask,
  output wire [45:0]   io_pop_payload_fragment_context,
  output wire [6:0]    io_pushOccupancy,
  output wire [6:0]    io_popOccupancy,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset,
  input  wire          io_memoryClk
);

  reg        [231:0]  ram_spinal_port1;
  wire       [6:0]    popToPushGray_buffercc_io_dataOut;
  wire                system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire       [6:0]    pushToPopGray_buffercc_io_dataOut;
  wire       [6:0]    _zz_pushCC_pushPtrGray;
  wire       [5:0]    _zz_ram_port;
  wire       [231:0]  _zz_ram_port_1;
  wire       [6:0]    _zz_popCC_popPtrGray;
  reg                 _zz_1;
  wire       [6:0]    popToPushGray;
  wire       [6:0]    pushToPopGray;
  reg        [6:0]    pushCC_pushPtr;
  wire       [6:0]    pushCC_pushPtrPlus;
  wire                io_push_fire;
  reg        [6:0]    pushCC_pushPtrGray;
  wire       [6:0]    pushCC_popPtrGray;
  wire                pushCC_full;
  wire                _zz_io_pushOccupancy;
  wire                _zz_io_pushOccupancy_1;
  wire                _zz_io_pushOccupancy_2;
  wire                _zz_io_pushOccupancy_3;
  wire                _zz_io_pushOccupancy_4;
  wire                _zz_io_pushOccupancy_5;
  wire                system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_synchronized;
  reg        [6:0]    popCC_popPtr;
  (* keep , syn_keep *) wire       [6:0]    popCC_popPtrPlus /* synthesis syn_keep = 1 */ ;
  wire       [6:0]    popCC_popPtrGray;
  wire       [6:0]    popCC_pushPtrGray;
  wire                popCC_addressGen_valid;
  reg                 popCC_addressGen_ready;
  wire       [5:0]    popCC_addressGen_payload;
  wire                popCC_empty;
  wire                popCC_addressGen_fire;
  wire                popCC_readArbitation_valid;
  wire                popCC_readArbitation_ready;
  wire       [5:0]    popCC_readArbitation_payload;
  reg                 popCC_addressGen_rValid;
  reg        [5:0]    popCC_addressGen_rData;
  wire                when_Stream_l375;
  wire                popCC_readPort_cmd_valid;
  wire       [5:0]    popCC_readPort_cmd_payload;
  wire                popCC_readPort_rsp_last;
  wire       [1:0]    popCC_readPort_rsp_fragment_source;
  wire       [0:0]    popCC_readPort_rsp_fragment_opcode;
  wire       [31:0]   popCC_readPort_rsp_fragment_address;
  wire       [5:0]    popCC_readPort_rsp_fragment_length;
  wire       [127:0]  popCC_readPort_rsp_fragment_data;
  wire       [15:0]   popCC_readPort_rsp_fragment_mask;
  wire       [45:0]   popCC_readPort_rsp_fragment_context;
  wire       [231:0]  _zz_popCC_readPort_rsp_last;
  wire       [230:0]  _zz_popCC_readPort_rsp_fragment_source;
  wire                popCC_readArbitation_translated_valid;
  wire                popCC_readArbitation_translated_ready;
  wire                popCC_readArbitation_translated_payload_last;
  wire       [1:0]    popCC_readArbitation_translated_payload_fragment_source;
  wire       [0:0]    popCC_readArbitation_translated_payload_fragment_opcode;
  wire       [31:0]   popCC_readArbitation_translated_payload_fragment_address;
  wire       [5:0]    popCC_readArbitation_translated_payload_fragment_length;
  wire       [127:0]  popCC_readArbitation_translated_payload_fragment_data;
  wire       [15:0]   popCC_readArbitation_translated_payload_fragment_mask;
  wire       [45:0]   popCC_readArbitation_translated_payload_fragment_context;
  wire                popCC_readArbitation_fire;
  reg        [6:0]    popCC_ptrToPush;
  reg        [6:0]    popCC_ptrToOccupancy;
  wire                _zz_io_popOccupancy;
  wire                _zz_io_popOccupancy_1;
  wire                _zz_io_popOccupancy_2;
  wire                _zz_io_popOccupancy_3;
  wire                _zz_io_popOccupancy_4;
  wire                _zz_io_popOccupancy_5;
  reg [231:0] ram [0:63];

  assign _zz_pushCC_pushPtrGray = (pushCC_pushPtrPlus >>> 1'b1);
  assign _zz_ram_port = pushCC_pushPtr[5:0];
  assign _zz_popCC_popPtrGray = (popCC_popPtr >>> 1'b1);
  assign _zz_ram_port_1 = {{io_push_payload_fragment_context,{io_push_payload_fragment_mask,{io_push_payload_fragment_data,{io_push_payload_fragment_length,{io_push_payload_fragment_address,{io_push_payload_fragment_opcode,io_push_payload_fragment_source}}}}}},io_push_payload_last};
  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      ram[_zz_ram_port] <= _zz_ram_port_1;
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_readPort_cmd_valid) begin
      ram_spinal_port1 <= ram[popCC_readPort_cmd_payload];
    end
  end

  (* keep_hierarchy = "TRUE" *) BufferCC_5 popToPushGray_buffercc (
    .io_dataIn                  (popToPushGray[6:0]                    ), //i
    .io_dataOut                 (popToPushGray_buffercc_io_dataOut[6:0]), //o
    .io_systemClk               (io_systemClk                          ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset            )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_6 system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn                  (system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut                 (system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .io_memoryClk               (io_memoryClk                                                                                               ), //i
    .systemCd_logic_outputReset (systemCd_logic_outputReset                                                                                 )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_7 pushToPopGray_buffercc (
    .io_dataIn                                                                    (pushToPopGray[6:0]                                                          ), //i
    .io_dataOut                                                                   (pushToPopGray_buffercc_io_dataOut[6:0]                                      ), //o
    .io_memoryClk                                                                 (io_memoryClk                                                                ), //i
    .system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_synchronized (system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_synchronized)  //i
  );
  always @(*) begin
    _zz_1 = 1'b0;
    if(io_push_fire) begin
      _zz_1 = 1'b1;
    end
  end

  assign pushCC_pushPtrPlus = (pushCC_pushPtr + 7'h01);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign pushCC_popPtrGray = popToPushGray_buffercc_io_dataOut;
  assign pushCC_full = ((pushCC_pushPtrGray[6 : 5] == (~ pushCC_popPtrGray[6 : 5])) && (pushCC_pushPtrGray[4 : 0] == pushCC_popPtrGray[4 : 0]));
  assign io_push_ready = (! pushCC_full);
  assign _zz_io_pushOccupancy = (pushCC_popPtrGray[1] ^ _zz_io_pushOccupancy_1);
  assign _zz_io_pushOccupancy_1 = (pushCC_popPtrGray[2] ^ _zz_io_pushOccupancy_2);
  assign _zz_io_pushOccupancy_2 = (pushCC_popPtrGray[3] ^ _zz_io_pushOccupancy_3);
  assign _zz_io_pushOccupancy_3 = (pushCC_popPtrGray[4] ^ _zz_io_pushOccupancy_4);
  assign _zz_io_pushOccupancy_4 = (pushCC_popPtrGray[5] ^ _zz_io_pushOccupancy_5);
  assign _zz_io_pushOccupancy_5 = pushCC_popPtrGray[6];
  assign io_pushOccupancy = (pushCC_pushPtr - {_zz_io_pushOccupancy_5,{_zz_io_pushOccupancy_4,{_zz_io_pushOccupancy_3,{_zz_io_pushOccupancy_2,{_zz_io_pushOccupancy_1,{_zz_io_pushOccupancy,(pushCC_popPtrGray[0] ^ _zz_io_pushOccupancy)}}}}}});
  assign system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_synchronized = system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign popCC_popPtrPlus = (popCC_popPtr + 7'h01);
  assign popCC_popPtrGray = (_zz_popCC_popPtrGray ^ popCC_popPtr);
  assign popCC_pushPtrGray = pushToPopGray_buffercc_io_dataOut;
  assign popCC_empty = (popCC_popPtrGray == popCC_pushPtrGray);
  assign popCC_addressGen_valid = (! popCC_empty);
  assign popCC_addressGen_payload = popCC_popPtr[5:0];
  assign popCC_addressGen_fire = (popCC_addressGen_valid && popCC_addressGen_ready);
  always @(*) begin
    popCC_addressGen_ready = popCC_readArbitation_ready;
    if(when_Stream_l375) begin
      popCC_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! popCC_readArbitation_valid);
  assign popCC_readArbitation_valid = popCC_addressGen_rValid;
  assign popCC_readArbitation_payload = popCC_addressGen_rData;
  assign _zz_popCC_readPort_rsp_last = ram_spinal_port1;
  assign _zz_popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_last[231 : 1];
  assign popCC_readPort_rsp_last = _zz_popCC_readPort_rsp_last[0];
  assign popCC_readPort_rsp_fragment_source = _zz_popCC_readPort_rsp_fragment_source[1 : 0];
  assign popCC_readPort_rsp_fragment_opcode = _zz_popCC_readPort_rsp_fragment_source[2 : 2];
  assign popCC_readPort_rsp_fragment_address = _zz_popCC_readPort_rsp_fragment_source[34 : 3];
  assign popCC_readPort_rsp_fragment_length = _zz_popCC_readPort_rsp_fragment_source[40 : 35];
  assign popCC_readPort_rsp_fragment_data = _zz_popCC_readPort_rsp_fragment_source[168 : 41];
  assign popCC_readPort_rsp_fragment_mask = _zz_popCC_readPort_rsp_fragment_source[184 : 169];
  assign popCC_readPort_rsp_fragment_context = _zz_popCC_readPort_rsp_fragment_source[230 : 185];
  assign popCC_readPort_cmd_valid = popCC_addressGen_fire;
  assign popCC_readPort_cmd_payload = popCC_addressGen_payload;
  assign popCC_readArbitation_translated_valid = popCC_readArbitation_valid;
  assign popCC_readArbitation_ready = popCC_readArbitation_translated_ready;
  assign popCC_readArbitation_translated_payload_last = popCC_readPort_rsp_last;
  assign popCC_readArbitation_translated_payload_fragment_source = popCC_readPort_rsp_fragment_source;
  assign popCC_readArbitation_translated_payload_fragment_opcode = popCC_readPort_rsp_fragment_opcode;
  assign popCC_readArbitation_translated_payload_fragment_address = popCC_readPort_rsp_fragment_address;
  assign popCC_readArbitation_translated_payload_fragment_length = popCC_readPort_rsp_fragment_length;
  assign popCC_readArbitation_translated_payload_fragment_data = popCC_readPort_rsp_fragment_data;
  assign popCC_readArbitation_translated_payload_fragment_mask = popCC_readPort_rsp_fragment_mask;
  assign popCC_readArbitation_translated_payload_fragment_context = popCC_readPort_rsp_fragment_context;
  assign io_pop_valid = popCC_readArbitation_translated_valid;
  assign popCC_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_last = popCC_readArbitation_translated_payload_last;
  assign io_pop_payload_fragment_source = popCC_readArbitation_translated_payload_fragment_source;
  assign io_pop_payload_fragment_opcode = popCC_readArbitation_translated_payload_fragment_opcode;
  assign io_pop_payload_fragment_address = popCC_readArbitation_translated_payload_fragment_address;
  assign io_pop_payload_fragment_length = popCC_readArbitation_translated_payload_fragment_length;
  assign io_pop_payload_fragment_data = popCC_readArbitation_translated_payload_fragment_data;
  assign io_pop_payload_fragment_mask = popCC_readArbitation_translated_payload_fragment_mask;
  assign io_pop_payload_fragment_context = popCC_readArbitation_translated_payload_fragment_context;
  assign popCC_readArbitation_fire = (popCC_readArbitation_valid && popCC_readArbitation_ready);
  assign _zz_io_popOccupancy = (popCC_pushPtrGray[1] ^ _zz_io_popOccupancy_1);
  assign _zz_io_popOccupancy_1 = (popCC_pushPtrGray[2] ^ _zz_io_popOccupancy_2);
  assign _zz_io_popOccupancy_2 = (popCC_pushPtrGray[3] ^ _zz_io_popOccupancy_3);
  assign _zz_io_popOccupancy_3 = (popCC_pushPtrGray[4] ^ _zz_io_popOccupancy_4);
  assign _zz_io_popOccupancy_4 = (popCC_pushPtrGray[5] ^ _zz_io_popOccupancy_5);
  assign _zz_io_popOccupancy_5 = popCC_pushPtrGray[6];
  assign io_popOccupancy = ({_zz_io_popOccupancy_5,{_zz_io_popOccupancy_4,{_zz_io_popOccupancy_3,{_zz_io_popOccupancy_2,{_zz_io_popOccupancy_1,{_zz_io_popOccupancy,(popCC_pushPtrGray[0] ^ _zz_io_popOccupancy)}}}}}} - popCC_ptrToOccupancy);
  assign pushToPopGray = pushCC_pushPtrGray;
  assign popToPushGray = popCC_ptrToPush;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      pushCC_pushPtr <= 7'h0;
      pushCC_pushPtrGray <= 7'h0;
    end else begin
      if(io_push_fire) begin
        pushCC_pushPtrGray <= (_zz_pushCC_pushPtrGray ^ pushCC_pushPtrPlus);
      end
      if(io_push_fire) begin
        pushCC_pushPtr <= pushCC_pushPtrPlus;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_synchronized) begin
      popCC_popPtr <= 7'h0;
      popCC_addressGen_rValid <= 1'b0;
      popCC_ptrToPush <= 7'h0;
      popCC_ptrToOccupancy <= 7'h0;
    end else begin
      if(popCC_addressGen_fire) begin
        popCC_popPtr <= popCC_popPtrPlus;
      end
      if(popCC_addressGen_ready) begin
        popCC_addressGen_rValid <= popCC_addressGen_valid;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToPush <= popCC_popPtrGray;
      end
      if(popCC_readArbitation_fire) begin
        popCC_ptrToOccupancy <= popCC_popPtr;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(popCC_addressGen_ready) begin
      popCC_addressGen_rData <= popCC_addressGen_payload;
    end
  end


endmodule

//StreamFifo_2 replaced by StreamFifo_1

module StreamFifo_1 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [1:0]    io_push_payload_source,
  input  wire [45:0]   io_push_payload_context,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [1:0]    io_pop_payload_source,
  output wire [45:0]   io_pop_payload_context,
  input  wire          io_flush,
  output wire [6:0]    io_occupancy,
  output wire [6:0]    io_availability,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  reg        [47:0]   logic_ram_spinal_port1;
  wire       [47:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [6:0]    logic_ptr_push;
  reg        [6:0]    logic_ptr_pop;
  wire       [6:0]    logic_ptr_occupancy;
  wire       [6:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [5:0]    logic_push_onRam_write_payload_address;
  wire       [1:0]    logic_push_onRam_write_payload_data_source;
  wire       [45:0]   logic_push_onRam_write_payload_data_context;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [5:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [5:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [5:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [5:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [1:0]    logic_pop_sync_readPort_rsp_source;
  wire       [45:0]   logic_pop_sync_readPort_rsp_context;
  wire       [47:0]   _zz_logic_pop_sync_readPort_rsp_source;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [1:0]    logic_pop_sync_readArbitation_translated_payload_source;
  wire       [45:0]   logic_pop_sync_readArbitation_translated_payload_context;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [6:0]    logic_pop_sync_popReg;
  reg [47:0] logic_ram [0:63];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_context,logic_push_onRam_write_payload_data_source};
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge io_memoryClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 7'h40) == 7'h0);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[5:0];
  assign logic_push_onRam_write_payload_data_source = io_push_payload_source;
  assign logic_push_onRam_write_payload_data_context = io_push_payload_context;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[5:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_source = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_source = _zz_logic_pop_sync_readPort_rsp_source[1 : 0];
  assign logic_pop_sync_readPort_rsp_context = _zz_logic_pop_sync_readPort_rsp_source[47 : 2];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_source = logic_pop_sync_readPort_rsp_source;
  assign logic_pop_sync_readArbitation_translated_payload_context = logic_pop_sync_readPort_rsp_context;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_source = logic_pop_sync_readArbitation_translated_payload_source;
  assign io_pop_payload_context = logic_pop_sync_readArbitation_translated_payload_context;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (7'h40 - logic_ptr_occupancy);
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      logic_ptr_push <= 7'h0;
      logic_ptr_pop <= 7'h0;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 7'h0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 7'h01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 7'h01);
      end
      if(io_flush) begin
        logic_ptr_push <= 7'h0;
        logic_ptr_pop <= 7'h0;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 7'h0;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module StreamArbiter_6 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire          io_inputs_0_payload_last,
  input  wire [1:0]    io_inputs_0_payload_fragment_source,
  input  wire [0:0]    io_inputs_0_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_0_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_payload_fragment_length,
  input  wire [63:0]   io_inputs_0_payload_fragment_data,
  input  wire [7:0]    io_inputs_0_payload_fragment_mask,
  input  wire [43:0]   io_inputs_0_payload_fragment_context,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire          io_inputs_1_payload_last,
  input  wire [1:0]    io_inputs_1_payload_fragment_source,
  input  wire [0:0]    io_inputs_1_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_1_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_payload_fragment_length,
  input  wire [63:0]   io_inputs_1_payload_fragment_data,
  input  wire [7:0]    io_inputs_1_payload_fragment_mask,
  input  wire [43:0]   io_inputs_1_payload_fragment_context,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [1:0]    io_output_payload_fragment_source,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire [31:0]   io_output_payload_fragment_address,
  output wire [5:0]    io_output_payload_fragment_length,
  output wire [63:0]   io_output_payload_fragment_data,
  output wire [7:0]    io_output_payload_fragment_mask,
  output wire [43:0]   io_output_payload_fragment_context,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                when_Stream_l683;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l683 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_output_payload_fragment_source = (maskRouted_0 ? io_inputs_0_payload_fragment_source : io_inputs_1_payload_fragment_source);
  assign io_output_payload_fragment_opcode = (maskRouted_0 ? io_inputs_0_payload_fragment_opcode : io_inputs_1_payload_fragment_opcode);
  assign io_output_payload_fragment_address = (maskRouted_0 ? io_inputs_0_payload_fragment_address : io_inputs_1_payload_fragment_address);
  assign io_output_payload_fragment_length = (maskRouted_0 ? io_inputs_0_payload_fragment_length : io_inputs_1_payload_fragment_length);
  assign io_output_payload_fragment_data = (maskRouted_0 ? io_inputs_0_payload_fragment_data : io_inputs_1_payload_fragment_data);
  assign io_output_payload_fragment_mask = (maskRouted_0 ? io_inputs_0_payload_fragment_mask : io_inputs_1_payload_fragment_mask);
  assign io_output_payload_fragment_context = (maskRouted_0 ? io_inputs_0_payload_fragment_context : io_inputs_1_payload_fragment_context);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l683) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamFork_2 (
  input  wire          io_input_valid,
  output reg           io_input_ready,
  input  wire          io_input_payload_all,
  input  wire [31:0]   io_input_payload_address,
  input  wire [5:0]    io_input_payload_length,
  input  wire [0:0]    io_input_payload_source,
  output wire          io_outputs_0_valid,
  input  wire          io_outputs_0_ready,
  output wire          io_outputs_0_payload_all,
  output wire [31:0]   io_outputs_0_payload_address,
  output wire [5:0]    io_outputs_0_payload_length,
  output wire [0:0]    io_outputs_0_payload_source,
  output wire          io_outputs_1_valid,
  input  wire          io_outputs_1_ready,
  output wire          io_outputs_1_payload_all,
  output wire [31:0]   io_outputs_1_payload_address,
  output wire [5:0]    io_outputs_1_payload_length,
  output wire [0:0]    io_outputs_1_payload_source,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg                 logic_linkEnable_0;
  reg                 logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                io_outputs_0_fire;
  wire                io_outputs_1_fire;

  always @(*) begin
    io_input_ready = 1'b1;
    if(when_Stream_l1063) begin
      io_input_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      io_input_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! io_outputs_0_ready) && logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! io_outputs_1_ready) && logic_linkEnable_1);
  assign io_outputs_0_valid = (io_input_valid && logic_linkEnable_0);
  assign io_outputs_0_payload_all = io_input_payload_all;
  assign io_outputs_0_payload_address = io_input_payload_address;
  assign io_outputs_0_payload_length = io_input_payload_length;
  assign io_outputs_0_payload_source = io_input_payload_source;
  assign io_outputs_0_fire = (io_outputs_0_valid && io_outputs_0_ready);
  assign io_outputs_1_valid = (io_input_valid && logic_linkEnable_1);
  assign io_outputs_1_payload_all = io_input_payload_all;
  assign io_outputs_1_payload_address = io_input_payload_address;
  assign io_outputs_1_payload_length = io_input_payload_length;
  assign io_outputs_1_payload_source = io_input_payload_source;
  assign io_outputs_1_fire = (io_outputs_1_valid && io_outputs_1_ready);
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      logic_linkEnable_0 <= 1'b1;
      logic_linkEnable_1 <= 1'b1;
    end else begin
      if(io_outputs_0_fire) begin
        logic_linkEnable_0 <= 1'b0;
      end
      if(io_outputs_1_fire) begin
        logic_linkEnable_1 <= 1'b0;
      end
      if(io_input_ready) begin
        logic_linkEnable_0 <= 1'b1;
        logic_linkEnable_1 <= 1'b1;
      end
    end
  end


endmodule

module StreamArbiter_5 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire          io_inputs_0_payload_last,
  input  wire [0:0]    io_inputs_0_payload_fragment_source,
  input  wire [0:0]    io_inputs_0_payload_fragment_opcode,
  input  wire          io_inputs_0_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_0_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_payload_fragment_length,
  input  wire [63:0]   io_inputs_0_payload_fragment_data,
  input  wire [7:0]    io_inputs_0_payload_fragment_mask,
  input  wire [3:0]    io_inputs_0_payload_fragment_context,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire          io_inputs_1_payload_last,
  input  wire [0:0]    io_inputs_1_payload_fragment_source,
  input  wire [0:0]    io_inputs_1_payload_fragment_opcode,
  input  wire          io_inputs_1_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_1_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_payload_fragment_length,
  input  wire [63:0]   io_inputs_1_payload_fragment_data,
  input  wire [7:0]    io_inputs_1_payload_fragment_mask,
  input  wire [3:0]    io_inputs_1_payload_fragment_context,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [0:0]    io_output_payload_fragment_source,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire          io_output_payload_fragment_exclusive,
  output wire [31:0]   io_output_payload_fragment_address,
  output wire [5:0]    io_output_payload_fragment_length,
  output wire [63:0]   io_output_payload_fragment_data,
  output wire [7:0]    io_output_payload_fragment_mask,
  output wire [3:0]    io_output_payload_fragment_context,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                when_Stream_l683;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l683 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_output_payload_fragment_source = (maskRouted_0 ? io_inputs_0_payload_fragment_source : io_inputs_1_payload_fragment_source);
  assign io_output_payload_fragment_opcode = (maskRouted_0 ? io_inputs_0_payload_fragment_opcode : io_inputs_1_payload_fragment_opcode);
  assign io_output_payload_fragment_exclusive = (maskRouted_0 ? io_inputs_0_payload_fragment_exclusive : io_inputs_1_payload_fragment_exclusive);
  assign io_output_payload_fragment_address = (maskRouted_0 ? io_inputs_0_payload_fragment_address : io_inputs_1_payload_fragment_address);
  assign io_output_payload_fragment_length = (maskRouted_0 ? io_inputs_0_payload_fragment_length : io_inputs_1_payload_fragment_length);
  assign io_output_payload_fragment_data = (maskRouted_0 ? io_inputs_0_payload_fragment_data : io_inputs_1_payload_fragment_data);
  assign io_output_payload_fragment_mask = (maskRouted_0 ? io_inputs_0_payload_fragment_mask : io_inputs_1_payload_fragment_mask);
  assign io_output_payload_fragment_context = (maskRouted_0 ? io_inputs_0_payload_fragment_context : io_inputs_1_payload_fragment_context);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l683) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamArbiter_4 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire          io_inputs_0_payload_last,
  input  wire [0:0]    io_inputs_0_payload_fragment_source,
  input  wire [0:0]    io_inputs_0_payload_fragment_opcode,
  input  wire          io_inputs_0_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_0_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_payload_fragment_length,
  input  wire [3:0]    io_inputs_0_payload_fragment_context,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire          io_inputs_1_payload_last,
  input  wire [0:0]    io_inputs_1_payload_fragment_source,
  input  wire [0:0]    io_inputs_1_payload_fragment_opcode,
  input  wire          io_inputs_1_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_1_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_payload_fragment_length,
  input  wire [3:0]    io_inputs_1_payload_fragment_context,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [0:0]    io_output_payload_fragment_source,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire          io_output_payload_fragment_exclusive,
  output wire [31:0]   io_output_payload_fragment_address,
  output wire [5:0]    io_output_payload_fragment_length,
  output wire [3:0]    io_output_payload_fragment_context,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [1:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_maskProposal_1_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_1;
  wire                io_output_fire;
  wire                when_Stream_l683;
  wire                _zz_io_chosen;

  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz_maskProposal_1_2));
  assign _zz_maskProposal_1_2 = (_zz_maskProposal_1 - 2'b01);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_1 = {io_inputs_1_valid,io_inputs_0_valid};
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l683 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_output_payload_fragment_source = (maskRouted_0 ? io_inputs_0_payload_fragment_source : io_inputs_1_payload_fragment_source);
  assign io_output_payload_fragment_opcode = (maskRouted_0 ? io_inputs_0_payload_fragment_opcode : io_inputs_1_payload_fragment_opcode);
  assign io_output_payload_fragment_exclusive = (maskRouted_0 ? io_inputs_0_payload_fragment_exclusive : io_inputs_1_payload_fragment_exclusive);
  assign io_output_payload_fragment_address = (maskRouted_0 ? io_inputs_0_payload_fragment_address : io_inputs_1_payload_fragment_address);
  assign io_output_payload_fragment_length = (maskRouted_0 ? io_inputs_0_payload_fragment_length : io_inputs_1_payload_fragment_length);
  assign io_output_payload_fragment_context = (maskRouted_0 ? io_inputs_0_payload_fragment_context : io_inputs_1_payload_fragment_context);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l683) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
    end
  end


endmodule

module StreamArbiter_3 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire          io_inputs_0_payload_last,
  input  wire [0:0]    io_inputs_0_payload_fragment_source,
  input  wire [0:0]    io_inputs_0_payload_fragment_opcode,
  input  wire          io_inputs_0_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_0_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_payload_fragment_length,
  input  wire [3:0]    io_inputs_0_payload_fragment_context,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire          io_inputs_1_payload_last,
  input  wire [0:0]    io_inputs_1_payload_fragment_source,
  input  wire [0:0]    io_inputs_1_payload_fragment_opcode,
  input  wire          io_inputs_1_payload_fragment_exclusive,
  input  wire [31:0]   io_inputs_1_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_payload_fragment_length,
  input  wire [3:0]    io_inputs_1_payload_fragment_context,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [0:0]    io_output_payload_fragment_source,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire          io_output_payload_fragment_exclusive,
  output wire [31:0]   io_output_payload_fragment_address,
  output wire [5:0]    io_output_payload_fragment_length,
  output wire [3:0]    io_output_payload_fragment_context,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_output_payload_fragment_source = (maskRouted_0 ? io_inputs_0_payload_fragment_source : io_inputs_1_payload_fragment_source);
  assign io_output_payload_fragment_opcode = (maskRouted_0 ? io_inputs_0_payload_fragment_opcode : io_inputs_1_payload_fragment_opcode);
  assign io_output_payload_fragment_exclusive = (maskRouted_0 ? io_inputs_0_payload_fragment_exclusive : io_inputs_1_payload_fragment_exclusive);
  assign io_output_payload_fragment_address = (maskRouted_0 ? io_inputs_0_payload_fragment_address : io_inputs_1_payload_fragment_address);
  assign io_output_payload_fragment_length = (maskRouted_0 ? io_inputs_0_payload_fragment_length : io_inputs_1_payload_fragment_length);
  assign io_output_payload_fragment_context = (maskRouted_0 ? io_inputs_0_payload_fragment_context : io_inputs_1_payload_fragment_context);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [0:0]    io_push_payload,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [0:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [4:0]    io_occupancy,
  output wire [4:0]    io_availability,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg        [0:0]    logic_ram_spinal_port1;
  wire       [0:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [4:0]    logic_ptr_push;
  reg        [4:0]    logic_ptr_pop;
  wire       [4:0]    logic_ptr_occupancy;
  wire       [4:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [3:0]    logic_push_onRam_write_payload_address;
  wire       [0:0]    logic_push_onRam_write_payload_data;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [3:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [3:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [3:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [3:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [0:0]    logic_pop_sync_readPort_rsp;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [0:0]    logic_pop_sync_readArbitation_translated_payload;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [4:0]    logic_pop_sync_popReg;
  reg [0:0] logic_ram [0:15];

  assign _zz_logic_ram_port = logic_push_onRam_write_payload_data;
  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge io_systemClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 5'h10) == 5'h0);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[3:0];
  assign logic_push_onRam_write_payload_data = io_push_payload;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[3:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign logic_pop_sync_readPort_rsp = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload = logic_pop_sync_readPort_rsp;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload = logic_pop_sync_readArbitation_translated_payload;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (5'h10 - logic_ptr_occupancy);
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      logic_ptr_push <= 5'h0;
      logic_ptr_pop <= 5'h0;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 5'h0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 5'h01);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 5'h01);
      end
      if(io_flush) begin
        logic_ptr_push <= 5'h0;
        logic_ptr_pop <= 5'h0;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 5'h0;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module StreamArbiter_2 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire          io_inputs_0_payload_last,
  input  wire [0:0]    io_inputs_0_payload_fragment_source,
  input  wire [0:0]    io_inputs_0_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_0_payload_fragment_address,
  input  wire [5:0]    io_inputs_0_payload_fragment_length,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire          io_inputs_1_payload_last,
  input  wire [0:0]    io_inputs_1_payload_fragment_source,
  input  wire [0:0]    io_inputs_1_payload_fragment_opcode,
  input  wire [31:0]   io_inputs_1_payload_fragment_address,
  input  wire [5:0]    io_inputs_1_payload_fragment_length,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire          io_output_payload_last,
  output wire [0:0]    io_output_payload_fragment_source,
  output wire [0:0]    io_output_payload_fragment_opcode,
  output wire [31:0]   io_output_payload_fragment_address,
  output wire [5:0]    io_output_payload_fragment_length,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                when_Stream_l683;
  wire                _zz_io_chosen;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_Stream_l683 = (io_output_fire && io_output_payload_last);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_last = (maskRouted_0 ? io_inputs_0_payload_last : io_inputs_1_payload_last);
  assign io_output_payload_fragment_source = (maskRouted_0 ? io_inputs_0_payload_fragment_source : io_inputs_1_payload_fragment_source);
  assign io_output_payload_fragment_opcode = (maskRouted_0 ? io_inputs_0_payload_fragment_opcode : io_inputs_1_payload_fragment_opcode);
  assign io_output_payload_fragment_address = (maskRouted_0 ? io_inputs_0_payload_fragment_address : io_inputs_1_payload_fragment_address);
  assign io_output_payload_fragment_length = (maskRouted_0 ? io_inputs_0_payload_fragment_length : io_inputs_1_payload_fragment_length);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(when_Stream_l683) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

module FlowCCByToggle_1 (
  input  wire          io_input_valid,
  input  wire          io_input_payload_error,
  input  wire [31:0]   io_input_payload_data,
  output wire          io_output_valid,
  output wire          io_output_payload_error,
  output wire [31:0]   io_output_payload_data,
  input  wire          io_systemClk,
  input  wire          debugCd_logic_outputReset,
  input  wire          jtagCtrl_tck
);

  wire                system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  wire                inputArea_target_buffercc_io_dataOut;
  wire                system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_asyncAssertSyncDeassert;
  wire                system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_synchronized;
  reg                 inputArea_target;
  reg                 inputArea_data_error;
  reg        [31:0]   inputArea_data_data;
  wire                outputArea_target;
  reg                 outputArea_hit;
  wire                outputArea_flow_valid;
  wire                outputArea_flow_payload_error;
  wire       [31:0]   outputArea_flow_payload_data;
  reg                 outputArea_flow_m2sPipe_valid;
  (* async_reg = "true" *) reg                 outputArea_flow_m2sPipe_payload_error;
  (* async_reg = "true" *) reg        [31:0]   outputArea_flow_m2sPipe_payload_data;

  (* keep_hierarchy = "TRUE" *) BufferCC_3 system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc (
    .io_dataIn                 (system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_asyncAssertSyncDeassert                    ), //i
    .io_dataOut                (system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut), //o
    .jtagCtrl_tck              (jtagCtrl_tck                                                                                                     ), //i
    .debugCd_logic_outputReset (debugCd_logic_outputReset                                                                                        )  //i
  );
  (* keep_hierarchy = "TRUE" *) BufferCC_4 inputArea_target_buffercc (
    .io_dataIn                                                                          (inputArea_target                                                                  ), //i
    .io_dataOut                                                                         (inputArea_target_buffercc_io_dataOut                                              ), //o
    .jtagCtrl_tck                                                                       (jtagCtrl_tck                                                                      ), //i
    .system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_synchronized (system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_synchronized)  //i
  );
  assign system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_asyncAssertSyncDeassert = (1'b0 ^ 1'b0);
  assign system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_synchronized = system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_asyncAssertSyncDeassert_buffercc_io_dataOut;
  assign outputArea_target = inputArea_target_buffercc_io_dataOut;
  assign outputArea_flow_valid = (outputArea_target != outputArea_hit);
  assign outputArea_flow_payload_error = inputArea_data_error;
  assign outputArea_flow_payload_data = inputArea_data_data;
  assign io_output_valid = outputArea_flow_m2sPipe_valid;
  assign io_output_payload_error = outputArea_flow_m2sPipe_payload_error;
  assign io_output_payload_data = outputArea_flow_m2sPipe_payload_data;
  always @(posedge io_systemClk) begin
    if(debugCd_logic_outputReset) begin
      inputArea_target <= 1'b0;
    end else begin
      if(io_input_valid) begin
        inputArea_target <= (! inputArea_target);
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_input_valid) begin
      inputArea_data_error <= io_input_payload_error;
      inputArea_data_data <= io_input_payload_data;
    end
  end

  always @(posedge jtagCtrl_tck) begin
    if(system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_synchronized) begin
      outputArea_flow_m2sPipe_valid <= 1'b0;
      outputArea_hit <= 1'b0;
    end else begin
      outputArea_hit <= outputArea_target;
      outputArea_flow_m2sPipe_valid <= outputArea_flow_valid;
    end
  end

  always @(posedge jtagCtrl_tck) begin
    if(outputArea_flow_valid) begin
      outputArea_flow_m2sPipe_payload_error <= outputArea_flow_payload_error;
      outputArea_flow_m2sPipe_payload_data <= outputArea_flow_payload_data;
    end
  end


endmodule

module FlowCCByToggle (
  input  wire          io_input_valid,
  input  wire          io_input_payload_write,
  input  wire [31:0]   io_input_payload_data,
  input  wire [6:0]    io_input_payload_address,
  output wire          io_output_valid,
  output wire          io_output_payload_write,
  output wire [31:0]   io_output_payload_data,
  output wire [6:0]    io_output_payload_address,
  input  wire          jtagCtrl_tck,
  input  wire          io_systemClk,
  input  wire          debugCd_logic_outputReset
);

  wire                inputArea_target_buffercc_io_dataOut;
  reg                 inputArea_target;
  reg                 inputArea_data_write;
  reg        [31:0]   inputArea_data_data;
  reg        [6:0]    inputArea_data_address;
  wire                outputArea_target;
  reg                 outputArea_hit;
  wire                outputArea_flow_valid;
  wire                outputArea_flow_payload_write;
  wire       [31:0]   outputArea_flow_payload_data;
  wire       [6:0]    outputArea_flow_payload_address;

  (* keep_hierarchy = "TRUE" *) BufferCC_2 inputArea_target_buffercc (
    .io_dataIn                 (inputArea_target                    ), //i
    .io_dataOut                (inputArea_target_buffercc_io_dataOut), //o
    .io_systemClk              (io_systemClk                        ), //i
    .debugCd_logic_outputReset (debugCd_logic_outputReset           )  //i
  );
  initial begin
  `ifndef SYNTHESIS
    inputArea_target = $urandom;
    outputArea_hit = $urandom;
  `endif
  end

  assign outputArea_target = inputArea_target_buffercc_io_dataOut;
  assign outputArea_flow_valid = (outputArea_target != outputArea_hit);
  assign outputArea_flow_payload_write = inputArea_data_write;
  assign outputArea_flow_payload_data = inputArea_data_data;
  assign outputArea_flow_payload_address = inputArea_data_address;
  assign io_output_valid = outputArea_flow_valid;
  assign io_output_payload_write = outputArea_flow_payload_write;
  assign io_output_payload_data = outputArea_flow_payload_data;
  assign io_output_payload_address = outputArea_flow_payload_address;
  always @(posedge jtagCtrl_tck) begin
    if(io_input_valid) begin
      inputArea_target <= (! inputArea_target);
      inputArea_data_write <= io_input_payload_write;
      inputArea_data_data <= io_input_payload_data;
      inputArea_data_address <= io_input_payload_address;
    end
  end

  always @(posedge io_systemClk) begin
    outputArea_hit <= outputArea_target;
  end


endmodule

module StreamArbiter_1 (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [0:0]    io_inputs_0_payload_source,
  input  wire [4:0]    io_inputs_0_payload_rd,
  input  wire [52:0]   io_inputs_0_payload_value_mantissa,
  input  wire [11:0]   io_inputs_0_payload_value_exponent,
  input  wire          io_inputs_0_payload_value_sign,
  input  wire          io_inputs_0_payload_value_special,
  input  wire          io_inputs_0_payload_scrap,
  input  wire [2:0]    io_inputs_0_payload_roundMode,
  input  wire [0:0]    io_inputs_0_payload_format,
  input  wire          io_inputs_0_payload_NV,
  input  wire          io_inputs_0_payload_DZ,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [0:0]    io_inputs_1_payload_source,
  input  wire [4:0]    io_inputs_1_payload_rd,
  input  wire [52:0]   io_inputs_1_payload_value_mantissa,
  input  wire [11:0]   io_inputs_1_payload_value_exponent,
  input  wire          io_inputs_1_payload_value_sign,
  input  wire          io_inputs_1_payload_value_special,
  input  wire          io_inputs_1_payload_scrap,
  input  wire [2:0]    io_inputs_1_payload_roundMode,
  input  wire [0:0]    io_inputs_1_payload_format,
  input  wire          io_inputs_1_payload_NV,
  input  wire          io_inputs_1_payload_DZ,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [0:0]    io_inputs_2_payload_source,
  input  wire [4:0]    io_inputs_2_payload_rd,
  input  wire [52:0]   io_inputs_2_payload_value_mantissa,
  input  wire [11:0]   io_inputs_2_payload_value_exponent,
  input  wire          io_inputs_2_payload_value_sign,
  input  wire          io_inputs_2_payload_value_special,
  input  wire          io_inputs_2_payload_scrap,
  input  wire [2:0]    io_inputs_2_payload_roundMode,
  input  wire [0:0]    io_inputs_2_payload_format,
  input  wire          io_inputs_2_payload_NV,
  input  wire          io_inputs_2_payload_DZ,
  input  wire          io_inputs_3_valid,
  output wire          io_inputs_3_ready,
  input  wire [0:0]    io_inputs_3_payload_source,
  input  wire [4:0]    io_inputs_3_payload_rd,
  input  wire [52:0]   io_inputs_3_payload_value_mantissa,
  input  wire [11:0]   io_inputs_3_payload_value_exponent,
  input  wire          io_inputs_3_payload_value_sign,
  input  wire          io_inputs_3_payload_value_special,
  input  wire          io_inputs_3_payload_scrap,
  input  wire [2:0]    io_inputs_3_payload_roundMode,
  input  wire [0:0]    io_inputs_3_payload_format,
  input  wire          io_inputs_3_payload_NV,
  input  wire          io_inputs_3_payload_DZ,
  input  wire          io_inputs_4_valid,
  output wire          io_inputs_4_ready,
  input  wire [0:0]    io_inputs_4_payload_source,
  input  wire [4:0]    io_inputs_4_payload_rd,
  input  wire [52:0]   io_inputs_4_payload_value_mantissa,
  input  wire [11:0]   io_inputs_4_payload_value_exponent,
  input  wire          io_inputs_4_payload_value_sign,
  input  wire          io_inputs_4_payload_value_special,
  input  wire          io_inputs_4_payload_scrap,
  input  wire [2:0]    io_inputs_4_payload_roundMode,
  input  wire [0:0]    io_inputs_4_payload_format,
  input  wire          io_inputs_4_payload_NV,
  input  wire          io_inputs_4_payload_DZ,
  input  wire          io_inputs_5_valid,
  output wire          io_inputs_5_ready,
  input  wire [0:0]    io_inputs_5_payload_source,
  input  wire [4:0]    io_inputs_5_payload_rd,
  input  wire [52:0]   io_inputs_5_payload_value_mantissa,
  input  wire [11:0]   io_inputs_5_payload_value_exponent,
  input  wire          io_inputs_5_payload_value_sign,
  input  wire          io_inputs_5_payload_value_special,
  input  wire          io_inputs_5_payload_scrap,
  input  wire [2:0]    io_inputs_5_payload_roundMode,
  input  wire [0:0]    io_inputs_5_payload_format,
  input  wire          io_inputs_5_payload_NV,
  input  wire          io_inputs_5_payload_DZ,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [0:0]    io_output_payload_source,
  output wire [4:0]    io_output_payload_rd,
  output wire [52:0]   io_output_payload_value_mantissa,
  output wire [11:0]   io_output_payload_value_exponent,
  output wire          io_output_payload_value_sign,
  output wire          io_output_payload_value_special,
  output wire          io_output_payload_scrap,
  output wire [2:0]    io_output_payload_roundMode,
  output wire [0:0]    io_output_payload_format,
  output wire          io_output_payload_NV,
  output wire          io_output_payload_DZ,
  output wire [2:0]    io_chosen,
  output wire [5:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);
  localparam FpuRoundMode_RNE = 3'd0;
  localparam FpuRoundMode_RTZ = 3'd1;
  localparam FpuRoundMode_RDN = 3'd2;
  localparam FpuRoundMode_RUP = 3'd3;
  localparam FpuRoundMode_RMM = 3'd4;
  localparam FpuFormat_FLOAT = 1'd0;
  localparam FpuFormat_DOUBLE = 1'd1;

  wire       [5:0]    _zz__zz_maskProposal_1_1;
  reg        [2:0]    _zz__zz_io_output_payload_roundMode;
  reg        [0:0]    _zz__zz_io_output_payload_format;
  reg        [0:0]    _zz_io_output_payload_source_4;
  reg        [4:0]    _zz_io_output_payload_rd;
  reg        [52:0]   _zz_io_output_payload_value_mantissa;
  reg        [11:0]   _zz_io_output_payload_value_exponent;
  reg                 _zz_io_output_payload_value_sign;
  reg                 _zz_io_output_payload_value_special;
  reg                 _zz_io_output_payload_scrap;
  reg                 _zz_io_output_payload_NV;
  reg                 _zz_io_output_payload_DZ;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  wire                maskProposal_3;
  wire                maskProposal_4;
  wire                maskProposal_5;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  reg                 maskLocked_3;
  reg                 maskLocked_4;
  reg                 maskLocked_5;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire                maskRouted_3;
  wire                maskRouted_4;
  wire                maskRouted_5;
  wire       [5:0]    _zz_maskProposal_1;
  wire       [5:0]    _zz_maskProposal_1_1;
  wire                _zz_io_output_payload_source;
  wire                _zz_io_output_payload_source_1;
  wire                _zz_io_output_payload_source_2;
  wire       [2:0]    _zz_io_output_payload_source_3;
  wire       [2:0]    _zz_io_output_payload_roundMode;
  wire       [0:0]    _zz_io_output_payload_format;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  wire                _zz_io_chosen_2;
  wire                _zz_io_chosen_3;
  wire                _zz_io_chosen_4;
  `ifndef SYNTHESIS
  reg [23:0] io_inputs_0_payload_roundMode_string;
  reg [47:0] io_inputs_0_payload_format_string;
  reg [23:0] io_inputs_1_payload_roundMode_string;
  reg [47:0] io_inputs_1_payload_format_string;
  reg [23:0] io_inputs_2_payload_roundMode_string;
  reg [47:0] io_inputs_2_payload_format_string;
  reg [23:0] io_inputs_3_payload_roundMode_string;
  reg [47:0] io_inputs_3_payload_format_string;
  reg [23:0] io_inputs_4_payload_roundMode_string;
  reg [47:0] io_inputs_4_payload_format_string;
  reg [23:0] io_inputs_5_payload_roundMode_string;
  reg [47:0] io_inputs_5_payload_format_string;
  reg [23:0] io_output_payload_roundMode_string;
  reg [47:0] io_output_payload_format_string;
  reg [23:0] _zz_io_output_payload_roundMode_string;
  reg [47:0] _zz_io_output_payload_format_string;
  `endif


  assign _zz__zz_maskProposal_1_1 = (_zz_maskProposal_1 - 6'h01);
  always @(*) begin
    case(_zz_io_output_payload_source_3)
      3'b000 : begin
        _zz__zz_io_output_payload_roundMode = io_inputs_0_payload_roundMode;
        _zz__zz_io_output_payload_format = io_inputs_0_payload_format;
        _zz_io_output_payload_source_4 = io_inputs_0_payload_source;
        _zz_io_output_payload_rd = io_inputs_0_payload_rd;
        _zz_io_output_payload_value_mantissa = io_inputs_0_payload_value_mantissa;
        _zz_io_output_payload_value_exponent = io_inputs_0_payload_value_exponent;
        _zz_io_output_payload_value_sign = io_inputs_0_payload_value_sign;
        _zz_io_output_payload_value_special = io_inputs_0_payload_value_special;
        _zz_io_output_payload_scrap = io_inputs_0_payload_scrap;
        _zz_io_output_payload_NV = io_inputs_0_payload_NV;
        _zz_io_output_payload_DZ = io_inputs_0_payload_DZ;
      end
      3'b001 : begin
        _zz__zz_io_output_payload_roundMode = io_inputs_1_payload_roundMode;
        _zz__zz_io_output_payload_format = io_inputs_1_payload_format;
        _zz_io_output_payload_source_4 = io_inputs_1_payload_source;
        _zz_io_output_payload_rd = io_inputs_1_payload_rd;
        _zz_io_output_payload_value_mantissa = io_inputs_1_payload_value_mantissa;
        _zz_io_output_payload_value_exponent = io_inputs_1_payload_value_exponent;
        _zz_io_output_payload_value_sign = io_inputs_1_payload_value_sign;
        _zz_io_output_payload_value_special = io_inputs_1_payload_value_special;
        _zz_io_output_payload_scrap = io_inputs_1_payload_scrap;
        _zz_io_output_payload_NV = io_inputs_1_payload_NV;
        _zz_io_output_payload_DZ = io_inputs_1_payload_DZ;
      end
      3'b010 : begin
        _zz__zz_io_output_payload_roundMode = io_inputs_2_payload_roundMode;
        _zz__zz_io_output_payload_format = io_inputs_2_payload_format;
        _zz_io_output_payload_source_4 = io_inputs_2_payload_source;
        _zz_io_output_payload_rd = io_inputs_2_payload_rd;
        _zz_io_output_payload_value_mantissa = io_inputs_2_payload_value_mantissa;
        _zz_io_output_payload_value_exponent = io_inputs_2_payload_value_exponent;
        _zz_io_output_payload_value_sign = io_inputs_2_payload_value_sign;
        _zz_io_output_payload_value_special = io_inputs_2_payload_value_special;
        _zz_io_output_payload_scrap = io_inputs_2_payload_scrap;
        _zz_io_output_payload_NV = io_inputs_2_payload_NV;
        _zz_io_output_payload_DZ = io_inputs_2_payload_DZ;
      end
      3'b011 : begin
        _zz__zz_io_output_payload_roundMode = io_inputs_3_payload_roundMode;
        _zz__zz_io_output_payload_format = io_inputs_3_payload_format;
        _zz_io_output_payload_source_4 = io_inputs_3_payload_source;
        _zz_io_output_payload_rd = io_inputs_3_payload_rd;
        _zz_io_output_payload_value_mantissa = io_inputs_3_payload_value_mantissa;
        _zz_io_output_payload_value_exponent = io_inputs_3_payload_value_exponent;
        _zz_io_output_payload_value_sign = io_inputs_3_payload_value_sign;
        _zz_io_output_payload_value_special = io_inputs_3_payload_value_special;
        _zz_io_output_payload_scrap = io_inputs_3_payload_scrap;
        _zz_io_output_payload_NV = io_inputs_3_payload_NV;
        _zz_io_output_payload_DZ = io_inputs_3_payload_DZ;
      end
      3'b100 : begin
        _zz__zz_io_output_payload_roundMode = io_inputs_4_payload_roundMode;
        _zz__zz_io_output_payload_format = io_inputs_4_payload_format;
        _zz_io_output_payload_source_4 = io_inputs_4_payload_source;
        _zz_io_output_payload_rd = io_inputs_4_payload_rd;
        _zz_io_output_payload_value_mantissa = io_inputs_4_payload_value_mantissa;
        _zz_io_output_payload_value_exponent = io_inputs_4_payload_value_exponent;
        _zz_io_output_payload_value_sign = io_inputs_4_payload_value_sign;
        _zz_io_output_payload_value_special = io_inputs_4_payload_value_special;
        _zz_io_output_payload_scrap = io_inputs_4_payload_scrap;
        _zz_io_output_payload_NV = io_inputs_4_payload_NV;
        _zz_io_output_payload_DZ = io_inputs_4_payload_DZ;
      end
      default : begin
        _zz__zz_io_output_payload_roundMode = io_inputs_5_payload_roundMode;
        _zz__zz_io_output_payload_format = io_inputs_5_payload_format;
        _zz_io_output_payload_source_4 = io_inputs_5_payload_source;
        _zz_io_output_payload_rd = io_inputs_5_payload_rd;
        _zz_io_output_payload_value_mantissa = io_inputs_5_payload_value_mantissa;
        _zz_io_output_payload_value_exponent = io_inputs_5_payload_value_exponent;
        _zz_io_output_payload_value_sign = io_inputs_5_payload_value_sign;
        _zz_io_output_payload_value_special = io_inputs_5_payload_value_special;
        _zz_io_output_payload_scrap = io_inputs_5_payload_scrap;
        _zz_io_output_payload_NV = io_inputs_5_payload_NV;
        _zz_io_output_payload_DZ = io_inputs_5_payload_DZ;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_0_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_0_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_0_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_0_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_0_payload_roundMode_string = "RMM";
      default : io_inputs_0_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_inputs_0_payload_format)
      FpuFormat_FLOAT : io_inputs_0_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_0_payload_format_string = "DOUBLE";
      default : io_inputs_0_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_1_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_1_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_1_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_1_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_1_payload_roundMode_string = "RMM";
      default : io_inputs_1_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_format)
      FpuFormat_FLOAT : io_inputs_1_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_1_payload_format_string = "DOUBLE";
      default : io_inputs_1_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_2_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_2_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_2_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_2_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_2_payload_roundMode_string = "RMM";
      default : io_inputs_2_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_inputs_2_payload_format)
      FpuFormat_FLOAT : io_inputs_2_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_2_payload_format_string = "DOUBLE";
      default : io_inputs_2_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_3_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_3_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_3_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_3_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_3_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_3_payload_roundMode_string = "RMM";
      default : io_inputs_3_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_inputs_3_payload_format)
      FpuFormat_FLOAT : io_inputs_3_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_3_payload_format_string = "DOUBLE";
      default : io_inputs_3_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_4_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_4_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_4_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_4_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_4_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_4_payload_roundMode_string = "RMM";
      default : io_inputs_4_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_inputs_4_payload_format)
      FpuFormat_FLOAT : io_inputs_4_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_4_payload_format_string = "DOUBLE";
      default : io_inputs_4_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_5_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_5_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_5_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_5_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_5_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_5_payload_roundMode_string = "RMM";
      default : io_inputs_5_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_inputs_5_payload_format)
      FpuFormat_FLOAT : io_inputs_5_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_5_payload_format_string = "DOUBLE";
      default : io_inputs_5_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_roundMode)
      FpuRoundMode_RNE : io_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_output_payload_roundMode_string = "RMM";
      default : io_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_output_payload_format)
      FpuFormat_FLOAT : io_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_output_payload_format_string = "DOUBLE";
      default : io_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_roundMode)
      FpuRoundMode_RNE : _zz_io_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : _zz_io_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : _zz_io_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : _zz_io_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : _zz_io_output_payload_roundMode_string = "RMM";
      default : _zz_io_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_format)
      FpuFormat_FLOAT : _zz_io_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_io_output_payload_format_string = "DOUBLE";
      default : _zz_io_output_payload_format_string = "??????";
    endcase
  end
  `endif

  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign maskRouted_3 = (locked ? maskLocked_3 : maskProposal_3);
  assign maskRouted_4 = (locked ? maskLocked_4 : maskProposal_4);
  assign maskRouted_5 = (locked ? maskLocked_5 : maskProposal_5);
  assign _zz_maskProposal_1 = {io_inputs_5_valid,{io_inputs_4_valid,{io_inputs_3_valid,{io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}}}}};
  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz__zz_maskProposal_1_1));
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign maskProposal_2 = _zz_maskProposal_1_1[2];
  assign maskProposal_3 = _zz_maskProposal_1_1[3];
  assign maskProposal_4 = _zz_maskProposal_1_1[4];
  assign maskProposal_5 = _zz_maskProposal_1_1[5];
  assign io_output_valid = ((((((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2)) || (io_inputs_3_valid && maskRouted_3)) || (io_inputs_4_valid && maskRouted_4)) || (io_inputs_5_valid && maskRouted_5));
  assign _zz_io_output_payload_source = ((maskRouted_1 || maskRouted_3) || maskRouted_5);
  assign _zz_io_output_payload_source_1 = (maskRouted_2 || maskRouted_3);
  assign _zz_io_output_payload_source_2 = (maskRouted_4 || maskRouted_5);
  assign _zz_io_output_payload_source_3 = {_zz_io_output_payload_source_2,{_zz_io_output_payload_source_1,_zz_io_output_payload_source}};
  assign _zz_io_output_payload_roundMode = _zz__zz_io_output_payload_roundMode;
  assign _zz_io_output_payload_format = _zz__zz_io_output_payload_format;
  assign io_output_payload_source = _zz_io_output_payload_source_4;
  assign io_output_payload_rd = _zz_io_output_payload_rd;
  assign io_output_payload_value_mantissa = _zz_io_output_payload_value_mantissa;
  assign io_output_payload_value_exponent = _zz_io_output_payload_value_exponent;
  assign io_output_payload_value_sign = _zz_io_output_payload_value_sign;
  assign io_output_payload_value_special = _zz_io_output_payload_value_special;
  assign io_output_payload_scrap = _zz_io_output_payload_scrap;
  assign io_output_payload_roundMode = _zz_io_output_payload_roundMode;
  assign io_output_payload_format = _zz_io_output_payload_format;
  assign io_output_payload_NV = _zz_io_output_payload_NV;
  assign io_output_payload_DZ = _zz_io_output_payload_DZ;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_inputs_3_ready = (maskRouted_3 && io_output_ready);
  assign io_inputs_4_ready = (maskRouted_4 && io_output_ready);
  assign io_inputs_5_ready = (maskRouted_5 && io_output_ready);
  assign io_chosenOH = {maskRouted_5,{maskRouted_4,{maskRouted_3,{maskRouted_2,{maskRouted_1,maskRouted_0}}}}};
  assign _zz_io_chosen = io_chosenOH[3];
  assign _zz_io_chosen_1 = io_chosenOH[5];
  assign _zz_io_chosen_2 = ((io_chosenOH[1] || _zz_io_chosen) || _zz_io_chosen_1);
  assign _zz_io_chosen_3 = (io_chosenOH[2] || _zz_io_chosen);
  assign _zz_io_chosen_4 = (io_chosenOH[4] || _zz_io_chosen_1);
  assign io_chosen = {_zz_io_chosen_4,{_zz_io_chosen_3,_zz_io_chosen_2}};
  always @(posedge io_systemClk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
      maskLocked_2 <= maskRouted_2;
      maskLocked_3 <= maskRouted_3;
      maskLocked_4 <= maskRouted_4;
      maskLocked_5 <= maskRouted_5;
    end
  end


endmodule

module FpuSqrt (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [53:0]   io_input_payload_a,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [52:0]   io_output_payload_result,
  output wire [56:0]   io_output_payload_remain,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [56:0]   _zz_t;
  wire       [54:0]   _zz_t_1;
  wire       [53:0]   _zz_q;
  wire       [58:0]   _zz_a_1;
  wire       [1:0]    _zz_a_2;
  reg        [5:0]    counter;
  reg                 busy;
  wire                io_output_fire;
  reg                 done;
  wire                when_FpuSqrt_l28;
  reg        [56:0]   a;
  reg        [51:0]   x;
  reg        [52:0]   q;
  wire       [56:0]   t;
  wire                when_FpuSqrt_l41;
  reg        [56:0]   _zz_a;
  wire                when_FpuSqrt_l44;
  wire                when_FpuSqrt_l52;

  assign _zz_t_1 = {q,2'b01};
  assign _zz_t = {2'd0, _zz_t_1};
  assign _zz_q = {q,(! t[56])};
  assign _zz_a_1 = {_zz_a,x[51 : 50]};
  assign _zz_a_2 = io_input_payload_a[53 : 52];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_FpuSqrt_l28 = (busy && (counter == 6'h35));
  assign t = (a - _zz_t);
  assign io_output_valid = done;
  assign io_output_payload_result = q;
  assign io_output_payload_remain = a;
  assign io_input_ready = (! busy);
  assign when_FpuSqrt_l41 = (! done);
  always @(*) begin
    _zz_a = a;
    if(when_FpuSqrt_l44) begin
      _zz_a = t;
    end
  end

  assign when_FpuSqrt_l44 = (! t[56]);
  assign when_FpuSqrt_l52 = (! busy);
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      busy <= 1'b0;
      done <= 1'b0;
    end else begin
      if(io_output_fire) begin
        busy <= 1'b0;
      end
      if(when_FpuSqrt_l28) begin
        done <= 1'b1;
      end
      if(io_output_fire) begin
        done <= 1'b0;
      end
      if(when_FpuSqrt_l52) begin
        if(io_input_valid) begin
          busy <= 1'b1;
        end
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(when_FpuSqrt_l41) begin
      counter <= (counter + 6'h01);
      q <= _zz_q[52:0];
      a <= _zz_a_1[56:0];
      x <= (x <<< 2);
    end
    if(when_FpuSqrt_l52) begin
      q <= 53'h0;
      a <= {55'd0, _zz_a_2};
      x <= io_input_payload_a[51:0];
      counter <= 6'h0;
    end
  end


endmodule

module FpuDiv (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [51:0]   io_input_payload_a,
  input  wire [51:0]   io_input_payload_b,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [54:0]   io_output_payload_result,
  output wire [52:0]   io_output_payload_remain,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  wire       [52:0]   _zz_shifter_1;
  wire       [52:0]   _zz_div1;
  wire       [54:0]   _zz_div3;
  wire       [53:0]   _zz_div3_1;
  wire       [53:0]   _zz_div3_2;
  reg        [4:0]    counter;
  reg                 busy;
  wire                io_output_fire;
  reg                 done;
  wire                when_FpuDiv_l31;
  reg        [54:0]   shifter;
  reg        [54:0]   result;
  reg        [54:0]   div1;
  reg        [54:0]   div3;
  wire       [54:0]   div2;
  wire       [55:0]   sub1;
  wire       [55:0]   sub2;
  wire       [55:0]   sub3;
  wire                when_FpuDiv_l48;
  reg        [54:0]   _zz_shifter;
  wire                when_FpuDiv_l52;
  wire                when_FpuDiv_l56;
  wire                when_FpuDiv_l60;
  wire                when_FpuDiv_l67;

  assign _zz_shifter_1 = {1'b1,io_input_payload_a};
  assign _zz_div1 = {1'b1,io_input_payload_b};
  assign _zz_div3_1 = {1'b0,{1'b1,io_input_payload_b}};
  assign _zz_div3 = {1'd0, _zz_div3_1};
  assign _zz_div3_2 = ({1'd0,{1'b1,io_input_payload_b}} <<< 1'd1);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_FpuDiv_l31 = (busy && (counter == 5'h1b));
  assign div2 = (div1 <<< 1);
  assign sub1 = ({1'b0,shifter} - {1'b0,div1});
  assign sub2 = ({1'b0,shifter} - {1'b0,div2});
  assign sub3 = ({1'b0,shifter} - {1'b0,div3});
  assign io_output_valid = done;
  assign io_output_payload_result = result;
  assign io_output_payload_remain = (shifter >>> 2'd2);
  assign io_input_ready = (! busy);
  assign when_FpuDiv_l48 = (! done);
  always @(*) begin
    _zz_shifter = shifter;
    if(when_FpuDiv_l52) begin
      _zz_shifter = sub1[54:0];
    end
    if(when_FpuDiv_l56) begin
      _zz_shifter = sub2[54:0];
    end
    if(when_FpuDiv_l60) begin
      _zz_shifter = sub3[54:0];
    end
  end

  assign when_FpuDiv_l52 = (! sub1[55]);
  assign when_FpuDiv_l56 = (! sub2[55]);
  assign when_FpuDiv_l60 = (! sub3[55]);
  assign when_FpuDiv_l67 = (! busy);
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      busy <= 1'b0;
      done <= 1'b0;
    end else begin
      if(io_output_fire) begin
        busy <= 1'b0;
      end
      if(when_FpuDiv_l31) begin
        done <= 1'b1;
      end
      if(io_output_fire) begin
        done <= 1'b0;
      end
      if(when_FpuDiv_l67) begin
        busy <= io_input_valid;
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(when_FpuDiv_l48) begin
      counter <= (counter + 5'h01);
      result <= (result <<< 2);
      if(when_FpuDiv_l52) begin
        result[1 : 0] <= 2'b01;
      end
      if(when_FpuDiv_l56) begin
        result[1 : 0] <= 2'b10;
      end
      if(when_FpuDiv_l60) begin
        result[1 : 0] <= 2'b11;
      end
      shifter <= (_zz_shifter <<< 2);
    end
    if(when_FpuDiv_l67) begin
      counter <= 5'h0;
      shifter <= {2'd0, _zz_shifter_1};
      div1 <= {2'd0, _zz_div1};
      div3 <= (_zz_div3 + {1'b0,_zz_div3_2});
    end
  end


endmodule

module StreamArbiter (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [3:0]    io_inputs_0_payload_opcode,
  input  wire [1:0]    io_inputs_0_payload_arg,
  input  wire [4:0]    io_inputs_0_payload_rs1,
  input  wire [4:0]    io_inputs_0_payload_rs2,
  input  wire [4:0]    io_inputs_0_payload_rs3,
  input  wire [4:0]    io_inputs_0_payload_rd,
  input  wire [0:0]    io_inputs_0_payload_format,
  input  wire [2:0]    io_inputs_0_payload_roundMode,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [3:0]    io_inputs_1_payload_opcode,
  input  wire [1:0]    io_inputs_1_payload_arg,
  input  wire [4:0]    io_inputs_1_payload_rs1,
  input  wire [4:0]    io_inputs_1_payload_rs2,
  input  wire [4:0]    io_inputs_1_payload_rs3,
  input  wire [4:0]    io_inputs_1_payload_rd,
  input  wire [0:0]    io_inputs_1_payload_format,
  input  wire [2:0]    io_inputs_1_payload_roundMode,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [3:0]    io_output_payload_opcode,
  output wire [1:0]    io_output_payload_arg,
  output wire [4:0]    io_output_payload_rs1,
  output wire [4:0]    io_output_payload_rs2,
  output wire [4:0]    io_output_payload_rs3,
  output wire [4:0]    io_output_payload_rd,
  output wire [0:0]    io_output_payload_format,
  output wire [2:0]    io_output_payload_roundMode,
  output wire [0:0]    io_chosen,
  output wire [1:0]    io_chosenOH,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);
  localparam FpuOpcode_LOAD = 4'd0;
  localparam FpuOpcode_STORE = 4'd1;
  localparam FpuOpcode_MUL = 4'd2;
  localparam FpuOpcode_ADD = 4'd3;
  localparam FpuOpcode_FMA = 4'd4;
  localparam FpuOpcode_I2F = 4'd5;
  localparam FpuOpcode_F2I = 4'd6;
  localparam FpuOpcode_CMP = 4'd7;
  localparam FpuOpcode_DIV = 4'd8;
  localparam FpuOpcode_SQRT = 4'd9;
  localparam FpuOpcode_MIN_MAX = 4'd10;
  localparam FpuOpcode_SGNJ = 4'd11;
  localparam FpuOpcode_FMV_X_W = 4'd12;
  localparam FpuOpcode_FMV_W_X = 4'd13;
  localparam FpuOpcode_FCLASS = 4'd14;
  localparam FpuOpcode_FCVT_X_X = 4'd15;
  localparam FpuFormat_FLOAT = 1'd0;
  localparam FpuFormat_DOUBLE = 1'd1;
  localparam FpuRoundMode_RNE = 3'd0;
  localparam FpuRoundMode_RTZ = 3'd1;
  localparam FpuRoundMode_RDN = 3'd2;
  localparam FpuRoundMode_RUP = 3'd3;
  localparam FpuRoundMode_RMM = 3'd4;

  wire       [3:0]    _zz__zz_maskProposal_0_2;
  wire       [3:0]    _zz__zz_maskProposal_0_2_1;
  wire       [1:0]    _zz__zz_maskProposal_0_2_2;
  wire                locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_0;
  wire       [3:0]    _zz_maskProposal_0_1;
  wire       [3:0]    _zz_maskProposal_0_2;
  wire       [1:0]    _zz_maskProposal_0_3;
  wire       [3:0]    _zz_io_output_payload_opcode;
  wire       [0:0]    _zz_io_output_payload_format;
  wire       [2:0]    _zz_io_output_payload_roundMode;
  wire                _zz_io_chosen;
  `ifndef SYNTHESIS
  reg [63:0] io_inputs_0_payload_opcode_string;
  reg [47:0] io_inputs_0_payload_format_string;
  reg [23:0] io_inputs_0_payload_roundMode_string;
  reg [63:0] io_inputs_1_payload_opcode_string;
  reg [47:0] io_inputs_1_payload_format_string;
  reg [23:0] io_inputs_1_payload_roundMode_string;
  reg [63:0] io_output_payload_opcode_string;
  reg [47:0] io_output_payload_format_string;
  reg [23:0] io_output_payload_roundMode_string;
  reg [63:0] _zz_io_output_payload_opcode_string;
  reg [47:0] _zz_io_output_payload_format_string;
  reg [23:0] _zz_io_output_payload_roundMode_string;
  `endif


  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_0,maskLocked_1};
  assign _zz__zz_maskProposal_0_2_1 = {2'd0, _zz__zz_maskProposal_0_2_2};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_inputs_0_payload_opcode)
      FpuOpcode_LOAD : io_inputs_0_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_inputs_0_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_inputs_0_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_inputs_0_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_inputs_0_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_inputs_0_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_inputs_0_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_inputs_0_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_inputs_0_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_inputs_0_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_inputs_0_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_inputs_0_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_inputs_0_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_inputs_0_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_inputs_0_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_inputs_0_payload_opcode_string = "FCVT_X_X";
      default : io_inputs_0_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_0_payload_format)
      FpuFormat_FLOAT : io_inputs_0_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_0_payload_format_string = "DOUBLE";
      default : io_inputs_0_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_0_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_0_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_0_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_0_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_0_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_0_payload_roundMode_string = "RMM";
      default : io_inputs_0_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_opcode)
      FpuOpcode_LOAD : io_inputs_1_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_inputs_1_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_inputs_1_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_inputs_1_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_inputs_1_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_inputs_1_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_inputs_1_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_inputs_1_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_inputs_1_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_inputs_1_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_inputs_1_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_inputs_1_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_inputs_1_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_inputs_1_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_inputs_1_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_inputs_1_payload_opcode_string = "FCVT_X_X";
      default : io_inputs_1_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_format)
      FpuFormat_FLOAT : io_inputs_1_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_inputs_1_payload_format_string = "DOUBLE";
      default : io_inputs_1_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_inputs_1_payload_roundMode)
      FpuRoundMode_RNE : io_inputs_1_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_inputs_1_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_inputs_1_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_inputs_1_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_inputs_1_payload_roundMode_string = "RMM";
      default : io_inputs_1_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(io_output_payload_opcode)
      FpuOpcode_LOAD : io_output_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_output_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_output_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_output_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_output_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_output_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_output_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_output_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_output_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_output_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_output_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_output_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_output_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_output_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_output_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_output_payload_opcode_string = "FCVT_X_X";
      default : io_output_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_format)
      FpuFormat_FLOAT : io_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : io_output_payload_format_string = "DOUBLE";
      default : io_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(io_output_payload_roundMode)
      FpuRoundMode_RNE : io_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : io_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : io_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : io_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : io_output_payload_roundMode_string = "RMM";
      default : io_output_payload_roundMode_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_opcode)
      FpuOpcode_LOAD : _zz_io_output_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : _zz_io_output_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : _zz_io_output_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : _zz_io_output_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : _zz_io_output_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : _zz_io_output_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : _zz_io_output_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : _zz_io_output_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : _zz_io_output_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : _zz_io_output_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : _zz_io_output_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : _zz_io_output_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : _zz_io_output_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : _zz_io_output_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : _zz_io_output_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : _zz_io_output_payload_opcode_string = "FCVT_X_X";
      default : _zz_io_output_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_format)
      FpuFormat_FLOAT : _zz_io_output_payload_format_string = "FLOAT ";
      FpuFormat_DOUBLE : _zz_io_output_payload_format_string = "DOUBLE";
      default : _zz_io_output_payload_format_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_io_output_payload_roundMode)
      FpuRoundMode_RNE : _zz_io_output_payload_roundMode_string = "RNE";
      FpuRoundMode_RTZ : _zz_io_output_payload_roundMode_string = "RTZ";
      FpuRoundMode_RDN : _zz_io_output_payload_roundMode_string = "RDN";
      FpuRoundMode_RUP : _zz_io_output_payload_roundMode_string = "RUP";
      FpuRoundMode_RMM : _zz_io_output_payload_roundMode_string = "RMM";
      default : _zz_io_output_payload_roundMode_string = "???";
    endcase
  end
  `endif

  assign locked = 1'b0;
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_0 = {io_inputs_1_valid,io_inputs_0_valid};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[3 : 2] | _zz_maskProposal_0_2[1 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign _zz_io_output_payload_opcode = (maskRouted_0 ? io_inputs_0_payload_opcode : io_inputs_1_payload_opcode);
  assign _zz_io_output_payload_format = (maskRouted_0 ? io_inputs_0_payload_format : io_inputs_1_payload_format);
  assign _zz_io_output_payload_roundMode = (maskRouted_0 ? io_inputs_0_payload_roundMode : io_inputs_1_payload_roundMode);
  assign io_output_payload_opcode = _zz_io_output_payload_opcode;
  assign io_output_payload_arg = (maskRouted_0 ? io_inputs_0_payload_arg : io_inputs_1_payload_arg);
  assign io_output_payload_rs1 = (maskRouted_0 ? io_inputs_0_payload_rs1 : io_inputs_1_payload_rs1);
  assign io_output_payload_rs2 = (maskRouted_0 ? io_inputs_0_payload_rs2 : io_inputs_1_payload_rs2);
  assign io_output_payload_rs3 = (maskRouted_0 ? io_inputs_0_payload_rs3 : io_inputs_1_payload_rs3);
  assign io_output_payload_rd = (maskRouted_0 ? io_inputs_0_payload_rd : io_inputs_1_payload_rd);
  assign io_output_payload_format = _zz_io_output_payload_format;
  assign io_output_payload_roundMode = _zz_io_output_payload_roundMode;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
      end
    end
  end


endmodule

//StreamFork_1 replaced by StreamFork

module StreamFork (
  input  wire          io_input_valid,
  output wire          io_input_ready,
  input  wire [3:0]    io_input_payload_opcode,
  input  wire [4:0]    io_input_payload_rd,
  input  wire          io_input_payload_write,
  input  wire [63:0]   io_input_payload_value,
  output wire          io_outputs_0_valid,
  input  wire          io_outputs_0_ready,
  output wire [3:0]    io_outputs_0_payload_opcode,
  output wire [4:0]    io_outputs_0_payload_rd,
  output wire          io_outputs_0_payload_write,
  output wire [63:0]   io_outputs_0_payload_value,
  output wire          io_outputs_1_valid,
  input  wire          io_outputs_1_ready,
  output wire [3:0]    io_outputs_1_payload_opcode,
  output wire [4:0]    io_outputs_1_payload_rd,
  output wire          io_outputs_1_payload_write,
  output wire [63:0]   io_outputs_1_payload_value
);
  localparam FpuOpcode_LOAD = 4'd0;
  localparam FpuOpcode_STORE = 4'd1;
  localparam FpuOpcode_MUL = 4'd2;
  localparam FpuOpcode_ADD = 4'd3;
  localparam FpuOpcode_FMA = 4'd4;
  localparam FpuOpcode_I2F = 4'd5;
  localparam FpuOpcode_F2I = 4'd6;
  localparam FpuOpcode_CMP = 4'd7;
  localparam FpuOpcode_DIV = 4'd8;
  localparam FpuOpcode_SQRT = 4'd9;
  localparam FpuOpcode_MIN_MAX = 4'd10;
  localparam FpuOpcode_SGNJ = 4'd11;
  localparam FpuOpcode_FMV_X_W = 4'd12;
  localparam FpuOpcode_FMV_W_X = 4'd13;
  localparam FpuOpcode_FCLASS = 4'd14;
  localparam FpuOpcode_FCVT_X_X = 4'd15;

  `ifndef SYNTHESIS
  reg [63:0] io_input_payload_opcode_string;
  reg [63:0] io_outputs_0_payload_opcode_string;
  reg [63:0] io_outputs_1_payload_opcode_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(io_input_payload_opcode)
      FpuOpcode_LOAD : io_input_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_input_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_input_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_input_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_input_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_input_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_input_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_input_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_input_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_input_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_input_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_input_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_input_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_input_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_input_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_input_payload_opcode_string = "FCVT_X_X";
      default : io_input_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_outputs_0_payload_opcode)
      FpuOpcode_LOAD : io_outputs_0_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_outputs_0_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_outputs_0_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_outputs_0_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_outputs_0_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_outputs_0_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_outputs_0_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_outputs_0_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_outputs_0_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_outputs_0_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_outputs_0_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_outputs_0_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_outputs_0_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_outputs_0_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_outputs_0_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_outputs_0_payload_opcode_string = "FCVT_X_X";
      default : io_outputs_0_payload_opcode_string = "????????";
    endcase
  end
  always @(*) begin
    case(io_outputs_1_payload_opcode)
      FpuOpcode_LOAD : io_outputs_1_payload_opcode_string = "LOAD    ";
      FpuOpcode_STORE : io_outputs_1_payload_opcode_string = "STORE   ";
      FpuOpcode_MUL : io_outputs_1_payload_opcode_string = "MUL     ";
      FpuOpcode_ADD : io_outputs_1_payload_opcode_string = "ADD     ";
      FpuOpcode_FMA : io_outputs_1_payload_opcode_string = "FMA     ";
      FpuOpcode_I2F : io_outputs_1_payload_opcode_string = "I2F     ";
      FpuOpcode_F2I : io_outputs_1_payload_opcode_string = "F2I     ";
      FpuOpcode_CMP : io_outputs_1_payload_opcode_string = "CMP     ";
      FpuOpcode_DIV : io_outputs_1_payload_opcode_string = "DIV     ";
      FpuOpcode_SQRT : io_outputs_1_payload_opcode_string = "SQRT    ";
      FpuOpcode_MIN_MAX : io_outputs_1_payload_opcode_string = "MIN_MAX ";
      FpuOpcode_SGNJ : io_outputs_1_payload_opcode_string = "SGNJ    ";
      FpuOpcode_FMV_X_W : io_outputs_1_payload_opcode_string = "FMV_X_W ";
      FpuOpcode_FMV_W_X : io_outputs_1_payload_opcode_string = "FMV_W_X ";
      FpuOpcode_FCLASS : io_outputs_1_payload_opcode_string = "FCLASS  ";
      FpuOpcode_FCVT_X_X : io_outputs_1_payload_opcode_string = "FCVT_X_X";
      default : io_outputs_1_payload_opcode_string = "????????";
    endcase
  end
  `endif

  assign io_input_ready = (io_outputs_0_ready && io_outputs_1_ready);
  assign io_outputs_0_valid = (io_input_valid && io_input_ready);
  assign io_outputs_1_valid = (io_input_valid && io_input_ready);
  assign io_outputs_0_payload_opcode = io_input_payload_opcode;
  assign io_outputs_0_payload_rd = io_input_payload_rd;
  assign io_outputs_0_payload_write = io_input_payload_write;
  assign io_outputs_0_payload_value = io_input_payload_value;
  assign io_outputs_1_payload_opcode = io_input_payload_opcode;
  assign io_outputs_1_payload_rd = io_input_payload_rd;
  assign io_outputs_1_payload_write = io_input_payload_write;
  assign io_outputs_1_payload_value = io_input_payload_value;

endmodule

//BufferCC_1 replaced by BufferCC

//DataCache_1 replaced by DataCache

//InstructionCache_1 replaced by InstructionCache

module BufferCC (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

module DataCache (
  input  wire          io_cpu_execute_isValid,
  input  wire [31:0]   io_cpu_execute_address,
  output reg           io_cpu_execute_haltIt,
  input  wire          io_cpu_execute_args_wr,
  input  wire [1:0]    io_cpu_execute_args_size,
  input  wire          io_cpu_execute_args_isLrsc,
  input  wire          io_cpu_execute_args_isAmo,
  input  wire          io_cpu_execute_args_amoCtrl_swap,
  input  wire [2:0]    io_cpu_execute_args_amoCtrl_alu,
  input  wire          io_cpu_execute_args_totalyConsistent,
  output wire          io_cpu_execute_refilling,
  input  wire          io_cpu_memory_isValid,
  input  wire          io_cpu_memory_isStuck,
  output wire          io_cpu_memory_isWrite,
  input  wire [31:0]   io_cpu_memory_address,
  input  wire [31:0]   io_cpu_memory_mmuRsp_physicalAddress,
  input  wire          io_cpu_memory_mmuRsp_isIoAccess,
  input  wire          io_cpu_memory_mmuRsp_isPaging,
  input  wire          io_cpu_memory_mmuRsp_allowRead,
  input  wire          io_cpu_memory_mmuRsp_allowWrite,
  input  wire          io_cpu_memory_mmuRsp_allowExecute,
  input  wire          io_cpu_memory_mmuRsp_exception,
  input  wire          io_cpu_memory_mmuRsp_refilling,
  input  wire          io_cpu_memory_mmuRsp_bypassTranslation,
  input  wire          io_cpu_writeBack_isValid,
  input  wire          io_cpu_writeBack_isStuck,
  input  wire          io_cpu_writeBack_isFiring,
  input  wire          io_cpu_writeBack_isUser,
  output reg           io_cpu_writeBack_haltIt,
  output wire          io_cpu_writeBack_isWrite,
  input  wire [63:0]   io_cpu_writeBack_storeData,
  output reg  [63:0]   io_cpu_writeBack_data,
  input  wire [31:0]   io_cpu_writeBack_address,
  output wire          io_cpu_writeBack_mmuException,
  output wire          io_cpu_writeBack_unalignedAccess,
  output reg           io_cpu_writeBack_accessError,
  output reg           io_cpu_writeBack_keepMemRspData,
  input  wire          io_cpu_writeBack_fence_SW,
  input  wire          io_cpu_writeBack_fence_SR,
  input  wire          io_cpu_writeBack_fence_SO,
  input  wire          io_cpu_writeBack_fence_SI,
  input  wire          io_cpu_writeBack_fence_PW,
  input  wire          io_cpu_writeBack_fence_PR,
  input  wire          io_cpu_writeBack_fence_PO,
  input  wire          io_cpu_writeBack_fence_PI,
  input  wire [3:0]    io_cpu_writeBack_fence_FM,
  output wire          io_cpu_writeBack_exclusiveOk,
  output reg           io_cpu_redo,
  input  wire          io_cpu_flush_valid,
  output wire          io_cpu_flush_ready,
  input  wire          io_cpu_flush_payload_singleLine,
  input  wire [5:0]    io_cpu_flush_payload_lineId,
  output wire          io_cpu_writesPending,
  output reg           io_mem_cmd_valid,
  input  wire          io_mem_cmd_ready,
  output reg           io_mem_cmd_payload_wr,
  output wire          io_mem_cmd_payload_uncached,
  output reg  [31:0]   io_mem_cmd_payload_address,
  output wire [63:0]   io_mem_cmd_payload_data,
  output wire [7:0]    io_mem_cmd_payload_mask,
  output reg  [2:0]    io_mem_cmd_payload_size,
  output wire          io_mem_cmd_payload_exclusive,
  output wire          io_mem_cmd_payload_last,
  input  wire          io_mem_rsp_valid,
  input  wire [3:0]    io_mem_rsp_payload_aggregated,
  input  wire          io_mem_rsp_payload_last,
  input  wire [63:0]   io_mem_rsp_payload_data,
  input  wire          io_mem_rsp_payload_error,
  input  wire          io_mem_rsp_payload_exclusive,
  input  wire          io_mem_inv_valid,
  output reg           io_mem_inv_ready,
  input  wire          io_mem_inv_payload_last,
  input  wire          io_mem_inv_payload_fragment_enable,
  input  wire [31:0]   io_mem_inv_payload_fragment_address,
  output wire          io_mem_ack_valid,
  input  wire          io_mem_ack_ready,
  output wire          io_mem_ack_payload_last,
  output wire          io_mem_ack_payload_fragment_hit,
  input  wire          io_mem_sync_valid,
  output wire          io_mem_sync_ready,
  input  wire [3:0]    io_mem_sync_payload_aggregated,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);
  localparam DataCacheExternalAmoStates_LR_CMD = 2'd0;
  localparam DataCacheExternalAmoStates_LR_RSP = 2'd1;
  localparam DataCacheExternalAmoStates_SC_CMD = 2'd2;
  localparam DataCacheExternalAmoStates_SC_RSP = 2'd3;

  reg        [21:0]   ways_0_tags_spinal_port0;
  reg        [21:0]   ways_0_tags_spinal_port1;
  reg        [63:0]   ways_0_data_spinal_port0;
  reg        [21:0]   ways_1_tags_spinal_port0;
  reg        [21:0]   ways_1_tags_spinal_port1;
  reg        [63:0]   ways_1_data_spinal_port0;
  wire       [0:0]    sync_syncContext_history_spinal_port1;
  wire       [21:0]   _zz_ways_0_tags_port;
  wire       [21:0]   _zz_ways_1_tags_port;
  wire       [6:0]    _zz_pending_counterNext;
  wire       [6:0]    _zz_pending_counterNext_1;
  wire       [0:0]    _zz_pending_counterNext_2;
  wire       [6:0]    _zz_pending_counterNext_3;
  wire       [4:0]    _zz_pending_counterNext_4;
  wire       [4:0]    _zz_pending_counterNext_5;
  wire       [4:0]    _zz_pending_counterNext_6;
  wire       [1:0]    _zz_pending_counterNext_7;
  wire       [4:0]    _zz_sync_syncCount;
  wire       [1:0]    _zz_sync_syncCount_1;
  wire       [5:0]    _zz_sync_syncContext_history_port;
  wire       [0:0]    _zz_sync_syncContext_history_port_1;
  wire       [6:0]    _zz_sync_syncContext_rPtr;
  wire       [5:0]    _zz_sync_syncContext_history_port_2;
  wire       [5:0]    _zz_sync_syncContext_uncached_1;
  wire       [6:0]    _zz_sync_syncContext_full;
  wire       [6:0]    _zz_sync_writeCached_pendingSyncNext;
  wire       [6:0]    _zz_sync_writeCached_pendingSyncNext_1;
  wire       [0:0]    _zz_sync_writeCached_pendingSyncNext_2;
  wire       [6:0]    _zz_sync_writeCached_pendingSyncNext_3;
  wire       [4:0]    _zz_sync_writeCached_pendingSyncNext_4;
  wire       [6:0]    _zz_sync_writeUncached_pendingSyncNext;
  wire       [6:0]    _zz_sync_writeUncached_pendingSyncNext_1;
  wire       [0:0]    _zz_sync_writeUncached_pendingSyncNext_2;
  wire       [6:0]    _zz_sync_writeUncached_pendingSyncNext_3;
  wire       [4:0]    _zz_sync_writeUncached_pendingSyncNext_4;
  wire       [6:0]    _zz_sync_w2w_counter;
  wire       [4:0]    _zz_sync_w2w_counter_1;
  wire       [6:0]    _zz_sync_w2r_counter;
  wire       [4:0]    _zz_sync_w2r_counter_1;
  wire       [6:0]    _zz_sync_w2i_counter;
  wire       [4:0]    _zz_sync_w2i_counter_1;
  wire       [6:0]    _zz_sync_w2o_counter;
  wire       [4:0]    _zz_sync_w2o_counter_1;
  wire       [6:0]    _zz_sync_o2w_counter;
  wire       [4:0]    _zz_sync_o2w_counter_1;
  wire       [6:0]    _zz_sync_o2r_counter;
  wire       [4:0]    _zz_sync_o2r_counter_1;
  wire       [31:0]   _zz_stageB_amo_addSub;
  wire       [31:0]   _zz_stageB_amo_addSub_1;
  wire       [31:0]   _zz_stageB_amo_addSub_2;
  wire       [31:0]   _zz_stageB_amo_addSub_3;
  reg        [31:0]   _zz_stageB_amo_addSub_4;
  wire       [0:0]    _zz_stageB_amo_addSub_5;
  reg        [31:0]   _zz_stageB_amo_addSub_6;
  wire       [0:0]    _zz_stageB_amo_addSub_7;
  wire       [31:0]   _zz_stageB_amo_addSub_8;
  wire       [1:0]    _zz_stageB_amo_addSub_9;
  reg        [31:0]   _zz_stageB_amo_less;
  wire       [0:0]    _zz_stageB_amo_less_1;
  reg        [31:0]   _zz_stageB_amo_less_2;
  wire       [0:0]    _zz_stageB_amo_less_3;
  reg        [31:0]   _zz_stageB_amo_result;
  wire       [0:0]    _zz_stageB_amo_result_1;
  reg        [31:0]   _zz_stageB_amo_result_2;
  wire       [0:0]    _zz_stageB_amo_result_3;
  reg        [31:0]   _zz_stageB_amo_result_4;
  wire       [0:0]    _zz_stageB_amo_result_5;
  reg        [31:0]   _zz_stageB_amo_result_6;
  wire       [0:0]    _zz_stageB_amo_result_7;
  wire       [0:0]    _zz_when;
  wire       [2:0]    _zz_loader_counter_valueNext;
  wire       [0:0]    _zz_loader_counter_valueNext_1;
  wire       [2:0]    _zz_loader_waysAllocator;
  reg        [1:0]    invalidate_s1_wayHits_1;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 _zz_3;
  reg                 _zz_4;
  reg                 _zz_5;
  wire                haltCpu;
  reg                 tagsReadCmd_valid;
  reg        [5:0]    tagsReadCmd_payload;
  wire                tagsInvReadCmd_valid;
  wire       [5:0]    tagsInvReadCmd_payload;
  reg                 tagsWriteCmd_valid;
  reg        [1:0]    tagsWriteCmd_payload_way;
  reg        [5:0]    tagsWriteCmd_payload_address;
  reg                 tagsWriteCmd_payload_data_valid;
  reg                 tagsWriteCmd_payload_data_error;
  reg        [19:0]   tagsWriteCmd_payload_data_address;
  reg                 tagsWriteLastCmd_valid;
  reg        [1:0]    tagsWriteLastCmd_payload_way;
  reg        [5:0]    tagsWriteLastCmd_payload_address;
  reg                 tagsWriteLastCmd_payload_data_valid;
  reg                 tagsWriteLastCmd_payload_data_error;
  reg        [19:0]   tagsWriteLastCmd_payload_data_address;
  reg                 dataReadCmd_valid;
  reg        [8:0]    dataReadCmd_payload;
  reg                 dataWriteCmd_valid;
  reg        [1:0]    dataWriteCmd_payload_way;
  reg        [8:0]    dataWriteCmd_payload_address;
  reg        [63:0]   dataWriteCmd_payload_data;
  reg        [7:0]    dataWriteCmd_payload_mask;
  wire                _zz_ways_0_tagsReadRsp_valid;
  wire                ways_0_tagsReadRsp_valid;
  wire                ways_0_tagsReadRsp_error;
  wire       [19:0]   ways_0_tagsReadRsp_address;
  wire       [21:0]   _zz_ways_0_tagsReadRsp_valid_1;
  wire                _zz_ways_0_dataReadRspMem;
  wire       [63:0]   ways_0_dataReadRspMem;
  wire       [63:0]   ways_0_dataReadRsp;
  wire                ways_0_tagsInvReadRsp_valid;
  wire                ways_0_tagsInvReadRsp_error;
  wire       [19:0]   ways_0_tagsInvReadRsp_address;
  wire       [21:0]   _zz_ways_0_tagsInvReadRsp_valid;
  wire                when_DataCache_l645;
  wire                when_DataCache_l648;
  wire                _zz_ways_1_tagsReadRsp_valid;
  wire                ways_1_tagsReadRsp_valid;
  wire                ways_1_tagsReadRsp_error;
  wire       [19:0]   ways_1_tagsReadRsp_address;
  wire       [21:0]   _zz_ways_1_tagsReadRsp_valid_1;
  wire                _zz_ways_1_dataReadRspMem;
  wire       [63:0]   ways_1_dataReadRspMem;
  wire       [63:0]   ways_1_dataReadRsp;
  wire                ways_1_tagsInvReadRsp_valid;
  wire                ways_1_tagsInvReadRsp_error;
  wire       [19:0]   ways_1_tagsInvReadRsp_address;
  wire       [21:0]   _zz_ways_1_tagsInvReadRsp_valid;
  wire                when_DataCache_l645_1;
  wire                when_DataCache_l648_1;
  wire                when_DataCache_l667;
  reg                 rspSync;
  reg                 rspLast;
  reg                 memCmdSent;
  wire                io_mem_cmd_fire;
  wire                when_DataCache_l689;
  reg        [6:0]    pending_counter;
  wire       [6:0]    pending_counterNext;
  reg                 pending_done;
  reg                 pending_full;
  reg                 pending_last;
  wire                when_DataCache_l703;
  wire                when_DataCache_l704;
  wire       [4:0]    sync_syncCount;
  reg        [6:0]    sync_syncContext_wPtr;
  reg        [6:0]    sync_syncContext_rPtr;
  wire                when_DataCache_l713;
  wire                io_mem_sync_fire;
  wire       [6:0]    _zz_sync_syncContext_uncached;
  wire                sync_syncContext_uncached;
  reg                 sync_syncContext_full;
  wire                sync_syncContext_empty;
  reg        [6:0]    sync_writeCached_pendingSync;
  wire       [6:0]    sync_writeCached_pendingSyncNext;
  reg        [6:0]    sync_writeUncached_pendingSync;
  wire       [6:0]    sync_writeUncached_pendingSyncNext;
  wire                when_DataCache_l740;
  reg        [6:0]    sync_w2w_counter;
  wire                sync_w2w_busy;
  wire                when_DataCache_l740_1;
  reg        [6:0]    sync_w2r_counter;
  wire                sync_w2r_busy;
  wire                when_DataCache_l740_2;
  reg        [6:0]    sync_w2i_counter;
  wire                sync_w2i_busy;
  wire                when_DataCache_l740_3;
  reg        [6:0]    sync_w2o_counter;
  wire                sync_w2o_busy;
  wire                when_DataCache_l740_4;
  reg        [6:0]    sync_o2w_counter;
  wire                sync_o2w_busy;
  wire                when_DataCache_l740_5;
  reg        [6:0]    sync_o2r_counter;
  wire                sync_o2r_busy;
  wire                sync_notTotalyConsistent;
  reg        [7:0]    _zz_stage0_mask;
  wire       [7:0]    stage0_mask;
  reg        [1:0]    stage0_dataColisions;
  wire       [8:0]    _zz_stage0_dataColisions;
  wire       [7:0]    _zz_stage0_dataColisions_1;
  reg        [1:0]    stage0_wayInvalidate;
  wire                when_DataCache_l776;
  reg                 stageA_request_wr;
  reg        [1:0]    stageA_request_size;
  reg                 stageA_request_isLrsc;
  reg                 stageA_request_isAmo;
  reg                 stageA_request_amoCtrl_swap;
  reg        [2:0]    stageA_request_amoCtrl_alu;
  reg                 stageA_request_totalyConsistent;
  wire                when_DataCache_l776_1;
  reg        [7:0]    stageA_mask;
  reg                 stageA_consistancyCheck_hazard;
  wire                stageA_consistancyCheck_w;
  wire                when_DataCache_l776_2;
  reg                 _zz_stageA_consistancyCheck_r;
  wire                stageA_consistancyCheck_r;
  wire                stageA_consistancyCheck_o;
  wire                stageA_consistancyCheck_i;
  wire                stageA_consistancyCheck_s;
  wire                stageA_consistancyCheck_l;
  wire                when_DataCache_l793;
  wire                when_DataCache_l796;
  wire       [1:0]    stageA_wayHits;
  wire                when_DataCache_l776_3;
  reg        [1:0]    stageA_wayInvalidate;
  wire                when_DataCache_l776_4;
  reg        [1:0]    stage0_dataColisions_regNextWhen;
  reg        [1:0]    _zz_stageA_dataColisions;
  wire       [8:0]    _zz_stageA_dataColisions_1;
  wire       [7:0]    _zz_stageA_dataColisions_2;
  wire       [1:0]    stageA_dataColisions;
  wire                when_DataCache_l827;
  reg                 stageB_request_wr;
  reg        [1:0]    stageB_request_size;
  reg                 stageB_request_isLrsc;
  reg                 stageB_request_isAmo;
  reg                 stageB_request_amoCtrl_swap;
  reg        [2:0]    stageB_request_amoCtrl_alu;
  reg                 stageB_request_totalyConsistent;
  reg                 stageB_mmuRspFreeze;
  wire                when_DataCache_l829;
  reg        [31:0]   stageB_mmuRsp_physicalAddress;
  reg                 stageB_mmuRsp_isIoAccess;
  reg                 stageB_mmuRsp_isPaging;
  reg                 stageB_mmuRsp_allowRead;
  reg                 stageB_mmuRsp_allowWrite;
  reg                 stageB_mmuRsp_allowExecute;
  reg                 stageB_mmuRsp_exception;
  reg                 stageB_mmuRsp_refilling;
  reg                 stageB_mmuRsp_bypassTranslation;
  wire                when_DataCache_l826;
  reg                 stageB_tagsReadRsp_0_valid;
  reg                 stageB_tagsReadRsp_0_error;
  reg        [19:0]   stageB_tagsReadRsp_0_address;
  wire                when_DataCache_l826_1;
  reg                 stageB_tagsReadRsp_1_valid;
  reg                 stageB_tagsReadRsp_1_error;
  reg        [19:0]   stageB_tagsReadRsp_1_address;
  wire                when_DataCache_l826_2;
  reg        [63:0]   stageB_dataReadRsp_0;
  wire                when_DataCache_l826_3;
  reg        [63:0]   stageB_dataReadRsp_1;
  wire                when_DataCache_l825;
  reg        [1:0]    stageB_wayInvalidate;
  wire                when_DataCache_l825_1;
  reg                 stageB_consistancyHazard;
  wire                when_DataCache_l825_2;
  reg        [1:0]    stageB_dataColisions;
  wire                when_DataCache_l825_3;
  reg                 stageB_unaligned;
  wire                when_DataCache_l825_4;
  reg        [1:0]    stageB_waysHitsBeforeInvalidate;
  wire       [1:0]    stageB_waysHits;
  wire                stageB_waysHit;
  wire       [63:0]   stageB_dataMux;
  wire                when_DataCache_l825_5;
  reg        [7:0]    stageB_mask;
  reg                 stageB_loaderValid;
  wire       [63:0]   stageB_ioMemRspMuxed;
  reg                 stageB_flusher_waitDone;
  reg                 stageB_flusher_hold;
  reg        [6:0]    stageB_flusher_counter;
  wire                when_DataCache_l855;
  wire                when_DataCache_l861;
  wire                when_DataCache_l863;
  reg                 stageB_flusher_start;
  wire                when_DataCache_l877;
  wire                stageB_isAmoCached;
  reg        [63:0]   stageB_requestDataBypass;
  wire                stageB_amo_compare;
  wire                stageB_amo_unsigned;
  wire       [31:0]   stageB_amo_addSub;
  wire                stageB_amo_less;
  wire                stageB_amo_selectRf;
  wire       [2:0]    switch_Misc_l241;
  reg        [31:0]   stageB_amo_result;
  reg        [31:0]   stageB_amo_resultReg;
  reg        [1:0]    stageB_amo_external_state;
  reg                 stageB_cpuWriteToCache;
  wire                when_DataCache_l931;
  wire                stageB_badPermissions;
  wire                stageB_loadStoreFault;
  wire                stageB_bypassCache;
  wire                when_DataCache_l974;
  reg                 _zz_when_DataCache_l1000;
  wire                when_DataCache_l1000;
  wire                when_DataCache_l1009;
  wire                when_DataCache_l1014;
  wire                when_DataCache_l1025;
  wire                when_DataCache_l1037;
  wire                when_DataCache_l996;
  wire                when_DataCache_l1059;
  wire                when_DataCache_l1061;
  wire                when_DataCache_l1072;
  wire                when_DataCache_l1081;
  reg                 loader_valid;
  reg                 loader_counter_willIncrement;
  wire                loader_counter_willClear;
  reg        [2:0]    loader_counter_valueNext;
  reg        [2:0]    loader_counter_value;
  wire                loader_counter_willOverflowIfInc;
  wire                loader_counter_willOverflow;
  reg        [1:0]    loader_waysAllocator;
  reg                 loader_error;
  reg                 loader_kill;
  reg                 loader_killReg;
  wire                when_DataCache_l1097;
  reg                 loader_done;
  wire                when_DataCache_l1108;
  wire                when_DataCache_l1125;
  reg                 loader_valid_regNext;
  wire                when_DataCache_l1129;
  wire                when_DataCache_l1132;
  wire                io_mem_inv_fire;
  wire                invalidate_s0_loaderTagHit;
  wire                invalidate_s0_loaderLineHit;
  wire                when_DataCache_l1143;
  wire                invalidate_s1_input_valid;
  reg                 invalidate_s1_input_ready;
  wire                invalidate_s1_input_payload_last;
  wire                invalidate_s1_input_payload_fragment_enable;
  wire       [31:0]   invalidate_s1_input_payload_fragment_address;
  reg                 io_mem_inv_rValid;
  reg                 io_mem_inv_rData_last;
  reg                 io_mem_inv_rData_fragment_enable;
  reg        [31:0]   io_mem_inv_rData_fragment_address;
  wire                when_Stream_l375;
  reg                 invalidate_s1_loaderValid;
  reg        [1:0]    invalidate_s1_loaderWay;
  reg                 invalidate_s1_loaderTagHit;
  reg                 invalidate_s1_loaderLineHit;
  wire       [1:0]    invalidate_s1_invalidations;
  wire       [1:0]    invalidate_s1_wayHits;
  wire                when_DataCache_l1158;
  wire                invalidate_s2_input_valid;
  wire                invalidate_s2_input_ready;
  wire                invalidate_s2_input_payload_last;
  wire                invalidate_s2_input_payload_fragment_enable;
  wire       [31:0]   invalidate_s2_input_payload_fragment_address;
  reg                 invalidate_s1_input_rValid;
  reg                 invalidate_s1_input_rData_last;
  reg                 invalidate_s1_input_rData_fragment_enable;
  reg        [31:0]   invalidate_s1_input_rData_fragment_address;
  wire                when_Stream_l375_1;
  reg        [1:0]    invalidate_s2_wayHits;
  wire                invalidate_s2_wayHit;
  wire                when_DataCache_l1167;
  wire                when_DataCache_l1169;
  reg        [1:0]    _zz_invalidate_s1_invalidations;
  `ifndef SYNTHESIS
  reg [47:0] stageB_amo_external_state_string;
  `endif

  reg [21:0] ways_0_tags [0:63];
  reg [7:0] ways_0_data_symbol0 [0:511];
  reg [7:0] ways_0_data_symbol1 [0:511];
  reg [7:0] ways_0_data_symbol2 [0:511];
  reg [7:0] ways_0_data_symbol3 [0:511];
  reg [7:0] ways_0_data_symbol4 [0:511];
  reg [7:0] ways_0_data_symbol5 [0:511];
  reg [7:0] ways_0_data_symbol6 [0:511];
  reg [7:0] ways_0_data_symbol7 [0:511];
  reg [7:0] _zz_ways_0_datasymbol_read;
  reg [7:0] _zz_ways_0_datasymbol_read_1;
  reg [7:0] _zz_ways_0_datasymbol_read_2;
  reg [7:0] _zz_ways_0_datasymbol_read_3;
  reg [7:0] _zz_ways_0_datasymbol_read_4;
  reg [7:0] _zz_ways_0_datasymbol_read_5;
  reg [7:0] _zz_ways_0_datasymbol_read_6;
  reg [7:0] _zz_ways_0_datasymbol_read_7;
  reg [21:0] ways_1_tags [0:63];
  reg [7:0] ways_1_data_symbol0 [0:511];
  reg [7:0] ways_1_data_symbol1 [0:511];
  reg [7:0] ways_1_data_symbol2 [0:511];
  reg [7:0] ways_1_data_symbol3 [0:511];
  reg [7:0] ways_1_data_symbol4 [0:511];
  reg [7:0] ways_1_data_symbol5 [0:511];
  reg [7:0] ways_1_data_symbol6 [0:511];
  reg [7:0] ways_1_data_symbol7 [0:511];
  reg [7:0] _zz_ways_1_datasymbol_read;
  reg [7:0] _zz_ways_1_datasymbol_read_1;
  reg [7:0] _zz_ways_1_datasymbol_read_2;
  reg [7:0] _zz_ways_1_datasymbol_read_3;
  reg [7:0] _zz_ways_1_datasymbol_read_4;
  reg [7:0] _zz_ways_1_datasymbol_read_5;
  reg [7:0] _zz_ways_1_datasymbol_read_6;
  reg [7:0] _zz_ways_1_datasymbol_read_7;
  (* ram_style = "distributed" *) reg [0:0] sync_syncContext_history [0:63];

  assign _zz_pending_counterNext = (pending_counter + _zz_pending_counterNext_1);
  assign _zz_pending_counterNext_2 = (io_mem_cmd_fire && io_mem_cmd_payload_last);
  assign _zz_pending_counterNext_1 = {6'd0, _zz_pending_counterNext_2};
  assign _zz_pending_counterNext_4 = ((io_mem_rsp_valid && io_mem_rsp_payload_last) ? _zz_pending_counterNext_5 : 5'h0);
  assign _zz_pending_counterNext_3 = {2'd0, _zz_pending_counterNext_4};
  assign _zz_pending_counterNext_5 = ({1'b0,io_mem_rsp_payload_aggregated} + _zz_pending_counterNext_6);
  assign _zz_pending_counterNext_7 = {1'b0,1'b1};
  assign _zz_pending_counterNext_6 = {3'd0, _zz_pending_counterNext_7};
  assign _zz_sync_syncCount_1 = {1'b0,1'b1};
  assign _zz_sync_syncCount = {3'd0, _zz_sync_syncCount_1};
  assign _zz_sync_syncContext_history_port = sync_syncContext_wPtr[5:0];
  assign _zz_sync_syncContext_rPtr = {2'd0, sync_syncCount};
  assign _zz_sync_syncContext_uncached_1 = _zz_sync_syncContext_uncached[5:0];
  assign _zz_sync_syncContext_full = (sync_syncContext_wPtr - sync_syncContext_rPtr);
  assign _zz_sync_writeCached_pendingSyncNext = (sync_writeCached_pendingSync + _zz_sync_writeCached_pendingSyncNext_1);
  assign _zz_sync_writeCached_pendingSyncNext_2 = ((io_mem_cmd_fire && io_mem_cmd_payload_wr) && (! io_mem_cmd_payload_uncached));
  assign _zz_sync_writeCached_pendingSyncNext_1 = {6'd0, _zz_sync_writeCached_pendingSyncNext_2};
  assign _zz_sync_writeCached_pendingSyncNext_4 = ((io_mem_sync_fire && (! sync_syncContext_uncached)) ? sync_syncCount : 5'h0);
  assign _zz_sync_writeCached_pendingSyncNext_3 = {2'd0, _zz_sync_writeCached_pendingSyncNext_4};
  assign _zz_sync_writeUncached_pendingSyncNext = (sync_writeUncached_pendingSync + _zz_sync_writeUncached_pendingSyncNext_1);
  assign _zz_sync_writeUncached_pendingSyncNext_2 = ((io_mem_cmd_fire && io_mem_cmd_payload_wr) && io_mem_cmd_payload_uncached);
  assign _zz_sync_writeUncached_pendingSyncNext_1 = {6'd0, _zz_sync_writeUncached_pendingSyncNext_2};
  assign _zz_sync_writeUncached_pendingSyncNext_4 = ((io_mem_sync_fire && sync_syncContext_uncached) ? sync_syncCount : 5'h0);
  assign _zz_sync_writeUncached_pendingSyncNext_3 = {2'd0, _zz_sync_writeUncached_pendingSyncNext_4};
  assign _zz_sync_w2w_counter_1 = (((io_mem_sync_fire && (sync_w2w_counter != 7'h0)) && (! sync_syncContext_uncached)) ? sync_syncCount : 5'h0);
  assign _zz_sync_w2w_counter = {2'd0, _zz_sync_w2w_counter_1};
  assign _zz_sync_w2r_counter_1 = (((io_mem_sync_fire && (sync_w2r_counter != 7'h0)) && (! sync_syncContext_uncached)) ? sync_syncCount : 5'h0);
  assign _zz_sync_w2r_counter = {2'd0, _zz_sync_w2r_counter_1};
  assign _zz_sync_w2i_counter_1 = (((io_mem_sync_fire && (sync_w2i_counter != 7'h0)) && (! sync_syncContext_uncached)) ? sync_syncCount : 5'h0);
  assign _zz_sync_w2i_counter = {2'd0, _zz_sync_w2i_counter_1};
  assign _zz_sync_w2o_counter_1 = (((io_mem_sync_fire && (sync_w2o_counter != 7'h0)) && (! sync_syncContext_uncached)) ? sync_syncCount : 5'h0);
  assign _zz_sync_w2o_counter = {2'd0, _zz_sync_w2o_counter_1};
  assign _zz_sync_o2w_counter_1 = (((io_mem_sync_fire && (sync_o2w_counter != 7'h0)) && sync_syncContext_uncached) ? sync_syncCount : 5'h0);
  assign _zz_sync_o2w_counter = {2'd0, _zz_sync_o2w_counter_1};
  assign _zz_sync_o2r_counter_1 = (((io_mem_sync_fire && (sync_o2r_counter != 7'h0)) && sync_syncContext_uncached) ? sync_syncCount : 5'h0);
  assign _zz_sync_o2r_counter = {2'd0, _zz_sync_o2r_counter_1};
  assign _zz_stageB_amo_addSub = ($signed(_zz_stageB_amo_addSub_1) + $signed(_zz_stageB_amo_addSub_8));
  assign _zz_stageB_amo_addSub_1 = ($signed(_zz_stageB_amo_addSub_2) + $signed(_zz_stageB_amo_addSub_3));
  assign _zz_stageB_amo_addSub_2 = io_cpu_writeBack_storeData[31 : 0];
  assign _zz_stageB_amo_addSub_3 = (stageB_amo_compare ? (~ _zz_stageB_amo_addSub_4) : _zz_stageB_amo_addSub_6);
  assign _zz_stageB_amo_addSub_9 = (stageB_amo_compare ? 2'b01 : 2'b00);
  assign _zz_stageB_amo_addSub_8 = {{30{_zz_stageB_amo_addSub_9[1]}}, _zz_stageB_amo_addSub_9};
  assign _zz_when = 1'b1;
  assign _zz_loader_counter_valueNext_1 = loader_counter_willIncrement;
  assign _zz_loader_counter_valueNext = {2'd0, _zz_loader_counter_valueNext_1};
  assign _zz_loader_waysAllocator = {loader_waysAllocator,loader_waysAllocator[1]};
  assign _zz_ways_0_tags_port = {tagsWriteCmd_payload_data_address,{tagsWriteCmd_payload_data_error,tagsWriteCmd_payload_data_valid}};
  assign _zz_ways_1_tags_port = {tagsWriteCmd_payload_data_address,{tagsWriteCmd_payload_data_error,tagsWriteCmd_payload_data_valid}};
  assign _zz_sync_syncContext_history_port_1 = io_mem_cmd_payload_uncached;
  assign _zz_stageB_amo_addSub_5 = io_cpu_writeBack_address[2 : 2];
  assign _zz_stageB_amo_addSub_7 = io_cpu_writeBack_address[2 : 2];
  assign _zz_stageB_amo_less_1 = io_cpu_writeBack_address[2 : 2];
  assign _zz_stageB_amo_less_3 = io_cpu_writeBack_address[2 : 2];
  assign _zz_stageB_amo_result_1 = io_cpu_writeBack_address[2 : 2];
  assign _zz_stageB_amo_result_3 = io_cpu_writeBack_address[2 : 2];
  assign _zz_stageB_amo_result_5 = io_cpu_writeBack_address[2 : 2];
  assign _zz_stageB_amo_result_7 = io_cpu_writeBack_address[2 : 2];
  always @(posedge io_systemClk) begin
    if(_zz_ways_0_tagsReadRsp_valid) begin
      ways_0_tags_spinal_port0 <= ways_0_tags[tagsReadCmd_payload];
    end
  end

  always @(posedge io_systemClk) begin
    if(tagsInvReadCmd_valid) begin
      ways_0_tags_spinal_port1 <= ways_0_tags[tagsInvReadCmd_payload];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_5) begin
      ways_0_tags[tagsWriteCmd_payload_address] <= _zz_ways_0_tags_port;
    end
  end

  always @(*) begin
    ways_0_data_spinal_port0 = {_zz_ways_0_datasymbol_read_7, _zz_ways_0_datasymbol_read_6, _zz_ways_0_datasymbol_read_5, _zz_ways_0_datasymbol_read_4, _zz_ways_0_datasymbol_read_3, _zz_ways_0_datasymbol_read_2, _zz_ways_0_datasymbol_read_1, _zz_ways_0_datasymbol_read};
  end
  always @(posedge io_systemClk) begin
    if(_zz_ways_0_dataReadRspMem) begin
      _zz_ways_0_datasymbol_read <= ways_0_data_symbol0[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_1 <= ways_0_data_symbol1[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_2 <= ways_0_data_symbol2[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_3 <= ways_0_data_symbol3[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_4 <= ways_0_data_symbol4[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_5 <= ways_0_data_symbol5[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_6 <= ways_0_data_symbol6[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_7 <= ways_0_data_symbol7[dataReadCmd_payload];
    end
  end

  always @(posedge io_systemClk) begin
    if(dataWriteCmd_payload_mask[0] && _zz_4) begin
      ways_0_data_symbol0[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[7 : 0];
    end
    if(dataWriteCmd_payload_mask[1] && _zz_4) begin
      ways_0_data_symbol1[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[15 : 8];
    end
    if(dataWriteCmd_payload_mask[2] && _zz_4) begin
      ways_0_data_symbol2[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[23 : 16];
    end
    if(dataWriteCmd_payload_mask[3] && _zz_4) begin
      ways_0_data_symbol3[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[31 : 24];
    end
    if(dataWriteCmd_payload_mask[4] && _zz_4) begin
      ways_0_data_symbol4[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[39 : 32];
    end
    if(dataWriteCmd_payload_mask[5] && _zz_4) begin
      ways_0_data_symbol5[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[47 : 40];
    end
    if(dataWriteCmd_payload_mask[6] && _zz_4) begin
      ways_0_data_symbol6[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[55 : 48];
    end
    if(dataWriteCmd_payload_mask[7] && _zz_4) begin
      ways_0_data_symbol7[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[63 : 56];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_ways_1_tagsReadRsp_valid) begin
      ways_1_tags_spinal_port0 <= ways_1_tags[tagsReadCmd_payload];
    end
  end

  always @(posedge io_systemClk) begin
    if(tagsInvReadCmd_valid) begin
      ways_1_tags_spinal_port1 <= ways_1_tags[tagsInvReadCmd_payload];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_3) begin
      ways_1_tags[tagsWriteCmd_payload_address] <= _zz_ways_1_tags_port;
    end
  end

  always @(*) begin
    ways_1_data_spinal_port0 = {_zz_ways_1_datasymbol_read_7, _zz_ways_1_datasymbol_read_6, _zz_ways_1_datasymbol_read_5, _zz_ways_1_datasymbol_read_4, _zz_ways_1_datasymbol_read_3, _zz_ways_1_datasymbol_read_2, _zz_ways_1_datasymbol_read_1, _zz_ways_1_datasymbol_read};
  end
  always @(posedge io_systemClk) begin
    if(_zz_ways_1_dataReadRspMem) begin
      _zz_ways_1_datasymbol_read <= ways_1_data_symbol0[dataReadCmd_payload];
      _zz_ways_1_datasymbol_read_1 <= ways_1_data_symbol1[dataReadCmd_payload];
      _zz_ways_1_datasymbol_read_2 <= ways_1_data_symbol2[dataReadCmd_payload];
      _zz_ways_1_datasymbol_read_3 <= ways_1_data_symbol3[dataReadCmd_payload];
      _zz_ways_1_datasymbol_read_4 <= ways_1_data_symbol4[dataReadCmd_payload];
      _zz_ways_1_datasymbol_read_5 <= ways_1_data_symbol5[dataReadCmd_payload];
      _zz_ways_1_datasymbol_read_6 <= ways_1_data_symbol6[dataReadCmd_payload];
      _zz_ways_1_datasymbol_read_7 <= ways_1_data_symbol7[dataReadCmd_payload];
    end
  end

  always @(posedge io_systemClk) begin
    if(dataWriteCmd_payload_mask[0] && _zz_2) begin
      ways_1_data_symbol0[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[7 : 0];
    end
    if(dataWriteCmd_payload_mask[1] && _zz_2) begin
      ways_1_data_symbol1[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[15 : 8];
    end
    if(dataWriteCmd_payload_mask[2] && _zz_2) begin
      ways_1_data_symbol2[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[23 : 16];
    end
    if(dataWriteCmd_payload_mask[3] && _zz_2) begin
      ways_1_data_symbol3[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[31 : 24];
    end
    if(dataWriteCmd_payload_mask[4] && _zz_2) begin
      ways_1_data_symbol4[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[39 : 32];
    end
    if(dataWriteCmd_payload_mask[5] && _zz_2) begin
      ways_1_data_symbol5[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[47 : 40];
    end
    if(dataWriteCmd_payload_mask[6] && _zz_2) begin
      ways_1_data_symbol6[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[55 : 48];
    end
    if(dataWriteCmd_payload_mask[7] && _zz_2) begin
      ways_1_data_symbol7[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[63 : 56];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      sync_syncContext_history[_zz_sync_syncContext_history_port] <= _zz_sync_syncContext_history_port_1;
    end
  end

  assign sync_syncContext_history_spinal_port1 = sync_syncContext_history[_zz_sync_syncContext_uncached_1];
  always @(*) begin
    case(_zz_stageB_amo_addSub_5)
      1'b0 : _zz_stageB_amo_addSub_4 = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_addSub_4 = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_stageB_amo_addSub_7)
      1'b0 : _zz_stageB_amo_addSub_6 = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_addSub_6 = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_stageB_amo_less_1)
      1'b0 : _zz_stageB_amo_less = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_less = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_stageB_amo_less_3)
      1'b0 : _zz_stageB_amo_less_2 = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_less_2 = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_stageB_amo_result_1)
      1'b0 : _zz_stageB_amo_result = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_result = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_stageB_amo_result_3)
      1'b0 : _zz_stageB_amo_result_2 = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_result_2 = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_stageB_amo_result_5)
      1'b0 : _zz_stageB_amo_result_4 = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_result_4 = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_stageB_amo_result_7)
      1'b0 : _zz_stageB_amo_result_6 = stageB_ioMemRspMuxed[31 : 0];
      default : _zz_stageB_amo_result_6 = stageB_ioMemRspMuxed[63 : 32];
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(stageB_amo_external_state)
      DataCacheExternalAmoStates_LR_CMD : stageB_amo_external_state_string = "LR_CMD";
      DataCacheExternalAmoStates_LR_RSP : stageB_amo_external_state_string = "LR_RSP";
      DataCacheExternalAmoStates_SC_CMD : stageB_amo_external_state_string = "SC_CMD";
      DataCacheExternalAmoStates_SC_RSP : stageB_amo_external_state_string = "SC_RSP";
      default : stageB_amo_external_state_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    invalidate_s1_wayHits_1 = invalidate_s1_wayHits;
    if(when_DataCache_l1158) begin
      invalidate_s1_wayHits_1 = (invalidate_s1_wayHits & (~ invalidate_s1_loaderWay));
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(when_DataCache_l713) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(when_DataCache_l648_1) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(when_DataCache_l645_1) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(when_DataCache_l648) begin
      _zz_4 = 1'b1;
    end
  end

  always @(*) begin
    _zz_5 = 1'b0;
    if(when_DataCache_l645) begin
      _zz_5 = 1'b1;
    end
  end

  assign haltCpu = 1'b0;
  assign _zz_ways_0_tagsReadRsp_valid = (tagsReadCmd_valid && (! io_cpu_memory_isStuck));
  assign _zz_ways_0_tagsReadRsp_valid_1 = ways_0_tags_spinal_port0;
  assign ways_0_tagsReadRsp_valid = _zz_ways_0_tagsReadRsp_valid_1[0];
  assign ways_0_tagsReadRsp_error = _zz_ways_0_tagsReadRsp_valid_1[1];
  assign ways_0_tagsReadRsp_address = _zz_ways_0_tagsReadRsp_valid_1[21 : 2];
  assign _zz_ways_0_dataReadRspMem = (dataReadCmd_valid && (! io_cpu_memory_isStuck));
  assign ways_0_dataReadRspMem = ways_0_data_spinal_port0;
  assign ways_0_dataReadRsp = ways_0_dataReadRspMem[63 : 0];
  assign _zz_ways_0_tagsInvReadRsp_valid = ways_0_tags_spinal_port1;
  assign ways_0_tagsInvReadRsp_valid = _zz_ways_0_tagsInvReadRsp_valid[0];
  assign ways_0_tagsInvReadRsp_error = _zz_ways_0_tagsInvReadRsp_valid[1];
  assign ways_0_tagsInvReadRsp_address = _zz_ways_0_tagsInvReadRsp_valid[21 : 2];
  assign when_DataCache_l645 = (tagsWriteCmd_valid && tagsWriteCmd_payload_way[0]);
  assign when_DataCache_l648 = (dataWriteCmd_valid && dataWriteCmd_payload_way[0]);
  assign _zz_ways_1_tagsReadRsp_valid = (tagsReadCmd_valid && (! io_cpu_memory_isStuck));
  assign _zz_ways_1_tagsReadRsp_valid_1 = ways_1_tags_spinal_port0;
  assign ways_1_tagsReadRsp_valid = _zz_ways_1_tagsReadRsp_valid_1[0];
  assign ways_1_tagsReadRsp_error = _zz_ways_1_tagsReadRsp_valid_1[1];
  assign ways_1_tagsReadRsp_address = _zz_ways_1_tagsReadRsp_valid_1[21 : 2];
  assign _zz_ways_1_dataReadRspMem = (dataReadCmd_valid && (! io_cpu_memory_isStuck));
  assign ways_1_dataReadRspMem = ways_1_data_spinal_port0;
  assign ways_1_dataReadRsp = ways_1_dataReadRspMem[63 : 0];
  assign _zz_ways_1_tagsInvReadRsp_valid = ways_1_tags_spinal_port1;
  assign ways_1_tagsInvReadRsp_valid = _zz_ways_1_tagsInvReadRsp_valid[0];
  assign ways_1_tagsInvReadRsp_error = _zz_ways_1_tagsInvReadRsp_valid[1];
  assign ways_1_tagsInvReadRsp_address = _zz_ways_1_tagsInvReadRsp_valid[21 : 2];
  assign when_DataCache_l645_1 = (tagsWriteCmd_valid && tagsWriteCmd_payload_way[1]);
  assign when_DataCache_l648_1 = (dataWriteCmd_valid && dataWriteCmd_payload_way[1]);
  always @(*) begin
    tagsReadCmd_valid = 1'b0;
    if(when_DataCache_l667) begin
      tagsReadCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    tagsReadCmd_payload = 6'bxxxxxx;
    if(when_DataCache_l667) begin
      tagsReadCmd_payload = io_cpu_execute_address[11 : 6];
    end
  end

  always @(*) begin
    dataReadCmd_valid = 1'b0;
    if(when_DataCache_l667) begin
      dataReadCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    dataReadCmd_payload = 9'bxxxxxxxxx;
    if(when_DataCache_l667) begin
      dataReadCmd_payload = io_cpu_execute_address[11 : 3];
    end
  end

  always @(*) begin
    tagsWriteCmd_valid = 1'b0;
    if(when_DataCache_l855) begin
      tagsWriteCmd_valid = 1'b1;
    end
    if(io_cpu_writeBack_isValid) begin
      if(when_DataCache_l1072) begin
        tagsWriteCmd_valid = 1'b0;
      end
    end
    if(loader_done) begin
      tagsWriteCmd_valid = 1'b1;
    end
    if(when_DataCache_l1167) begin
      if(invalidate_s2_wayHit) begin
        tagsWriteCmd_valid = 1'b1;
      end
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_way = 2'bxx;
    if(when_DataCache_l855) begin
      tagsWriteCmd_payload_way = 2'b11;
    end
    if(loader_done) begin
      tagsWriteCmd_payload_way = loader_waysAllocator;
    end
    if(when_DataCache_l1167) begin
      if(invalidate_s2_wayHit) begin
        tagsWriteCmd_payload_way = invalidate_s2_wayHits;
      end
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_address = 6'bxxxxxx;
    if(when_DataCache_l855) begin
      tagsWriteCmd_payload_address = stageB_flusher_counter[5:0];
    end
    if(loader_done) begin
      tagsWriteCmd_payload_address = stageB_mmuRsp_physicalAddress[11 : 6];
    end
    if(when_DataCache_l1167) begin
      if(invalidate_s2_wayHit) begin
        tagsWriteCmd_payload_address = invalidate_s2_input_payload_fragment_address[11 : 6];
      end
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_data_valid = 1'bx;
    if(when_DataCache_l855) begin
      tagsWriteCmd_payload_data_valid = 1'b0;
    end
    if(loader_done) begin
      tagsWriteCmd_payload_data_valid = (! (loader_kill || loader_killReg));
    end
    if(when_DataCache_l1167) begin
      if(invalidate_s2_wayHit) begin
        tagsWriteCmd_payload_data_valid = 1'b0;
      end
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_data_error = 1'bx;
    if(loader_done) begin
      tagsWriteCmd_payload_data_error = (loader_error || (io_mem_rsp_valid && io_mem_rsp_payload_error));
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_data_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(loader_done) begin
      tagsWriteCmd_payload_data_address = stageB_mmuRsp_physicalAddress[31 : 12];
    end
  end

  always @(*) begin
    dataWriteCmd_valid = 1'b0;
    if(stageB_cpuWriteToCache) begin
      if(when_DataCache_l931) begin
        dataWriteCmd_valid = 1'b1;
      end
    end
    if(io_cpu_writeBack_isValid) begin
      if(when_DataCache_l1072) begin
        dataWriteCmd_valid = 1'b0;
      end
    end
    if(when_DataCache_l1097) begin
      dataWriteCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    dataWriteCmd_payload_way = 2'bxx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_way = stageB_waysHits;
    end
    if(when_DataCache_l1097) begin
      dataWriteCmd_payload_way = loader_waysAllocator;
    end
  end

  always @(*) begin
    dataWriteCmd_payload_address = 9'bxxxxxxxxx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_address = stageB_mmuRsp_physicalAddress[11 : 3];
    end
    if(when_DataCache_l1097) begin
      dataWriteCmd_payload_address = {stageB_mmuRsp_physicalAddress[11 : 6],loader_counter_value};
    end
  end

  always @(*) begin
    dataWriteCmd_payload_data = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_data[63 : 0] = stageB_requestDataBypass;
    end
    if(when_DataCache_l1097) begin
      dataWriteCmd_payload_data = io_mem_rsp_payload_data;
    end
  end

  always @(*) begin
    dataWriteCmd_payload_mask = 8'bxxxxxxxx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_mask = 8'h0;
      if(_zz_when[0]) begin
        dataWriteCmd_payload_mask[7 : 0] = stageB_mask;
      end
    end
    if(when_DataCache_l1097) begin
      dataWriteCmd_payload_mask = 8'hff;
    end
  end

  assign when_DataCache_l667 = (io_cpu_execute_isValid && (! io_cpu_memory_isStuck));
  always @(*) begin
    io_cpu_execute_haltIt = 1'b0;
    if(sync_syncContext_full) begin
      io_cpu_execute_haltIt = 1'b1;
    end
    if(when_DataCache_l855) begin
      io_cpu_execute_haltIt = 1'b1;
    end
  end

  always @(*) begin
    rspSync = 1'b1;
    if(when_DataCache_l703) begin
      rspSync = 1'b0;
    end
  end

  always @(*) begin
    rspLast = 1'b1;
    if(when_DataCache_l704) begin
      rspLast = 1'b0;
    end
  end

  assign io_mem_cmd_fire = (io_mem_cmd_valid && io_mem_cmd_ready);
  assign when_DataCache_l689 = (! io_cpu_writeBack_isStuck);
  assign pending_counterNext = (_zz_pending_counterNext - _zz_pending_counterNext_3);
  assign when_DataCache_l703 = ((! pending_last) || (! memCmdSent));
  assign when_DataCache_l704 = (! pending_last);
  assign io_mem_sync_ready = 1'b1;
  assign sync_syncCount = ({1'b0,io_mem_sync_payload_aggregated} + _zz_sync_syncCount);
  assign when_DataCache_l713 = (io_mem_cmd_fire && io_mem_cmd_payload_wr);
  assign io_mem_sync_fire = (io_mem_sync_valid && io_mem_sync_ready);
  assign _zz_sync_syncContext_uncached = sync_syncContext_rPtr;
  assign sync_syncContext_uncached = sync_syncContext_history_spinal_port1[0];
  assign sync_syncContext_empty = (sync_syncContext_wPtr == sync_syncContext_rPtr);
  assign io_cpu_writesPending = (! sync_syncContext_empty);
  assign sync_writeCached_pendingSyncNext = (_zz_sync_writeCached_pendingSyncNext - _zz_sync_writeCached_pendingSyncNext_3);
  assign sync_writeUncached_pendingSyncNext = (_zz_sync_writeUncached_pendingSyncNext - _zz_sync_writeUncached_pendingSyncNext_3);
  assign when_DataCache_l740 = (io_cpu_writeBack_fence_PW && io_cpu_writeBack_fence_SW);
  assign sync_w2w_busy = (sync_w2w_counter != 7'h0);
  assign when_DataCache_l740_1 = (io_cpu_writeBack_fence_PW && io_cpu_writeBack_fence_SR);
  assign sync_w2r_busy = (sync_w2r_counter != 7'h0);
  assign when_DataCache_l740_2 = (io_cpu_writeBack_fence_PW && io_cpu_writeBack_fence_SI);
  assign sync_w2i_busy = (sync_w2i_counter != 7'h0);
  assign when_DataCache_l740_3 = (io_cpu_writeBack_fence_PW && io_cpu_writeBack_fence_SO);
  assign sync_w2o_busy = (sync_w2o_counter != 7'h0);
  assign when_DataCache_l740_4 = (io_cpu_writeBack_fence_PO && io_cpu_writeBack_fence_SW);
  assign sync_o2w_busy = (sync_o2w_counter != 7'h0);
  assign when_DataCache_l740_5 = (io_cpu_writeBack_fence_PO && io_cpu_writeBack_fence_SR);
  assign sync_o2r_busy = (sync_o2r_counter != 7'h0);
  assign sync_notTotalyConsistent = (((((sync_w2w_busy || sync_w2r_busy) || sync_w2i_busy) || sync_w2o_busy) || sync_o2w_busy) || sync_o2r_busy);
  always @(*) begin
    _zz_stage0_mask = 8'bxxxxxxxx;
    case(io_cpu_execute_args_size)
      2'b00 : begin
        _zz_stage0_mask = 8'h01;
      end
      2'b01 : begin
        _zz_stage0_mask = 8'h03;
      end
      2'b10 : begin
        _zz_stage0_mask = 8'h0f;
      end
      default : begin
        _zz_stage0_mask = 8'hff;
      end
    endcase
  end

  assign stage0_mask = (_zz_stage0_mask <<< io_cpu_execute_address[2 : 0]);
  assign _zz_stage0_dataColisions = io_cpu_execute_address[11 : 3];
  assign _zz_stage0_dataColisions_1 = dataWriteCmd_payload_mask[7 : 0];
  always @(*) begin
    stage0_dataColisions[0] = (((dataWriteCmd_valid && dataWriteCmd_payload_way[0]) && (dataWriteCmd_payload_address == _zz_stage0_dataColisions)) && ((stage0_mask & _zz_stage0_dataColisions_1) != 8'h0));
    stage0_dataColisions[1] = (((dataWriteCmd_valid && dataWriteCmd_payload_way[1]) && (dataWriteCmd_payload_address == _zz_stage0_dataColisions)) && ((stage0_mask & _zz_stage0_dataColisions_1) != 8'h0));
  end

  always @(*) begin
    stage0_wayInvalidate = 2'b00;
    if(when_DataCache_l1167) begin
      if(when_DataCache_l1169) begin
        stage0_wayInvalidate = invalidate_s2_wayHits;
      end
    end
  end

  assign when_DataCache_l776 = (! io_cpu_memory_isStuck);
  assign when_DataCache_l776_1 = (! io_cpu_memory_isStuck);
  assign io_cpu_memory_isWrite = stageA_request_wr;
  always @(*) begin
    stageA_consistancyCheck_hazard = 1'b0;
    if(when_DataCache_l793) begin
      stageA_consistancyCheck_hazard = 1'b1;
    end
    if(when_DataCache_l796) begin
      stageA_consistancyCheck_hazard = 1'b1;
    end
  end

  assign stageA_consistancyCheck_w = (sync_w2w_busy || sync_o2w_busy);
  assign when_DataCache_l776_2 = (! io_cpu_memory_isStuck);
  assign stageA_consistancyCheck_r = ((_zz_stageA_consistancyCheck_r || sync_w2r_busy) || sync_o2r_busy);
  assign stageA_consistancyCheck_o = sync_w2o_busy;
  assign stageA_consistancyCheck_i = sync_w2i_busy;
  assign stageA_consistancyCheck_s = (io_cpu_memory_mmuRsp_isIoAccess ? stageA_consistancyCheck_o : stageA_consistancyCheck_w);
  assign stageA_consistancyCheck_l = (io_cpu_memory_mmuRsp_isIoAccess ? stageA_consistancyCheck_i : stageA_consistancyCheck_r);
  assign when_DataCache_l793 = (stageA_request_isAmo ? (stageA_consistancyCheck_s || stageA_consistancyCheck_l) : (stageA_request_wr ? stageA_consistancyCheck_s : stageA_consistancyCheck_l));
  assign when_DataCache_l796 = (stageA_request_totalyConsistent && (sync_notTotalyConsistent || (io_cpu_writeBack_isValid && io_cpu_writeBack_isWrite)));
  assign stageA_wayHits = {((io_cpu_memory_mmuRsp_physicalAddress[31 : 12] == ways_1_tagsReadRsp_address) && ways_1_tagsReadRsp_valid),((io_cpu_memory_mmuRsp_physicalAddress[31 : 12] == ways_0_tagsReadRsp_address) && ways_0_tagsReadRsp_valid)};
  assign when_DataCache_l776_3 = (! io_cpu_memory_isStuck);
  assign when_DataCache_l776_4 = (! io_cpu_memory_isStuck);
  assign _zz_stageA_dataColisions_1 = io_cpu_memory_address[11 : 3];
  assign _zz_stageA_dataColisions_2 = dataWriteCmd_payload_mask[7 : 0];
  always @(*) begin
    _zz_stageA_dataColisions[0] = (((dataWriteCmd_valid && dataWriteCmd_payload_way[0]) && (dataWriteCmd_payload_address == _zz_stageA_dataColisions_1)) && ((stageA_mask & _zz_stageA_dataColisions_2) != 8'h0));
    _zz_stageA_dataColisions[1] = (((dataWriteCmd_valid && dataWriteCmd_payload_way[1]) && (dataWriteCmd_payload_address == _zz_stageA_dataColisions_1)) && ((stageA_mask & _zz_stageA_dataColisions_2) != 8'h0));
  end

  assign stageA_dataColisions = (stage0_dataColisions_regNextWhen | _zz_stageA_dataColisions);
  assign when_DataCache_l827 = (! io_cpu_writeBack_isStuck);
  always @(*) begin
    stageB_mmuRspFreeze = 1'b0;
    if(when_DataCache_l1132) begin
      stageB_mmuRspFreeze = 1'b1;
    end
  end

  assign when_DataCache_l829 = ((! io_cpu_writeBack_isStuck) && (! stageB_mmuRspFreeze));
  assign when_DataCache_l826 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l826_1 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l826_2 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l826_3 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l825 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l825_1 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l825_2 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l825_3 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l825_4 = (! io_cpu_writeBack_isStuck);
  assign stageB_waysHits = (stageB_waysHitsBeforeInvalidate & (~ stageB_wayInvalidate));
  assign stageB_waysHit = (|stageB_waysHits);
  assign stageB_dataMux = (stageB_waysHits[0] ? stageB_dataReadRsp_0 : stageB_dataReadRsp_1);
  assign when_DataCache_l825_5 = (! io_cpu_writeBack_isStuck);
  always @(*) begin
    stageB_loaderValid = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_request_isAmo) begin
        if(!when_DataCache_l996) begin
          if(!when_DataCache_l1009) begin
            if(io_mem_cmd_ready) begin
              stageB_loaderValid = 1'b1;
            end
          end
        end
      end
    end
    if(io_cpu_writeBack_isValid) begin
      if(when_DataCache_l1072) begin
        stageB_loaderValid = 1'b0;
      end
    end
  end

  assign stageB_ioMemRspMuxed = io_mem_rsp_payload_data[63 : 0];
  always @(*) begin
    io_cpu_writeBack_haltIt = 1'b1;
    if(io_cpu_writeBack_isValid) begin
      if(stageB_request_isAmo) begin
        case(stageB_amo_external_state)
          DataCacheExternalAmoStates_LR_CMD : begin
          end
          DataCacheExternalAmoStates_LR_RSP : begin
          end
          DataCacheExternalAmoStates_SC_CMD : begin
          end
          default : begin
            if(io_mem_rsp_valid) begin
              if(io_mem_rsp_payload_exclusive) begin
                io_cpu_writeBack_haltIt = 1'b0;
              end
            end
          end
        endcase
      end else begin
        if(when_DataCache_l996) begin
          if(when_DataCache_l1000) begin
            io_cpu_writeBack_haltIt = 1'b0;
          end
        end else begin
          if(when_DataCache_l1009) begin
            if(when_DataCache_l1014) begin
              io_cpu_writeBack_haltIt = 1'b0;
            end
          end
        end
      end
    end
    if(io_cpu_writeBack_isValid) begin
      if(when_DataCache_l1072) begin
        io_cpu_writeBack_haltIt = 1'b0;
      end
    end
  end

  always @(*) begin
    stageB_flusher_hold = 1'b0;
    if(when_DataCache_l1167) begin
      if(invalidate_s2_wayHit) begin
        stageB_flusher_hold = 1'b1;
      end
    end
  end

  assign when_DataCache_l855 = (! stageB_flusher_counter[6]);
  assign when_DataCache_l861 = (! stageB_flusher_hold);
  assign when_DataCache_l863 = (io_cpu_flush_valid && io_cpu_flush_payload_singleLine);
  assign io_cpu_flush_ready = (stageB_flusher_waitDone && stageB_flusher_counter[6]);
  assign when_DataCache_l877 = (io_cpu_flush_valid && io_cpu_flush_payload_singleLine);
  assign stageB_isAmoCached = 1'b0;
  always @(*) begin
    stageB_requestDataBypass = io_cpu_writeBack_storeData;
    if(stageB_request_isAmo) begin
      stageB_requestDataBypass[31 : 0] = stageB_amo_resultReg;
      stageB_requestDataBypass[63 : 32] = stageB_amo_resultReg;
    end
  end

  assign stageB_amo_compare = stageB_request_amoCtrl_alu[2];
  assign stageB_amo_unsigned = (stageB_request_amoCtrl_alu[2 : 1] == 2'b11);
  assign stageB_amo_addSub = _zz_stageB_amo_addSub;
  assign stageB_amo_less = ((io_cpu_writeBack_storeData[31] == _zz_stageB_amo_less[31]) ? stageB_amo_addSub[31] : (stageB_amo_unsigned ? _zz_stageB_amo_less_2[31] : io_cpu_writeBack_storeData[31]));
  assign stageB_amo_selectRf = (stageB_request_amoCtrl_swap ? 1'b1 : (stageB_request_amoCtrl_alu[0] ^ stageB_amo_less));
  assign switch_Misc_l241 = (stageB_request_amoCtrl_alu | {stageB_request_amoCtrl_swap,2'b00});
  always @(*) begin
    case(switch_Misc_l241)
      3'b000 : begin
        stageB_amo_result = stageB_amo_addSub;
      end
      3'b001 : begin
        stageB_amo_result = (io_cpu_writeBack_storeData[31 : 0] ^ _zz_stageB_amo_result);
      end
      3'b010 : begin
        stageB_amo_result = (io_cpu_writeBack_storeData[31 : 0] | _zz_stageB_amo_result_2);
      end
      3'b011 : begin
        stageB_amo_result = (io_cpu_writeBack_storeData[31 : 0] & _zz_stageB_amo_result_4);
      end
      default : begin
        stageB_amo_result = (stageB_amo_selectRf ? io_cpu_writeBack_storeData[31 : 0] : _zz_stageB_amo_result_6);
      end
    endcase
  end

  always @(*) begin
    stageB_cpuWriteToCache = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(stageB_request_isAmo) begin
        case(stageB_amo_external_state)
          DataCacheExternalAmoStates_LR_CMD : begin
          end
          DataCacheExternalAmoStates_LR_RSP : begin
          end
          DataCacheExternalAmoStates_SC_CMD : begin
          end
          default : begin
            if(io_mem_rsp_valid) begin
              if(io_mem_rsp_payload_exclusive) begin
                stageB_cpuWriteToCache = 1'b1;
              end
            end
          end
        endcase
      end else begin
        if(!when_DataCache_l996) begin
          if(when_DataCache_l1009) begin
            stageB_cpuWriteToCache = 1'b1;
          end
        end
      end
    end
    if(when_DataCache_l1059) begin
      if(when_DataCache_l1061) begin
        stageB_cpuWriteToCache = 1'b1;
      end
    end
  end

  assign when_DataCache_l931 = (stageB_request_wr && stageB_waysHit);
  assign stageB_badPermissions = (((! stageB_mmuRsp_allowWrite) && stageB_request_wr) || ((! stageB_mmuRsp_allowRead) && ((! stageB_request_wr) || stageB_request_isAmo)));
  assign stageB_loadStoreFault = (io_cpu_writeBack_isValid && (stageB_mmuRsp_exception || stageB_badPermissions));
  always @(*) begin
    io_cpu_redo = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_request_isAmo) begin
        if(!when_DataCache_l996) begin
          if(when_DataCache_l1009) begin
            if(when_DataCache_l1025) begin
              io_cpu_redo = 1'b1;
            end
          end
        end
      end
    end
    if(io_cpu_writeBack_isValid) begin
      if(when_DataCache_l1081) begin
        io_cpu_redo = 1'b1;
      end
    end
    if(when_DataCache_l1129) begin
      io_cpu_redo = 1'b1;
    end
  end

  always @(*) begin
    io_cpu_writeBack_accessError = 1'b0;
    if(stageB_bypassCache) begin
      io_cpu_writeBack_accessError = ((((! stageB_request_wr) && pending_last) && io_mem_rsp_valid) && io_mem_rsp_payload_error);
    end else begin
      io_cpu_writeBack_accessError = (((stageB_waysHits & {stageB_tagsReadRsp_1_error,stageB_tagsReadRsp_0_error}) != 2'b00) || (stageB_loadStoreFault && (! stageB_mmuRsp_isPaging)));
    end
  end

  assign io_cpu_writeBack_mmuException = (stageB_loadStoreFault && stageB_mmuRsp_isPaging);
  assign io_cpu_writeBack_unalignedAccess = (io_cpu_writeBack_isValid && stageB_unaligned);
  assign io_cpu_writeBack_isWrite = stageB_request_wr;
  always @(*) begin
    io_mem_cmd_valid = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(stageB_request_isAmo) begin
        case(stageB_amo_external_state)
          DataCacheExternalAmoStates_LR_CMD : begin
            io_mem_cmd_valid = 1'b1;
          end
          DataCacheExternalAmoStates_LR_RSP : begin
          end
          DataCacheExternalAmoStates_SC_CMD : begin
            io_mem_cmd_valid = 1'b1;
          end
          default : begin
          end
        endcase
      end else begin
        if(when_DataCache_l996) begin
          io_mem_cmd_valid = (! memCmdSent);
        end else begin
          if(when_DataCache_l1009) begin
            if(stageB_request_wr) begin
              io_mem_cmd_valid = 1'b1;
            end
            if(when_DataCache_l1025) begin
              io_mem_cmd_valid = 1'b0;
            end
          end else begin
            if(when_DataCache_l1037) begin
              io_mem_cmd_valid = 1'b1;
            end
          end
        end
      end
    end
    if(io_cpu_writeBack_isValid) begin
      if(when_DataCache_l1072) begin
        io_mem_cmd_valid = 1'b0;
      end
    end
  end

  always @(*) begin
    io_mem_cmd_payload_address = stageB_mmuRsp_physicalAddress;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_request_isAmo) begin
        if(!when_DataCache_l996) begin
          if(!when_DataCache_l1009) begin
            io_mem_cmd_payload_address[5 : 0] = 6'h0;
          end
        end
      end
    end
  end

  assign io_mem_cmd_payload_last = 1'b1;
  always @(*) begin
    io_mem_cmd_payload_wr = stageB_request_wr;
    if(io_cpu_writeBack_isValid) begin
      if(stageB_request_isAmo) begin
        case(stageB_amo_external_state)
          DataCacheExternalAmoStates_LR_CMD : begin
            io_mem_cmd_payload_wr = 1'b0;
          end
          DataCacheExternalAmoStates_LR_RSP : begin
          end
          DataCacheExternalAmoStates_SC_CMD : begin
          end
          default : begin
          end
        endcase
      end else begin
        if(!when_DataCache_l996) begin
          if(!when_DataCache_l1009) begin
            io_mem_cmd_payload_wr = 1'b0;
          end
        end
      end
    end
  end

  assign io_mem_cmd_payload_mask = stageB_mask;
  assign io_mem_cmd_payload_data = stageB_requestDataBypass;
  assign io_mem_cmd_payload_uncached = stageB_mmuRsp_isIoAccess;
  always @(*) begin
    io_mem_cmd_payload_size = {1'd0, stageB_request_size};
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_request_isAmo) begin
        if(!when_DataCache_l996) begin
          if(!when_DataCache_l1009) begin
            io_mem_cmd_payload_size = 3'b110;
          end
        end
      end
    end
  end

  assign io_mem_cmd_payload_exclusive = (stageB_request_isLrsc || stageB_request_isAmo);
  assign stageB_bypassCache = ((stageB_mmuRsp_isIoAccess || stageB_request_isLrsc) || stageB_request_isAmo);
  always @(*) begin
    io_cpu_writeBack_keepMemRspData = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(stageB_request_isAmo) begin
        case(stageB_amo_external_state)
          DataCacheExternalAmoStates_LR_CMD : begin
          end
          DataCacheExternalAmoStates_LR_RSP : begin
          end
          DataCacheExternalAmoStates_SC_CMD : begin
          end
          default : begin
            io_cpu_writeBack_keepMemRspData = 1'b1;
          end
        endcase
      end
    end
  end

  assign when_DataCache_l974 = (io_mem_rsp_valid && pending_last);
  always @(*) begin
    _zz_when_DataCache_l1000 = (! stageB_request_wr);
    if(stageB_request_isLrsc) begin
      _zz_when_DataCache_l1000 = 1'b1;
    end
  end

  assign when_DataCache_l1000 = (_zz_when_DataCache_l1000 ? (io_mem_rsp_valid && rspSync) : io_mem_cmd_ready);
  assign when_DataCache_l1009 = (stageB_waysHit || (stageB_request_wr && (! stageB_isAmoCached)));
  assign when_DataCache_l1014 = ((! stageB_request_wr) || io_mem_cmd_ready);
  assign when_DataCache_l1025 = (((! stageB_request_wr) || stageB_isAmoCached) && ((stageB_dataColisions & stageB_waysHits) != 2'b00));
  assign when_DataCache_l1037 = (! memCmdSent);
  assign when_DataCache_l996 = (stageB_mmuRsp_isIoAccess || stageB_request_isLrsc);
  always @(*) begin
    if(stageB_bypassCache) begin
      io_cpu_writeBack_data = stageB_ioMemRspMuxed;
    end else begin
      io_cpu_writeBack_data = stageB_dataMux;
    end
  end

  assign io_cpu_writeBack_exclusiveOk = io_mem_rsp_payload_exclusive;
  assign when_DataCache_l1059 = (stageB_request_isLrsc && stageB_request_wr);
  assign when_DataCache_l1061 = ((((io_cpu_writeBack_isValid && io_mem_rsp_valid) && rspSync) && io_mem_rsp_payload_exclusive) && stageB_waysHit);
  assign when_DataCache_l1072 = ((((stageB_consistancyHazard || stageB_mmuRsp_refilling) || io_cpu_writeBack_accessError) || io_cpu_writeBack_mmuException) || io_cpu_writeBack_unalignedAccess);
  assign when_DataCache_l1081 = (stageB_mmuRsp_refilling || stageB_consistancyHazard);
  always @(*) begin
    loader_counter_willIncrement = 1'b0;
    if(when_DataCache_l1097) begin
      loader_counter_willIncrement = 1'b1;
    end
  end

  assign loader_counter_willClear = 1'b0;
  assign loader_counter_willOverflowIfInc = (loader_counter_value == 3'b111);
  assign loader_counter_willOverflow = (loader_counter_willOverflowIfInc && loader_counter_willIncrement);
  always @(*) begin
    loader_counter_valueNext = (loader_counter_value + _zz_loader_counter_valueNext);
    if(loader_counter_willClear) begin
      loader_counter_valueNext = 3'b000;
    end
  end

  always @(*) begin
    loader_kill = 1'b0;
    if(when_DataCache_l1143) begin
      loader_kill = 1'b1;
    end
  end

  assign when_DataCache_l1097 = ((loader_valid && io_mem_rsp_valid) && rspLast);
  always @(*) begin
    loader_done = loader_counter_willOverflow;
    if(when_DataCache_l1108) begin
      loader_done = 1'b1;
    end
    if(when_DataCache_l1167) begin
      if(invalidate_s2_wayHit) begin
        loader_done = 1'b0;
      end
    end
  end

  assign when_DataCache_l1108 = (loader_valid && (pending_counter == 7'h0));
  assign when_DataCache_l1125 = (! loader_valid);
  assign when_DataCache_l1129 = (loader_valid && (! loader_valid_regNext));
  assign io_cpu_execute_refilling = loader_valid;
  assign when_DataCache_l1132 = (stageB_loaderValid || loader_valid);
  assign io_mem_inv_fire = (io_mem_inv_valid && io_mem_inv_ready);
  assign tagsInvReadCmd_valid = io_mem_inv_fire;
  assign tagsInvReadCmd_payload = io_mem_inv_payload_fragment_address[11 : 6];
  assign invalidate_s0_loaderTagHit = (io_mem_inv_payload_fragment_address[31 : 12] == stageB_mmuRsp_physicalAddress[31 : 12]);
  assign invalidate_s0_loaderLineHit = (io_mem_inv_payload_fragment_address[11 : 6] == stageB_mmuRsp_physicalAddress[11 : 6]);
  assign when_DataCache_l1143 = ((((io_mem_inv_valid && io_mem_inv_payload_fragment_enable) && loader_valid) && invalidate_s0_loaderLineHit) && invalidate_s0_loaderTagHit);
  always @(*) begin
    io_mem_inv_ready = invalidate_s1_input_ready;
    if(when_Stream_l375) begin
      io_mem_inv_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! invalidate_s1_input_valid);
  assign invalidate_s1_input_valid = io_mem_inv_rValid;
  assign invalidate_s1_input_payload_last = io_mem_inv_rData_last;
  assign invalidate_s1_input_payload_fragment_enable = io_mem_inv_rData_fragment_enable;
  assign invalidate_s1_input_payload_fragment_address = io_mem_inv_rData_fragment_address;
  assign invalidate_s1_wayHits = ({((invalidate_s1_input_payload_fragment_address[31 : 12] == ways_1_tagsInvReadRsp_address) && ways_1_tagsInvReadRsp_valid),((invalidate_s1_input_payload_fragment_address[31 : 12] == ways_0_tagsInvReadRsp_address) && ways_0_tagsInvReadRsp_valid)} & (~ invalidate_s1_invalidations));
  assign when_DataCache_l1158 = ((invalidate_s1_loaderValid && invalidate_s1_loaderLineHit) && (! invalidate_s1_loaderTagHit));
  always @(*) begin
    invalidate_s1_input_ready = invalidate_s2_input_ready;
    if(when_Stream_l375_1) begin
      invalidate_s1_input_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! invalidate_s2_input_valid);
  assign invalidate_s2_input_valid = invalidate_s1_input_rValid;
  assign invalidate_s2_input_payload_last = invalidate_s1_input_rData_last;
  assign invalidate_s2_input_payload_fragment_enable = invalidate_s1_input_rData_fragment_enable;
  assign invalidate_s2_input_payload_fragment_address = invalidate_s1_input_rData_fragment_address;
  assign invalidate_s2_wayHit = (|invalidate_s2_wayHits);
  assign when_DataCache_l1167 = (invalidate_s2_input_valid && invalidate_s2_input_payload_fragment_enable);
  assign when_DataCache_l1169 = (invalidate_s2_input_payload_fragment_address[11 : 6] == io_cpu_execute_address[11 : 6]);
  assign io_mem_ack_valid = invalidate_s2_input_valid;
  assign invalidate_s2_input_ready = io_mem_ack_ready;
  assign io_mem_ack_payload_fragment_hit = invalidate_s2_wayHit;
  assign io_mem_ack_payload_last = invalidate_s2_input_payload_last;
  assign invalidate_s1_invalidations = _zz_invalidate_s1_invalidations;
  always @(posedge io_systemClk) begin
    tagsWriteLastCmd_valid <= tagsWriteCmd_valid;
    tagsWriteLastCmd_payload_way <= tagsWriteCmd_payload_way;
    tagsWriteLastCmd_payload_address <= tagsWriteCmd_payload_address;
    tagsWriteLastCmd_payload_data_valid <= tagsWriteCmd_payload_data_valid;
    tagsWriteLastCmd_payload_data_error <= tagsWriteCmd_payload_data_error;
    tagsWriteLastCmd_payload_data_address <= tagsWriteCmd_payload_data_address;
    pending_done <= (pending_counterNext == 7'h0);
    pending_full <= pending_counter[6];
    pending_last <= (pending_counterNext == 7'h01);
    sync_syncContext_full <= (7'h3f <= _zz_sync_syncContext_full);
    if(when_DataCache_l776) begin
      stageA_request_wr <= io_cpu_execute_args_wr;
      stageA_request_size <= io_cpu_execute_args_size;
      stageA_request_isLrsc <= io_cpu_execute_args_isLrsc;
      stageA_request_isAmo <= io_cpu_execute_args_isAmo;
      stageA_request_amoCtrl_swap <= io_cpu_execute_args_amoCtrl_swap;
      stageA_request_amoCtrl_alu <= io_cpu_execute_args_amoCtrl_alu;
      stageA_request_totalyConsistent <= io_cpu_execute_args_totalyConsistent;
    end
    if(when_DataCache_l776_1) begin
      stageA_mask <= stage0_mask;
    end
    if(when_DataCache_l776_2) begin
      _zz_stageA_consistancyCheck_r <= (sync_w2r_busy || sync_o2r_busy);
    end
    if(when_DataCache_l776_3) begin
      stageA_wayInvalidate <= stage0_wayInvalidate;
    end
    if(when_DataCache_l776_4) begin
      stage0_dataColisions_regNextWhen <= stage0_dataColisions;
    end
    if(when_DataCache_l827) begin
      stageB_request_wr <= stageA_request_wr;
      stageB_request_size <= stageA_request_size;
      stageB_request_isLrsc <= stageA_request_isLrsc;
      stageB_request_isAmo <= stageA_request_isAmo;
      stageB_request_amoCtrl_swap <= stageA_request_amoCtrl_swap;
      stageB_request_amoCtrl_alu <= stageA_request_amoCtrl_alu;
      stageB_request_totalyConsistent <= stageA_request_totalyConsistent;
    end
    if(when_DataCache_l829) begin
      stageB_mmuRsp_physicalAddress <= io_cpu_memory_mmuRsp_physicalAddress;
      stageB_mmuRsp_isIoAccess <= io_cpu_memory_mmuRsp_isIoAccess;
      stageB_mmuRsp_isPaging <= io_cpu_memory_mmuRsp_isPaging;
      stageB_mmuRsp_allowRead <= io_cpu_memory_mmuRsp_allowRead;
      stageB_mmuRsp_allowWrite <= io_cpu_memory_mmuRsp_allowWrite;
      stageB_mmuRsp_allowExecute <= io_cpu_memory_mmuRsp_allowExecute;
      stageB_mmuRsp_exception <= io_cpu_memory_mmuRsp_exception;
      stageB_mmuRsp_refilling <= io_cpu_memory_mmuRsp_refilling;
      stageB_mmuRsp_bypassTranslation <= io_cpu_memory_mmuRsp_bypassTranslation;
    end
    if(when_DataCache_l826) begin
      stageB_tagsReadRsp_0_valid <= ways_0_tagsReadRsp_valid;
      stageB_tagsReadRsp_0_error <= ways_0_tagsReadRsp_error;
      stageB_tagsReadRsp_0_address <= ways_0_tagsReadRsp_address;
    end
    if(when_DataCache_l826_1) begin
      stageB_tagsReadRsp_1_valid <= ways_1_tagsReadRsp_valid;
      stageB_tagsReadRsp_1_error <= ways_1_tagsReadRsp_error;
      stageB_tagsReadRsp_1_address <= ways_1_tagsReadRsp_address;
    end
    if(when_DataCache_l826_2) begin
      stageB_dataReadRsp_0 <= ways_0_dataReadRsp;
    end
    if(when_DataCache_l826_3) begin
      stageB_dataReadRsp_1 <= ways_1_dataReadRsp;
    end
    if(when_DataCache_l825) begin
      stageB_wayInvalidate <= stageA_wayInvalidate;
    end
    if(when_DataCache_l825_1) begin
      stageB_consistancyHazard <= stageA_consistancyCheck_hazard;
    end
    if(when_DataCache_l825_2) begin
      stageB_dataColisions <= stageA_dataColisions;
    end
    if(when_DataCache_l825_3) begin
      stageB_unaligned <= (|{((stageA_request_size == 2'b11) && (io_cpu_memory_address[2 : 0] != 3'b000)),{((stageA_request_size == 2'b10) && (io_cpu_memory_address[1 : 0] != 2'b00)),((stageA_request_size == 2'b01) && (io_cpu_memory_address[0 : 0] != 1'b0))}});
    end
    if(when_DataCache_l825_4) begin
      stageB_waysHitsBeforeInvalidate <= stageA_wayHits;
    end
    if(when_DataCache_l825_5) begin
      stageB_mask <= stageA_mask;
    end
    if(io_cpu_writeBack_isValid) begin
      if(stageB_request_isAmo) begin
        case(stageB_amo_external_state)
          DataCacheExternalAmoStates_LR_CMD : begin
          end
          DataCacheExternalAmoStates_LR_RSP : begin
            if(when_DataCache_l974) begin
              stageB_amo_resultReg <= stageB_amo_result;
            end
          end
          DataCacheExternalAmoStates_SC_CMD : begin
          end
          default : begin
          end
        endcase
      end
    end
    loader_valid_regNext <= loader_valid;
    if(io_mem_inv_ready) begin
      io_mem_inv_rData_last <= io_mem_inv_payload_last;
      io_mem_inv_rData_fragment_enable <= io_mem_inv_payload_fragment_enable;
      io_mem_inv_rData_fragment_address <= io_mem_inv_payload_fragment_address;
    end
    if(io_mem_inv_ready) begin
      invalidate_s1_loaderValid <= loader_valid;
    end
    if(io_mem_inv_ready) begin
      invalidate_s1_loaderWay <= loader_waysAllocator;
    end
    if(io_mem_inv_ready) begin
      invalidate_s1_loaderTagHit <= invalidate_s0_loaderTagHit;
    end
    if(io_mem_inv_ready) begin
      invalidate_s1_loaderLineHit <= invalidate_s0_loaderLineHit;
    end
    if(invalidate_s1_input_ready) begin
      invalidate_s1_input_rData_last <= invalidate_s1_input_payload_last;
      invalidate_s1_input_rData_fragment_enable <= invalidate_s1_input_payload_fragment_enable;
      invalidate_s1_input_rData_fragment_address <= invalidate_s1_input_payload_fragment_address;
    end
    if(invalidate_s1_input_ready) begin
      invalidate_s2_wayHits <= invalidate_s1_wayHits_1;
    end
    if(io_mem_inv_ready) begin
      _zz_invalidate_s1_invalidations <= (((invalidate_s2_input_valid && invalidate_s2_input_payload_fragment_enable) && (invalidate_s2_input_payload_fragment_address[11 : 6] == io_mem_inv_payload_fragment_address[11 : 6])) ? invalidate_s2_wayHits : 2'b00);
    end
  end

  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      memCmdSent <= 1'b0;
      pending_counter <= 7'h0;
      sync_syncContext_wPtr <= 7'h0;
      sync_syncContext_rPtr <= 7'h0;
      sync_writeCached_pendingSync <= 7'h0;
      sync_writeUncached_pendingSync <= 7'h0;
      sync_w2w_counter <= 7'h0;
      sync_w2r_counter <= 7'h0;
      sync_w2i_counter <= 7'h0;
      sync_w2o_counter <= 7'h0;
      sync_o2w_counter <= 7'h0;
      sync_o2r_counter <= 7'h0;
      stageB_flusher_waitDone <= 1'b0;
      stageB_flusher_counter <= 7'h0;
      stageB_flusher_start <= 1'b1;
      stageB_amo_external_state <= DataCacheExternalAmoStates_LR_CMD;
      loader_valid <= 1'b0;
      loader_counter_value <= 3'b000;
      loader_waysAllocator <= 2'b01;
      loader_error <= 1'b0;
      loader_killReg <= 1'b0;
      io_mem_inv_rValid <= 1'b0;
      invalidate_s1_input_rValid <= 1'b0;
    end else begin
      if(io_mem_cmd_fire) begin
        memCmdSent <= 1'b1;
      end
      if(when_DataCache_l689) begin
        memCmdSent <= 1'b0;
      end
      pending_counter <= pending_counterNext;
      if(when_DataCache_l713) begin
        sync_syncContext_wPtr <= (sync_syncContext_wPtr + 7'h01);
      end
      if(io_mem_sync_fire) begin
        sync_syncContext_rPtr <= (sync_syncContext_rPtr + _zz_sync_syncContext_rPtr);
      end
      sync_writeCached_pendingSync <= sync_writeCached_pendingSyncNext;
      sync_writeUncached_pendingSync <= sync_writeUncached_pendingSyncNext;
      sync_w2w_counter <= (sync_w2w_counter - _zz_sync_w2w_counter);
      if(when_DataCache_l740) begin
        sync_w2w_counter <= sync_writeCached_pendingSyncNext;
      end
      sync_w2r_counter <= (sync_w2r_counter - _zz_sync_w2r_counter);
      if(when_DataCache_l740_1) begin
        sync_w2r_counter <= sync_writeCached_pendingSyncNext;
      end
      sync_w2i_counter <= (sync_w2i_counter - _zz_sync_w2i_counter);
      if(when_DataCache_l740_2) begin
        sync_w2i_counter <= sync_writeCached_pendingSyncNext;
      end
      sync_w2o_counter <= (sync_w2o_counter - _zz_sync_w2o_counter);
      if(when_DataCache_l740_3) begin
        sync_w2o_counter <= sync_writeCached_pendingSyncNext;
      end
      sync_o2w_counter <= (sync_o2w_counter - _zz_sync_o2w_counter);
      if(when_DataCache_l740_4) begin
        sync_o2w_counter <= sync_writeUncached_pendingSyncNext;
      end
      sync_o2r_counter <= (sync_o2r_counter - _zz_sync_o2r_counter);
      if(when_DataCache_l740_5) begin
        sync_o2r_counter <= sync_writeUncached_pendingSyncNext;
      end
      if(io_cpu_flush_ready) begin
        stageB_flusher_waitDone <= 1'b0;
      end
      if(when_DataCache_l855) begin
        if(when_DataCache_l861) begin
          stageB_flusher_counter <= (stageB_flusher_counter + 7'h01);
          if(when_DataCache_l863) begin
            stageB_flusher_counter[6] <= 1'b1;
          end
        end
      end
      stageB_flusher_start <= (((((((! stageB_flusher_waitDone) && (! stageB_flusher_start)) && io_cpu_flush_valid) && (! io_cpu_execute_isValid)) && (! io_cpu_memory_isValid)) && (! io_cpu_writeBack_isValid)) && (! io_cpu_redo));
      if(stageB_flusher_start) begin
        stageB_flusher_waitDone <= 1'b1;
        stageB_flusher_counter <= 7'h0;
        if(when_DataCache_l877) begin
          stageB_flusher_counter <= {1'b0,io_cpu_flush_payload_lineId};
        end
      end
      if(io_cpu_writeBack_isValid) begin
        if(stageB_request_isAmo) begin
          case(stageB_amo_external_state)
            DataCacheExternalAmoStates_LR_CMD : begin
              if(io_mem_cmd_ready) begin
                stageB_amo_external_state <= DataCacheExternalAmoStates_LR_RSP;
              end
            end
            DataCacheExternalAmoStates_LR_RSP : begin
              if(when_DataCache_l974) begin
                stageB_amo_external_state <= DataCacheExternalAmoStates_SC_CMD;
              end
            end
            DataCacheExternalAmoStates_SC_CMD : begin
              if(io_mem_cmd_ready) begin
                stageB_amo_external_state <= DataCacheExternalAmoStates_SC_RSP;
              end
            end
            default : begin
              if(io_mem_rsp_valid) begin
                stageB_amo_external_state <= DataCacheExternalAmoStates_LR_CMD;
              end
            end
          endcase
        end
      end
      if(io_cpu_writeBack_isValid) begin
        if(when_DataCache_l1072) begin
          stageB_amo_external_state <= DataCacheExternalAmoStates_LR_CMD;
        end
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((io_cpu_writeBack_isValid && (! io_cpu_writeBack_haltIt)) && io_cpu_writeBack_isStuck))); // DataCache.scala:L1084
        `else
          if(!(! ((io_cpu_writeBack_isValid && (! io_cpu_writeBack_haltIt)) && io_cpu_writeBack_isStuck))) begin
            $display("ERROR writeBack stuck by another plugin is not allowed"); // DataCache.scala:L1084
          end
        `endif
      `endif
      if(stageB_loaderValid) begin
        loader_valid <= 1'b1;
      end
      loader_counter_value <= loader_counter_valueNext;
      if(loader_kill) begin
        loader_killReg <= 1'b1;
      end
      if(when_DataCache_l1097) begin
        loader_error <= (loader_error || io_mem_rsp_payload_error);
      end
      if(loader_done) begin
        loader_valid <= 1'b0;
        loader_error <= 1'b0;
        loader_killReg <= 1'b0;
      end
      if(when_DataCache_l1125) begin
        loader_waysAllocator <= _zz_loader_waysAllocator[1:0];
      end
      if(io_mem_inv_ready) begin
        io_mem_inv_rValid <= io_mem_inv_valid;
      end
      if(invalidate_s1_input_ready) begin
        invalidate_s1_input_rValid <= invalidate_s1_input_valid;
      end
    end
  end


endmodule

module InstructionCache (
  input  wire          io_flush,
  input  wire          io_cpu_prefetch_isValid,
  output reg           io_cpu_prefetch_haltIt,
  input  wire [31:0]   io_cpu_prefetch_pc,
  input  wire          io_cpu_fetch_isValid,
  input  wire          io_cpu_fetch_isStuck,
  input  wire          io_cpu_fetch_isRemoved,
  input  wire [31:0]   io_cpu_fetch_pc,
  output wire [31:0]   io_cpu_fetch_data,
  input  wire [31:0]   io_cpu_fetch_mmuRsp_physicalAddress,
  input  wire          io_cpu_fetch_mmuRsp_isIoAccess,
  input  wire          io_cpu_fetch_mmuRsp_isPaging,
  input  wire          io_cpu_fetch_mmuRsp_allowRead,
  input  wire          io_cpu_fetch_mmuRsp_allowWrite,
  input  wire          io_cpu_fetch_mmuRsp_allowExecute,
  input  wire          io_cpu_fetch_mmuRsp_exception,
  input  wire          io_cpu_fetch_mmuRsp_refilling,
  input  wire          io_cpu_fetch_mmuRsp_bypassTranslation,
  output wire [31:0]   io_cpu_fetch_physicalAddress,
  input  wire          io_cpu_decode_isValid,
  input  wire          io_cpu_decode_isStuck,
  input  wire [31:0]   io_cpu_decode_pc,
  output wire [31:0]   io_cpu_decode_physicalAddress,
  output wire [31:0]   io_cpu_decode_data,
  output wire          io_cpu_decode_cacheMiss,
  output wire          io_cpu_decode_error,
  output wire          io_cpu_decode_mmuRefilling,
  output wire          io_cpu_decode_mmuException,
  input  wire          io_cpu_decode_isUser,
  input  wire          io_cpu_fill_valid,
  input  wire [31:0]   io_cpu_fill_payload,
  output wire          io_mem_cmd_valid,
  input  wire          io_mem_cmd_ready,
  output wire [31:0]   io_mem_cmd_payload_address,
  output wire [2:0]    io_mem_cmd_payload_size,
  input  wire          io_mem_rsp_valid,
  input  wire [63:0]   io_mem_rsp_payload_data,
  input  wire          io_mem_rsp_payload_error,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  reg        [31:0]   banks_0_spinal_port1;
  reg        [31:0]   banks_1_spinal_port1;
  reg        [21:0]   ways_0_tags_spinal_port1;
  reg        [21:0]   ways_1_tags_spinal_port1;
  wire       [21:0]   _zz_ways_0_tags_port;
  wire       [21:0]   _zz_ways_1_tags_port;
  wire       [0:0]    _zz__zz_lineLoader_write_data_0_payload_address;
  reg        [31:0]   _zz_lineLoader_write_data_0_payload_data;
  wire       [0:0]    _zz__zz_lineLoader_write_data_1_payload_address;
  reg        [31:0]   _zz_lineLoader_write_data_1_payload_data;
  wire       [0:0]    _zz_fetchStage_hit_bankId;
  reg                 _zz_fetchStage_hit_error;
  reg        [31:0]   _zz_fetchStage_hit_data;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 _zz_3;
  reg                 _zz_4;
  reg                 lineLoader_fire;
  reg                 lineLoader_valid;
  (* keep , syn_keep *) reg        [31:0]   lineLoader_address /* synthesis syn_keep = 1 */ ;
  reg                 lineLoader_hadError;
  reg                 lineLoader_flushPending;
  reg        [6:0]    lineLoader_flushCounter;
  wire                when_InstructionCache_l338;
  reg                 _zz_when_InstructionCache_l342;
  wire                when_InstructionCache_l342;
  wire                when_InstructionCache_l351;
  reg                 lineLoader_cmdSent;
  wire                io_mem_cmd_fire;
  wire                when_Utils_l578;
  reg                 lineLoader_wayToAllocate_willIncrement;
  wire                lineLoader_wayToAllocate_willClear;
  reg        [0:0]    lineLoader_wayToAllocate_valueNext;
  reg        [0:0]    lineLoader_wayToAllocate_value;
  wire                lineLoader_wayToAllocate_willOverflowIfInc;
  wire                lineLoader_wayToAllocate_willOverflow;
  (* keep , syn_keep *) reg        [2:0]    lineLoader_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                lineLoader_write_tag_0_valid;
  wire       [5:0]    lineLoader_write_tag_0_payload_address;
  wire                lineLoader_write_tag_0_payload_data_valid;
  wire                lineLoader_write_tag_0_payload_data_error;
  wire       [19:0]   lineLoader_write_tag_0_payload_data_address;
  wire                lineLoader_write_tag_1_valid;
  wire       [5:0]    lineLoader_write_tag_1_payload_address;
  wire                lineLoader_write_tag_1_payload_data_valid;
  wire                lineLoader_write_tag_1_payload_data_error;
  wire       [19:0]   lineLoader_write_tag_1_payload_data_address;
  wire                lineLoader_write_data_0_valid;
  wire       [9:0]    lineLoader_write_data_0_payload_address;
  wire       [31:0]   lineLoader_write_data_0_payload_data;
  wire                lineLoader_write_data_1_valid;
  wire       [9:0]    lineLoader_write_data_1_payload_address;
  wire       [31:0]   lineLoader_write_data_1_payload_data;
  wire       [0:0]    _zz_lineLoader_write_data_0_payload_address;
  wire       [0:0]    _zz_lineLoader_write_data_1_payload_address;
  wire                when_InstructionCache_l401;
  wire       [9:0]    _zz_fetchStage_read_banksValue_0_dataMem;
  wire                _zz_fetchStage_read_banksValue_0_dataMem_1;
  wire       [31:0]   fetchStage_read_banksValue_0_dataMem;
  wire       [31:0]   fetchStage_read_banksValue_0_data;
  wire       [9:0]    _zz_fetchStage_read_banksValue_1_dataMem;
  wire                _zz_fetchStage_read_banksValue_1_dataMem_1;
  wire       [31:0]   fetchStage_read_banksValue_1_dataMem;
  wire       [31:0]   fetchStage_read_banksValue_1_data;
  wire       [5:0]    _zz_fetchStage_read_waysValues_0_tag_valid;
  wire                _zz_fetchStage_read_waysValues_0_tag_valid_1;
  wire                fetchStage_read_waysValues_0_tag_valid;
  wire                fetchStage_read_waysValues_0_tag_error;
  wire       [19:0]   fetchStage_read_waysValues_0_tag_address;
  wire       [21:0]   _zz_fetchStage_read_waysValues_0_tag_valid_2;
  wire       [5:0]    _zz_fetchStage_read_waysValues_1_tag_valid;
  wire                _zz_fetchStage_read_waysValues_1_tag_valid_1;
  wire                fetchStage_read_waysValues_1_tag_valid;
  wire                fetchStage_read_waysValues_1_tag_error;
  wire       [19:0]   fetchStage_read_waysValues_1_tag_address;
  wire       [21:0]   _zz_fetchStage_read_waysValues_1_tag_valid_2;
  wire                fetchStage_hit_hits_0;
  wire                fetchStage_hit_hits_1;
  wire                fetchStage_hit_valid;
  wire       [0:0]    fetchStage_hit_wayId;
  wire       [0:0]    fetchStage_hit_bankId;
  wire                fetchStage_hit_error;
  wire       [31:0]   fetchStage_hit_data;
  wire       [31:0]   fetchStage_hit_word;
  wire                when_InstructionCache_l435;
  reg        [31:0]   io_cpu_fetch_data_regNextWhen;
  wire                when_InstructionCache_l459;
  reg        [31:0]   decodeStage_mmuRsp_physicalAddress;
  reg                 decodeStage_mmuRsp_isIoAccess;
  reg                 decodeStage_mmuRsp_isPaging;
  reg                 decodeStage_mmuRsp_allowRead;
  reg                 decodeStage_mmuRsp_allowWrite;
  reg                 decodeStage_mmuRsp_allowExecute;
  reg                 decodeStage_mmuRsp_exception;
  reg                 decodeStage_mmuRsp_refilling;
  reg                 decodeStage_mmuRsp_bypassTranslation;
  wire                when_InstructionCache_l459_1;
  reg                 decodeStage_hit_valid;
  wire                when_InstructionCache_l459_2;
  reg                 decodeStage_hit_error;
  reg [31:0] banks_0 [0:1023];
  reg [31:0] banks_1 [0:1023];
  reg [21:0] ways_0_tags [0:63];
  reg [21:0] ways_1_tags [0:63];

  assign _zz__zz_lineLoader_write_data_0_payload_address = (1'b0 - lineLoader_wayToAllocate_value);
  assign _zz__zz_lineLoader_write_data_1_payload_address = (1'b1 - lineLoader_wayToAllocate_value);
  assign _zz_fetchStage_hit_bankId = (fetchStage_hit_wayId + io_cpu_fetch_mmuRsp_physicalAddress[2 : 2]);
  assign _zz_ways_0_tags_port = {lineLoader_write_tag_0_payload_data_address,{lineLoader_write_tag_0_payload_data_error,lineLoader_write_tag_0_payload_data_valid}};
  assign _zz_ways_1_tags_port = {lineLoader_write_tag_1_payload_data_address,{lineLoader_write_tag_1_payload_data_error,lineLoader_write_tag_1_payload_data_valid}};
  always @(posedge io_systemClk) begin
    if(_zz_2) begin
      banks_0[lineLoader_write_data_0_payload_address] <= lineLoader_write_data_0_payload_data;
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_fetchStage_read_banksValue_0_dataMem_1) begin
      banks_0_spinal_port1 <= banks_0[_zz_fetchStage_read_banksValue_0_dataMem];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_1) begin
      banks_1[lineLoader_write_data_1_payload_address] <= lineLoader_write_data_1_payload_data;
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_fetchStage_read_banksValue_1_dataMem_1) begin
      banks_1_spinal_port1 <= banks_1[_zz_fetchStage_read_banksValue_1_dataMem];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_4) begin
      ways_0_tags[lineLoader_write_tag_0_payload_address] <= _zz_ways_0_tags_port;
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_fetchStage_read_waysValues_0_tag_valid_1) begin
      ways_0_tags_spinal_port1 <= ways_0_tags[_zz_fetchStage_read_waysValues_0_tag_valid];
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_3) begin
      ways_1_tags[lineLoader_write_tag_1_payload_address] <= _zz_ways_1_tags_port;
    end
  end

  always @(posedge io_systemClk) begin
    if(_zz_fetchStage_read_waysValues_1_tag_valid_1) begin
      ways_1_tags_spinal_port1 <= ways_1_tags[_zz_fetchStage_read_waysValues_1_tag_valid];
    end
  end

  always @(*) begin
    case(_zz_lineLoader_write_data_0_payload_address)
      1'b0 : _zz_lineLoader_write_data_0_payload_data = io_mem_rsp_payload_data[31 : 0];
      default : _zz_lineLoader_write_data_0_payload_data = io_mem_rsp_payload_data[63 : 32];
    endcase
  end

  always @(*) begin
    case(_zz_lineLoader_write_data_1_payload_address)
      1'b0 : _zz_lineLoader_write_data_1_payload_data = io_mem_rsp_payload_data[31 : 0];
      default : _zz_lineLoader_write_data_1_payload_data = io_mem_rsp_payload_data[63 : 32];
    endcase
  end

  always @(*) begin
    case(fetchStage_hit_wayId)
      1'b0 : _zz_fetchStage_hit_error = fetchStage_read_waysValues_0_tag_error;
      default : _zz_fetchStage_hit_error = fetchStage_read_waysValues_1_tag_error;
    endcase
  end

  always @(*) begin
    case(fetchStage_hit_bankId)
      1'b0 : _zz_fetchStage_hit_data = fetchStage_read_banksValue_0_data;
      default : _zz_fetchStage_hit_data = fetchStage_read_banksValue_1_data;
    endcase
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(lineLoader_write_data_1_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(lineLoader_write_data_0_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    _zz_3 = 1'b0;
    if(lineLoader_write_tag_1_valid) begin
      _zz_3 = 1'b1;
    end
  end

  always @(*) begin
    _zz_4 = 1'b0;
    if(lineLoader_write_tag_0_valid) begin
      _zz_4 = 1'b1;
    end
  end

  always @(*) begin
    lineLoader_fire = 1'b0;
    if(io_mem_rsp_valid) begin
      if(when_InstructionCache_l401) begin
        lineLoader_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    io_cpu_prefetch_haltIt = (lineLoader_valid || lineLoader_flushPending);
    if(when_InstructionCache_l338) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(when_InstructionCache_l342) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(io_flush) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
  end

  assign when_InstructionCache_l338 = (! lineLoader_flushCounter[6]);
  assign when_InstructionCache_l342 = (! _zz_when_InstructionCache_l342);
  assign when_InstructionCache_l351 = (lineLoader_flushPending && (! (lineLoader_valid || io_cpu_fetch_isValid)));
  assign io_mem_cmd_fire = (io_mem_cmd_valid && io_mem_cmd_ready);
  assign io_mem_cmd_valid = (lineLoader_valid && (! lineLoader_cmdSent));
  assign io_mem_cmd_payload_address = {lineLoader_address[31 : 6],6'h0};
  assign io_mem_cmd_payload_size = 3'b110;
  assign when_Utils_l578 = (! lineLoader_valid);
  always @(*) begin
    lineLoader_wayToAllocate_willIncrement = 1'b0;
    if(when_Utils_l578) begin
      lineLoader_wayToAllocate_willIncrement = 1'b1;
    end
  end

  assign lineLoader_wayToAllocate_willClear = 1'b0;
  assign lineLoader_wayToAllocate_willOverflowIfInc = (lineLoader_wayToAllocate_value == 1'b1);
  assign lineLoader_wayToAllocate_willOverflow = (lineLoader_wayToAllocate_willOverflowIfInc && lineLoader_wayToAllocate_willIncrement);
  always @(*) begin
    lineLoader_wayToAllocate_valueNext = (lineLoader_wayToAllocate_value + lineLoader_wayToAllocate_willIncrement);
    if(lineLoader_wayToAllocate_willClear) begin
      lineLoader_wayToAllocate_valueNext = 1'b0;
    end
  end

  assign lineLoader_write_tag_0_valid = (((lineLoader_wayToAllocate_value == 1'b0) && lineLoader_fire) || (! lineLoader_flushCounter[6]));
  assign lineLoader_write_tag_0_payload_address = (lineLoader_flushCounter[6] ? lineLoader_address[11 : 6] : lineLoader_flushCounter[5 : 0]);
  assign lineLoader_write_tag_0_payload_data_valid = lineLoader_flushCounter[6];
  assign lineLoader_write_tag_0_payload_data_error = (lineLoader_hadError || io_mem_rsp_payload_error);
  assign lineLoader_write_tag_0_payload_data_address = lineLoader_address[31 : 12];
  assign lineLoader_write_tag_1_valid = (((lineLoader_wayToAllocate_value == 1'b1) && lineLoader_fire) || (! lineLoader_flushCounter[6]));
  assign lineLoader_write_tag_1_payload_address = (lineLoader_flushCounter[6] ? lineLoader_address[11 : 6] : lineLoader_flushCounter[5 : 0]);
  assign lineLoader_write_tag_1_payload_data_valid = lineLoader_flushCounter[6];
  assign lineLoader_write_tag_1_payload_data_error = (lineLoader_hadError || io_mem_rsp_payload_error);
  assign lineLoader_write_tag_1_payload_data_address = lineLoader_address[31 : 12];
  assign _zz_lineLoader_write_data_0_payload_address = _zz__zz_lineLoader_write_data_0_payload_address[0 : 0];
  assign lineLoader_write_data_0_valid = (io_mem_rsp_valid && 1'b1);
  assign lineLoader_write_data_0_payload_address = {{lineLoader_address[11 : 6],lineLoader_wordIndex},_zz_lineLoader_write_data_0_payload_address};
  assign lineLoader_write_data_0_payload_data = _zz_lineLoader_write_data_0_payload_data;
  assign _zz_lineLoader_write_data_1_payload_address = _zz__zz_lineLoader_write_data_1_payload_address[0 : 0];
  assign lineLoader_write_data_1_valid = (io_mem_rsp_valid && 1'b1);
  assign lineLoader_write_data_1_payload_address = {{lineLoader_address[11 : 6],lineLoader_wordIndex},_zz_lineLoader_write_data_1_payload_address};
  assign lineLoader_write_data_1_payload_data = _zz_lineLoader_write_data_1_payload_data;
  assign when_InstructionCache_l401 = (lineLoader_wordIndex == 3'b111);
  assign _zz_fetchStage_read_banksValue_0_dataMem = io_cpu_prefetch_pc[11 : 2];
  assign _zz_fetchStage_read_banksValue_0_dataMem_1 = (! io_cpu_fetch_isStuck);
  assign fetchStage_read_banksValue_0_dataMem = banks_0_spinal_port1;
  assign fetchStage_read_banksValue_0_data = fetchStage_read_banksValue_0_dataMem[31 : 0];
  assign _zz_fetchStage_read_banksValue_1_dataMem = io_cpu_prefetch_pc[11 : 2];
  assign _zz_fetchStage_read_banksValue_1_dataMem_1 = (! io_cpu_fetch_isStuck);
  assign fetchStage_read_banksValue_1_dataMem = banks_1_spinal_port1;
  assign fetchStage_read_banksValue_1_data = fetchStage_read_banksValue_1_dataMem[31 : 0];
  assign _zz_fetchStage_read_waysValues_0_tag_valid = io_cpu_prefetch_pc[11 : 6];
  assign _zz_fetchStage_read_waysValues_0_tag_valid_1 = (! io_cpu_fetch_isStuck);
  assign _zz_fetchStage_read_waysValues_0_tag_valid_2 = ways_0_tags_spinal_port1;
  assign fetchStage_read_waysValues_0_tag_valid = _zz_fetchStage_read_waysValues_0_tag_valid_2[0];
  assign fetchStage_read_waysValues_0_tag_error = _zz_fetchStage_read_waysValues_0_tag_valid_2[1];
  assign fetchStage_read_waysValues_0_tag_address = _zz_fetchStage_read_waysValues_0_tag_valid_2[21 : 2];
  assign _zz_fetchStage_read_waysValues_1_tag_valid = io_cpu_prefetch_pc[11 : 6];
  assign _zz_fetchStage_read_waysValues_1_tag_valid_1 = (! io_cpu_fetch_isStuck);
  assign _zz_fetchStage_read_waysValues_1_tag_valid_2 = ways_1_tags_spinal_port1;
  assign fetchStage_read_waysValues_1_tag_valid = _zz_fetchStage_read_waysValues_1_tag_valid_2[0];
  assign fetchStage_read_waysValues_1_tag_error = _zz_fetchStage_read_waysValues_1_tag_valid_2[1];
  assign fetchStage_read_waysValues_1_tag_address = _zz_fetchStage_read_waysValues_1_tag_valid_2[21 : 2];
  assign fetchStage_hit_hits_0 = (fetchStage_read_waysValues_0_tag_valid && (fetchStage_read_waysValues_0_tag_address == io_cpu_fetch_mmuRsp_physicalAddress[31 : 12]));
  assign fetchStage_hit_hits_1 = (fetchStage_read_waysValues_1_tag_valid && (fetchStage_read_waysValues_1_tag_address == io_cpu_fetch_mmuRsp_physicalAddress[31 : 12]));
  assign fetchStage_hit_valid = (|{fetchStage_hit_hits_1,fetchStage_hit_hits_0});
  assign fetchStage_hit_wayId = fetchStage_hit_hits_1;
  assign fetchStage_hit_bankId = _zz_fetchStage_hit_bankId;
  assign fetchStage_hit_error = _zz_fetchStage_hit_error;
  assign fetchStage_hit_data = _zz_fetchStage_hit_data;
  assign fetchStage_hit_word = fetchStage_hit_data;
  assign io_cpu_fetch_data = fetchStage_hit_word;
  assign when_InstructionCache_l435 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_data = io_cpu_fetch_data_regNextWhen;
  assign io_cpu_fetch_physicalAddress = io_cpu_fetch_mmuRsp_physicalAddress;
  assign when_InstructionCache_l459 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_1 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_2 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_cacheMiss = (! decodeStage_hit_valid);
  assign io_cpu_decode_error = (decodeStage_hit_error || ((! decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute))));
  assign io_cpu_decode_mmuRefilling = decodeStage_mmuRsp_refilling;
  assign io_cpu_decode_mmuException = (((! decodeStage_mmuRsp_refilling) && decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute)));
  assign io_cpu_decode_physicalAddress = decodeStage_mmuRsp_physicalAddress;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      lineLoader_valid <= 1'b0;
      lineLoader_hadError <= 1'b0;
      lineLoader_flushPending <= 1'b1;
      lineLoader_cmdSent <= 1'b0;
      lineLoader_wayToAllocate_value <= 1'b0;
      lineLoader_wordIndex <= 3'b000;
    end else begin
      if(lineLoader_fire) begin
        lineLoader_valid <= 1'b0;
      end
      if(lineLoader_fire) begin
        lineLoader_hadError <= 1'b0;
      end
      if(io_cpu_fill_valid) begin
        lineLoader_valid <= 1'b1;
      end
      if(io_flush) begin
        lineLoader_flushPending <= 1'b1;
      end
      if(when_InstructionCache_l351) begin
        lineLoader_flushPending <= 1'b0;
      end
      if(io_mem_cmd_fire) begin
        lineLoader_cmdSent <= 1'b1;
      end
      if(lineLoader_fire) begin
        lineLoader_cmdSent <= 1'b0;
      end
      lineLoader_wayToAllocate_value <= lineLoader_wayToAllocate_valueNext;
      if(io_mem_rsp_valid) begin
        lineLoader_wordIndex <= (lineLoader_wordIndex + 3'b001);
        if(io_mem_rsp_payload_error) begin
          lineLoader_hadError <= 1'b1;
        end
      end
    end
  end

  always @(posedge io_systemClk) begin
    if(io_cpu_fill_valid) begin
      lineLoader_address <= io_cpu_fill_payload;
    end
    if(when_InstructionCache_l338) begin
      lineLoader_flushCounter <= (lineLoader_flushCounter + 7'h01);
    end
    _zz_when_InstructionCache_l342 <= lineLoader_flushCounter[6];
    if(when_InstructionCache_l351) begin
      lineLoader_flushCounter <= 7'h0;
    end
    if(when_InstructionCache_l435) begin
      io_cpu_fetch_data_regNextWhen <= io_cpu_fetch_data;
    end
    if(when_InstructionCache_l459) begin
      decodeStage_mmuRsp_physicalAddress <= io_cpu_fetch_mmuRsp_physicalAddress;
      decodeStage_mmuRsp_isIoAccess <= io_cpu_fetch_mmuRsp_isIoAccess;
      decodeStage_mmuRsp_isPaging <= io_cpu_fetch_mmuRsp_isPaging;
      decodeStage_mmuRsp_allowRead <= io_cpu_fetch_mmuRsp_allowRead;
      decodeStage_mmuRsp_allowWrite <= io_cpu_fetch_mmuRsp_allowWrite;
      decodeStage_mmuRsp_allowExecute <= io_cpu_fetch_mmuRsp_allowExecute;
      decodeStage_mmuRsp_exception <= io_cpu_fetch_mmuRsp_exception;
      decodeStage_mmuRsp_refilling <= io_cpu_fetch_mmuRsp_refilling;
      decodeStage_mmuRsp_bypassTranslation <= io_cpu_fetch_mmuRsp_bypassTranslation;
    end
    if(when_InstructionCache_l459_1) begin
      decodeStage_hit_valid <= fetchStage_hit_valid;
    end
    if(when_InstructionCache_l459_2) begin
      decodeStage_hit_error <= fetchStage_hit_error;
    end
  end


endmodule

//BufferCC_51 replaced by BufferCC_46

//BufferCC_50 replaced by BufferCC_46

//BufferCC_49 replaced by BufferCC_46

//BufferCC_48 replaced by BufferCC_46

//BufferCC_47 replaced by BufferCC_46

module BufferCC_46 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module UartCtrlRx (
  input  wire [2:0]    io_configFrame_dataLength,
  input  wire [0:0]    io_configFrame_stop,
  input  wire [1:0]    io_configFrame_parity,
  input  wire          io_samplingTick,
  output wire          io_read_valid,
  input  wire          io_read_ready,
  output wire [7:0]    io_read_payload,
  input  wire          io_rxd,
  output wire          io_rts,
  output reg           io_error,
  output wire          io_break,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;
  localparam UartCtrlRxState_IDLE = 3'd0;
  localparam UartCtrlRxState_START = 3'd1;
  localparam UartCtrlRxState_DATA = 3'd2;
  localparam UartCtrlRxState_PARITY = 3'd3;
  localparam UartCtrlRxState_STOP = 3'd4;

  wire                io_rxd_buffercc_io_dataOut;
  wire                _zz_sampler_value;
  wire                _zz_sampler_value_1;
  wire                _zz_sampler_value_2;
  wire                _zz_sampler_value_3;
  wire                _zz_sampler_value_4;
  wire                _zz_sampler_value_5;
  wire                _zz_sampler_value_6;
  wire       [2:0]    _zz_when_UartCtrlRx_l139;
  wire       [0:0]    _zz_when_UartCtrlRx_l139_1;
  reg                 _zz_io_rts;
  wire                sampler_synchroniser;
  wire                sampler_samples_0;
  reg                 sampler_samples_1;
  reg                 sampler_samples_2;
  reg                 sampler_samples_3;
  reg                 sampler_samples_4;
  reg                 sampler_value;
  reg                 sampler_tick;
  reg        [2:0]    bitTimer_counter;
  reg                 bitTimer_tick;
  wire                when_UartCtrlRx_l43;
  reg        [2:0]    bitCounter_value;
  reg        [6:0]    break_counter;
  wire                break_valid;
  wire                when_UartCtrlRx_l69;
  reg        [2:0]    stateMachine_state;
  reg                 stateMachine_parity;
  reg        [7:0]    stateMachine_shifter;
  reg                 stateMachine_validReg;
  wire                when_UartCtrlRx_l93;
  wire                when_UartCtrlRx_l103;
  wire                when_UartCtrlRx_l111;
  wire                when_UartCtrlRx_l113;
  wire                when_UartCtrlRx_l125;
  wire                when_UartCtrlRx_l136;
  wire                when_UartCtrlRx_l139;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  `endif


  assign _zz_when_UartCtrlRx_l139_1 = ((io_configFrame_stop == UartStopType_ONE) ? 1'b0 : 1'b1);
  assign _zz_when_UartCtrlRx_l139 = {2'd0, _zz_when_UartCtrlRx_l139_1};
  assign _zz_sampler_value = ((((1'b0 || ((_zz_sampler_value_1 && sampler_samples_1) && sampler_samples_2)) || (((_zz_sampler_value_2 && sampler_samples_0) && sampler_samples_1) && sampler_samples_3)) || (((1'b1 && sampler_samples_0) && sampler_samples_2) && sampler_samples_3)) || (((1'b1 && sampler_samples_1) && sampler_samples_2) && sampler_samples_3));
  assign _zz_sampler_value_3 = (((1'b1 && sampler_samples_0) && sampler_samples_1) && sampler_samples_4);
  assign _zz_sampler_value_4 = ((1'b1 && sampler_samples_0) && sampler_samples_2);
  assign _zz_sampler_value_5 = (1'b1 && sampler_samples_1);
  assign _zz_sampler_value_6 = 1'b1;
  assign _zz_sampler_value_1 = (1'b1 && sampler_samples_0);
  assign _zz_sampler_value_2 = 1'b1;
  (* keep_hierarchy = "TRUE" *) BufferCC_45 io_rxd_buffercc (
    .io_dataIn                      (io_rxd                        ), //i
    .io_dataOut                     (io_rxd_buffercc_io_dataOut    ), //o
    .io_peripheralClk               (io_peripheralClk              ), //i
    .peripheralCd_logic_outputReset (peripheralCd_logic_outputReset)  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      UartStopType_ONE : io_configFrame_stop_string = "ONE";
      UartStopType_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      UartParityType_NONE : io_configFrame_parity_string = "NONE";
      UartParityType_EVEN : io_configFrame_parity_string = "EVEN";
      UartParityType_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      UartCtrlRxState_IDLE : stateMachine_state_string = "IDLE  ";
      UartCtrlRxState_START : stateMachine_state_string = "START ";
      UartCtrlRxState_DATA : stateMachine_state_string = "DATA  ";
      UartCtrlRxState_PARITY : stateMachine_state_string = "PARITY";
      UartCtrlRxState_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    io_error = 1'b0;
    case(stateMachine_state)
      UartCtrlRxState_IDLE : begin
      end
      UartCtrlRxState_START : begin
      end
      UartCtrlRxState_DATA : begin
      end
      UartCtrlRxState_PARITY : begin
        if(bitTimer_tick) begin
          if(!when_UartCtrlRx_l125) begin
            io_error = 1'b1;
          end
        end
      end
      default : begin
        if(bitTimer_tick) begin
          if(when_UartCtrlRx_l136) begin
            io_error = 1'b1;
          end
        end
      end
    endcase
  end

  assign io_rts = _zz_io_rts;
  assign sampler_synchroniser = io_rxd_buffercc_io_dataOut;
  assign sampler_samples_0 = sampler_synchroniser;
  always @(*) begin
    bitTimer_tick = 1'b0;
    if(sampler_tick) begin
      if(when_UartCtrlRx_l43) begin
        bitTimer_tick = 1'b1;
      end
    end
  end

  assign when_UartCtrlRx_l43 = (bitTimer_counter == 3'b000);
  assign break_valid = (break_counter == 7'h68);
  assign when_UartCtrlRx_l69 = (io_samplingTick && (! break_valid));
  assign io_break = break_valid;
  assign io_read_valid = stateMachine_validReg;
  assign when_UartCtrlRx_l93 = ((sampler_tick && (! sampler_value)) && (! break_valid));
  assign when_UartCtrlRx_l103 = (sampler_value == 1'b1);
  assign when_UartCtrlRx_l111 = (bitCounter_value == io_configFrame_dataLength);
  assign when_UartCtrlRx_l113 = (io_configFrame_parity == UartParityType_NONE);
  assign when_UartCtrlRx_l125 = (stateMachine_parity == sampler_value);
  assign when_UartCtrlRx_l136 = (! sampler_value);
  assign when_UartCtrlRx_l139 = (bitCounter_value == _zz_when_UartCtrlRx_l139);
  assign io_read_payload = stateMachine_shifter;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      _zz_io_rts <= 1'b0;
      sampler_samples_1 <= 1'b1;
      sampler_samples_2 <= 1'b1;
      sampler_samples_3 <= 1'b1;
      sampler_samples_4 <= 1'b1;
      sampler_value <= 1'b1;
      sampler_tick <= 1'b0;
      break_counter <= 7'h0;
      stateMachine_state <= UartCtrlRxState_IDLE;
      stateMachine_validReg <= 1'b0;
    end else begin
      _zz_io_rts <= (! io_read_ready);
      if(io_samplingTick) begin
        sampler_samples_1 <= sampler_samples_0;
      end
      if(io_samplingTick) begin
        sampler_samples_2 <= sampler_samples_1;
      end
      if(io_samplingTick) begin
        sampler_samples_3 <= sampler_samples_2;
      end
      if(io_samplingTick) begin
        sampler_samples_4 <= sampler_samples_3;
      end
      sampler_value <= ((((((_zz_sampler_value || _zz_sampler_value_3) || (_zz_sampler_value_4 && sampler_samples_4)) || ((_zz_sampler_value_5 && sampler_samples_2) && sampler_samples_4)) || (((_zz_sampler_value_6 && sampler_samples_0) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_1) && sampler_samples_3) && sampler_samples_4)) || (((1'b1 && sampler_samples_2) && sampler_samples_3) && sampler_samples_4));
      sampler_tick <= io_samplingTick;
      if(sampler_value) begin
        break_counter <= 7'h0;
      end else begin
        if(when_UartCtrlRx_l69) begin
          break_counter <= (break_counter + 7'h01);
        end
      end
      stateMachine_validReg <= 1'b0;
      case(stateMachine_state)
        UartCtrlRxState_IDLE : begin
          if(when_UartCtrlRx_l93) begin
            stateMachine_state <= UartCtrlRxState_START;
          end
        end
        UartCtrlRxState_START : begin
          if(bitTimer_tick) begin
            stateMachine_state <= UartCtrlRxState_DATA;
            if(when_UartCtrlRx_l103) begin
              stateMachine_state <= UartCtrlRxState_IDLE;
            end
          end
        end
        UartCtrlRxState_DATA : begin
          if(bitTimer_tick) begin
            if(when_UartCtrlRx_l111) begin
              if(when_UartCtrlRx_l113) begin
                stateMachine_state <= UartCtrlRxState_STOP;
                stateMachine_validReg <= 1'b1;
              end else begin
                stateMachine_state <= UartCtrlRxState_PARITY;
              end
            end
          end
        end
        UartCtrlRxState_PARITY : begin
          if(bitTimer_tick) begin
            if(when_UartCtrlRx_l125) begin
              stateMachine_state <= UartCtrlRxState_STOP;
              stateMachine_validReg <= 1'b1;
            end else begin
              stateMachine_state <= UartCtrlRxState_IDLE;
            end
          end
        end
        default : begin
          if(bitTimer_tick) begin
            if(when_UartCtrlRx_l136) begin
              stateMachine_state <= UartCtrlRxState_IDLE;
            end else begin
              if(when_UartCtrlRx_l139) begin
                stateMachine_state <= UartCtrlRxState_IDLE;
              end
            end
          end
        end
      endcase
    end
  end

  always @(posedge io_peripheralClk) begin
    if(sampler_tick) begin
      bitTimer_counter <= (bitTimer_counter - 3'b001);
    end
    if(bitTimer_tick) begin
      bitCounter_value <= (bitCounter_value + 3'b001);
    end
    if(bitTimer_tick) begin
      stateMachine_parity <= (stateMachine_parity ^ sampler_value);
    end
    case(stateMachine_state)
      UartCtrlRxState_IDLE : begin
        if(when_UartCtrlRx_l93) begin
          bitTimer_counter <= 3'b010;
        end
      end
      UartCtrlRxState_START : begin
        if(bitTimer_tick) begin
          bitCounter_value <= 3'b000;
          stateMachine_parity <= (io_configFrame_parity == UartParityType_ODD);
        end
      end
      UartCtrlRxState_DATA : begin
        if(bitTimer_tick) begin
          stateMachine_shifter[bitCounter_value] <= sampler_value;
          if(when_UartCtrlRx_l111) begin
            bitCounter_value <= 3'b000;
          end
        end
      end
      UartCtrlRxState_PARITY : begin
        if(bitTimer_tick) begin
          bitCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module UartCtrlTx (
  input  wire [2:0]    io_configFrame_dataLength,
  input  wire [0:0]    io_configFrame_stop,
  input  wire [1:0]    io_configFrame_parity,
  input  wire          io_samplingTick,
  input  wire          io_write_valid,
  output reg           io_write_ready,
  input  wire [7:0]    io_write_payload,
  input  wire          io_cts,
  output wire          io_txd,
  input  wire          io_break,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);
  localparam UartStopType_ONE = 1'd0;
  localparam UartStopType_TWO = 1'd1;
  localparam UartParityType_NONE = 2'd0;
  localparam UartParityType_EVEN = 2'd1;
  localparam UartParityType_ODD = 2'd2;
  localparam UartCtrlTxState_IDLE = 3'd0;
  localparam UartCtrlTxState_START = 3'd1;
  localparam UartCtrlTxState_DATA = 3'd2;
  localparam UartCtrlTxState_PARITY = 3'd3;
  localparam UartCtrlTxState_STOP = 3'd4;

  wire       [2:0]    _zz_clockDivider_counter_valueNext;
  wire       [0:0]    _zz_clockDivider_counter_valueNext_1;
  wire       [2:0]    _zz_when_UartCtrlTx_l93;
  wire       [0:0]    _zz_when_UartCtrlTx_l93_1;
  reg                 clockDivider_counter_willIncrement;
  wire                clockDivider_counter_willClear;
  reg        [2:0]    clockDivider_counter_valueNext;
  reg        [2:0]    clockDivider_counter_value;
  wire                clockDivider_counter_willOverflowIfInc;
  wire                clockDivider_counter_willOverflow;
  reg        [2:0]    tickCounter_value;
  reg        [2:0]    stateMachine_state;
  reg                 stateMachine_parity;
  reg                 stateMachine_txd;
  wire                when_UartCtrlTx_l58;
  wire                when_UartCtrlTx_l73;
  wire                when_UartCtrlTx_l76;
  wire                when_UartCtrlTx_l93;
  wire       [2:0]    _zz_stateMachine_state;
  reg                 _zz_io_txd;
  `ifndef SYNTHESIS
  reg [23:0] io_configFrame_stop_string;
  reg [31:0] io_configFrame_parity_string;
  reg [47:0] stateMachine_state_string;
  reg [47:0] _zz_stateMachine_state_string;
  `endif


  assign _zz_clockDivider_counter_valueNext_1 = clockDivider_counter_willIncrement;
  assign _zz_clockDivider_counter_valueNext = {2'd0, _zz_clockDivider_counter_valueNext_1};
  assign _zz_when_UartCtrlTx_l93_1 = ((io_configFrame_stop == UartStopType_ONE) ? 1'b0 : 1'b1);
  assign _zz_when_UartCtrlTx_l93 = {2'd0, _zz_when_UartCtrlTx_l93_1};
  `ifndef SYNTHESIS
  always @(*) begin
    case(io_configFrame_stop)
      UartStopType_ONE : io_configFrame_stop_string = "ONE";
      UartStopType_TWO : io_configFrame_stop_string = "TWO";
      default : io_configFrame_stop_string = "???";
    endcase
  end
  always @(*) begin
    case(io_configFrame_parity)
      UartParityType_NONE : io_configFrame_parity_string = "NONE";
      UartParityType_EVEN : io_configFrame_parity_string = "EVEN";
      UartParityType_ODD : io_configFrame_parity_string = "ODD ";
      default : io_configFrame_parity_string = "????";
    endcase
  end
  always @(*) begin
    case(stateMachine_state)
      UartCtrlTxState_IDLE : stateMachine_state_string = "IDLE  ";
      UartCtrlTxState_START : stateMachine_state_string = "START ";
      UartCtrlTxState_DATA : stateMachine_state_string = "DATA  ";
      UartCtrlTxState_PARITY : stateMachine_state_string = "PARITY";
      UartCtrlTxState_STOP : stateMachine_state_string = "STOP  ";
      default : stateMachine_state_string = "??????";
    endcase
  end
  always @(*) begin
    case(_zz_stateMachine_state)
      UartCtrlTxState_IDLE : _zz_stateMachine_state_string = "IDLE  ";
      UartCtrlTxState_START : _zz_stateMachine_state_string = "START ";
      UartCtrlTxState_DATA : _zz_stateMachine_state_string = "DATA  ";
      UartCtrlTxState_PARITY : _zz_stateMachine_state_string = "PARITY";
      UartCtrlTxState_STOP : _zz_stateMachine_state_string = "STOP  ";
      default : _zz_stateMachine_state_string = "??????";
    endcase
  end
  `endif

  always @(*) begin
    clockDivider_counter_willIncrement = 1'b0;
    if(io_samplingTick) begin
      clockDivider_counter_willIncrement = 1'b1;
    end
  end

  assign clockDivider_counter_willClear = 1'b0;
  assign clockDivider_counter_willOverflowIfInc = (clockDivider_counter_value == 3'b111);
  assign clockDivider_counter_willOverflow = (clockDivider_counter_willOverflowIfInc && clockDivider_counter_willIncrement);
  always @(*) begin
    clockDivider_counter_valueNext = (clockDivider_counter_value + _zz_clockDivider_counter_valueNext);
    if(clockDivider_counter_willClear) begin
      clockDivider_counter_valueNext = 3'b000;
    end
  end

  always @(*) begin
    stateMachine_txd = 1'b1;
    case(stateMachine_state)
      UartCtrlTxState_IDLE : begin
      end
      UartCtrlTxState_START : begin
        stateMachine_txd = 1'b0;
      end
      UartCtrlTxState_DATA : begin
        stateMachine_txd = io_write_payload[tickCounter_value];
      end
      UartCtrlTxState_PARITY : begin
        stateMachine_txd = stateMachine_parity;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_write_ready = io_break;
    case(stateMachine_state)
      UartCtrlTxState_IDLE : begin
      end
      UartCtrlTxState_START : begin
      end
      UartCtrlTxState_DATA : begin
        if(clockDivider_counter_willOverflow) begin
          if(when_UartCtrlTx_l73) begin
            io_write_ready = 1'b1;
          end
        end
      end
      UartCtrlTxState_PARITY : begin
      end
      default : begin
      end
    endcase
  end

  assign when_UartCtrlTx_l58 = ((io_write_valid && (! io_cts)) && clockDivider_counter_willOverflow);
  assign when_UartCtrlTx_l73 = (tickCounter_value == io_configFrame_dataLength);
  assign when_UartCtrlTx_l76 = (io_configFrame_parity == UartParityType_NONE);
  assign when_UartCtrlTx_l93 = (tickCounter_value == _zz_when_UartCtrlTx_l93);
  assign _zz_stateMachine_state = (io_write_valid ? UartCtrlTxState_START : UartCtrlTxState_IDLE);
  assign io_txd = _zz_io_txd;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      clockDivider_counter_value <= 3'b000;
      stateMachine_state <= UartCtrlTxState_IDLE;
      _zz_io_txd <= 1'b1;
    end else begin
      clockDivider_counter_value <= clockDivider_counter_valueNext;
      case(stateMachine_state)
        UartCtrlTxState_IDLE : begin
          if(when_UartCtrlTx_l58) begin
            stateMachine_state <= UartCtrlTxState_START;
          end
        end
        UartCtrlTxState_START : begin
          if(clockDivider_counter_willOverflow) begin
            stateMachine_state <= UartCtrlTxState_DATA;
          end
        end
        UartCtrlTxState_DATA : begin
          if(clockDivider_counter_willOverflow) begin
            if(when_UartCtrlTx_l73) begin
              if(when_UartCtrlTx_l76) begin
                stateMachine_state <= UartCtrlTxState_STOP;
              end else begin
                stateMachine_state <= UartCtrlTxState_PARITY;
              end
            end
          end
        end
        UartCtrlTxState_PARITY : begin
          if(clockDivider_counter_willOverflow) begin
            stateMachine_state <= UartCtrlTxState_STOP;
          end
        end
        default : begin
          if(clockDivider_counter_willOverflow) begin
            if(when_UartCtrlTx_l93) begin
              stateMachine_state <= _zz_stateMachine_state;
            end
          end
        end
      endcase
      _zz_io_txd <= (stateMachine_txd && (! io_break));
    end
  end

  always @(posedge io_peripheralClk) begin
    if(clockDivider_counter_willOverflow) begin
      tickCounter_value <= (tickCounter_value + 3'b001);
    end
    if(clockDivider_counter_willOverflow) begin
      stateMachine_parity <= (stateMachine_parity ^ stateMachine_txd);
    end
    case(stateMachine_state)
      UartCtrlTxState_IDLE : begin
      end
      UartCtrlTxState_START : begin
        if(clockDivider_counter_willOverflow) begin
          stateMachine_parity <= (io_configFrame_parity == UartParityType_ODD);
          tickCounter_value <= 3'b000;
        end
      end
      UartCtrlTxState_DATA : begin
        if(clockDivider_counter_willOverflow) begin
          if(when_UartCtrlTx_l73) begin
            tickCounter_value <= 3'b000;
          end
        end
      end
      UartCtrlTxState_PARITY : begin
        if(clockDivider_counter_willOverflow) begin
          tickCounter_value <= 3'b000;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module BufferCC_44 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_systemClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    if(system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized_1) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_43 replaced by BufferCC_45

module BufferCC_42 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk) begin
    if(system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized_1) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_41 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_40 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_systemClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    if(system_bridge_bmb_crossClock_toplevel_peripheralCd_logic_outputReset_synchronized) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_39 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_systemClk,
  input  wire          peripheralCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk or posedge peripheralCd_logic_outputReset) begin
    if(peripheralCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_38 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_37 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk) begin
    if(system_bridge_bmb_crossClock_toplevel_systemCd_logic_outputReset_synchronized) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_36 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          systemCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk or posedge systemCd_logic_outputReset) begin
    if(systemCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_35 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//StreamFifo_5 replaced by StreamFifo_4

module BufferCC_34 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_ddrMasters_0_clk,
  input  wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_0_clk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_33 replaced by BufferCC_14

//BufferCC_32 replaced by BufferCC_30

//BufferCC_31 replaced by BufferCC_23

module BufferCC_30 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized_1) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_29 replaced by BufferCC_23

module BufferCC_28 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_ddrMasters_0_clk,
  input  wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_0_clk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_ddrCd_logic_outputReset_synchronized) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_27 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_ddrMasters_0_clk,
  input  wire          ddrCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_0_clk or posedge ddrCd_logic_outputReset) begin
    if(ddrCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_26 replaced by BufferCC_14

module BufferCC_25 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_1_bridge_toplevel_io_ddrMasters_0_reset_synchronized) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_24 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_memoryClk,
  input  wire          io_ddrMasters_0_reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk or posedge io_ddrMasters_0_reset) begin
    if(io_ddrMasters_0_reset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_23 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_ddrMasters_0_clk,
  input  wire          io_ddrMasters_0_reset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_0_clk) begin
    if(io_ddrMasters_0_reset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module StreamFifo_4 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [3:0]    io_push_payload_startAt,
  input  wire [3:0]    io_push_payload_endAt,
  input  wire [2:0]    io_push_payload_size,
  input  wire [3:0]    io_push_payload_id,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [3:0]    io_pop_payload_startAt,
  output wire [3:0]    io_pop_payload_endAt,
  output wire [2:0]    io_pop_payload_size,
  output wire [3:0]    io_pop_payload_id,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  reg        [14:0]   logic_ram_spinal_port1;
  wire       [14:0]   _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [3:0]    logic_push_onRam_write_payload_data_startAt;
  wire       [3:0]    logic_push_onRam_write_payload_data_endAt;
  wire       [2:0]    logic_push_onRam_write_payload_data_size;
  wire       [3:0]    logic_push_onRam_write_payload_data_id;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [1:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [1:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [1:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [3:0]    logic_pop_sync_readPort_rsp_startAt;
  wire       [3:0]    logic_pop_sync_readPort_rsp_endAt;
  wire       [2:0]    logic_pop_sync_readPort_rsp_size;
  wire       [3:0]    logic_pop_sync_readPort_rsp_id;
  wire       [14:0]   _zz_logic_pop_sync_readPort_rsp_startAt;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_startAt;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_endAt;
  wire       [2:0]    logic_pop_sync_readArbitation_translated_payload_size;
  wire       [3:0]    logic_pop_sync_readArbitation_translated_payload_id;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [2:0]    logic_pop_sync_popReg;
  reg [14:0] logic_ram [0:3];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_id,{logic_push_onRam_write_payload_data_size,{logic_push_onRam_write_payload_data_endAt,logic_push_onRam_write_payload_data_startAt}}};
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge io_memoryClk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 3'b100) == 3'b000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[1:0];
  assign logic_push_onRam_write_payload_data_startAt = io_push_payload_startAt;
  assign logic_push_onRam_write_payload_data_endAt = io_push_payload_endAt;
  assign logic_push_onRam_write_payload_data_size = io_push_payload_size;
  assign logic_push_onRam_write_payload_data_id = io_push_payload_id;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[1:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_startAt = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_startAt = _zz_logic_pop_sync_readPort_rsp_startAt[3 : 0];
  assign logic_pop_sync_readPort_rsp_endAt = _zz_logic_pop_sync_readPort_rsp_startAt[7 : 4];
  assign logic_pop_sync_readPort_rsp_size = _zz_logic_pop_sync_readPort_rsp_startAt[10 : 8];
  assign logic_pop_sync_readPort_rsp_id = _zz_logic_pop_sync_readPort_rsp_startAt[14 : 11];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_startAt = logic_pop_sync_readPort_rsp_startAt;
  assign logic_pop_sync_readArbitation_translated_payload_endAt = logic_pop_sync_readPort_rsp_endAt;
  assign logic_pop_sync_readArbitation_translated_payload_size = logic_pop_sync_readPort_rsp_size;
  assign logic_pop_sync_readArbitation_translated_payload_id = logic_pop_sync_readPort_rsp_id;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_startAt = logic_pop_sync_readArbitation_translated_payload_startAt;
  assign io_pop_payload_endAt = logic_pop_sync_readArbitation_translated_payload_endAt;
  assign io_pop_payload_size = logic_pop_sync_readArbitation_translated_payload_size;
  assign io_pop_payload_id = logic_pop_sync_readArbitation_translated_payload_id;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b100 - logic_ptr_occupancy);
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 3'b000;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 3'b000;
      end
    end
  end

  always @(posedge io_memoryClk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule

module BufferCC_22 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_ddrMasters_1_clk,
  input  wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_1_clk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized_1) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_21 replaced by BufferCC_14

//BufferCC_20 replaced by BufferCC_18

//BufferCC_19 replaced by BufferCC_11

module BufferCC_18 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized_1) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

//BufferCC_17 replaced by BufferCC_11

module BufferCC_16 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_ddrMasters_1_clk,
  input  wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_1_clk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_ddrCd_logic_outputReset_synchronized) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_15 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_ddrMasters_1_clk,
  input  wire          ddrCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_1_clk or posedge ddrCd_logic_outputReset) begin
    if(ddrCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_14 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_13 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_userAdapters_0_bridge_toplevel_io_ddrMasters_1_reset_synchronized) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_12 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_memoryClk,
  input  wire          io_ddrMasters_1_reset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk or posedge io_ddrMasters_1_reset) begin
    if(io_ddrMasters_1_reset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_11 (
  input  wire [4:0]    io_dataIn,
  output wire [4:0]    io_dataOut,
  input  wire          io_ddrMasters_1_clk,
  input  wire          io_ddrMasters_1_reset
);

  (* async_reg = "true" *) reg        [4:0]    buffers_0;
  (* async_reg = "true" *) reg        [4:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_ddrMasters_1_clk) begin
    if(io_ddrMasters_1_reset) begin
      buffers_0 <= 5'h0;
      buffers_1 <= 5'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module StreamFifo_3 (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [1:0]    io_push_payload,
  output reg           io_pop_valid,
  input  wire          io_pop_ready,
  output reg  [1:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  wire       [1:0]    logic_ram_spinal_port1;
  wire       [1:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  reg                 logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [1:0]    logic_push_onRam_write_payload_data;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [1:0]    logic_pop_async_readed;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [1:0]    logic_pop_addressGen_translated_payload;
  (* ram_style = "distributed" *) reg [1:0] logic_ram [0:3];

  assign _zz_logic_ram_port = logic_push_onRam_write_payload_data;
  always @(posedge io_memoryClk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  assign logic_ram_spinal_port1 = logic_ram[logic_pop_addressGen_payload];
  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 3'b100) == 3'b000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  always @(*) begin
    logic_ptr_doPush = io_push_fire;
    if(logic_ptr_empty) begin
      if(io_pop_ready) begin
        logic_ptr_doPush = 1'b0;
      end
    end
  end

  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[1:0];
  assign logic_push_onRam_write_payload_data = io_push_payload;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[1:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign logic_pop_async_readed = logic_ram_spinal_port1;
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload = logic_pop_async_readed;
  always @(*) begin
    io_pop_valid = logic_pop_addressGen_translated_valid;
    if(logic_ptr_empty) begin
      io_pop_valid = io_push_valid;
    end
  end

  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  always @(*) begin
    io_pop_payload = logic_pop_addressGen_translated_payload;
    if(logic_ptr_empty) begin
      io_pop_payload = io_push_payload;
    end
  end

  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b100 - logic_ptr_occupancy);
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
    end
  end


endmodule

module BufferCC_10 (
  input  wire [6:0]    io_dataIn,
  output wire [6:0]    io_dataOut,
  input  wire          io_systemClk,
  input  wire          system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_synchronized
);

  (* async_reg = "true" *) reg        [6:0]    buffers_0;
  (* async_reg = "true" *) reg        [6:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    if(system_ddr_ddrLogic_cc_fifo_toplevel_ddrCd_logic_outputReset_synchronized) begin
      buffers_0 <= 7'h0;
      buffers_1 <= 7'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_9 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_systemClk,
  input  wire          ddrCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk or posedge ddrCd_logic_outputReset) begin
    if(ddrCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_8 (
  input  wire [6:0]    io_dataIn,
  output wire [6:0]    io_dataOut,
  input  wire          io_memoryClk,
  input  wire          ddrCd_logic_outputReset
);

  (* async_reg = "true" *) reg        [6:0]    buffers_0;
  (* async_reg = "true" *) reg        [6:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk) begin
    if(ddrCd_logic_outputReset) begin
      buffers_0 <= 7'h0;
      buffers_1 <= 7'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_7 (
  input  wire [6:0]    io_dataIn,
  output wire [6:0]    io_dataOut,
  input  wire          io_memoryClk,
  input  wire          system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_synchronized
);

  (* async_reg = "true" *) reg        [6:0]    buffers_0;
  (* async_reg = "true" *) reg        [6:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk) begin
    if(system_ddr_ddrLogic_cc_fifo_toplevel_systemCd_logic_outputReset_synchronized) begin
      buffers_0 <= 7'h0;
      buffers_1 <= 7'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_6 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_memoryClk,
  input  wire          systemCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_memoryClk or posedge systemCd_logic_outputReset) begin
    if(systemCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_5 (
  input  wire [6:0]    io_dataIn,
  output wire [6:0]    io_dataOut,
  input  wire          io_systemClk,
  input  wire          systemCd_logic_outputReset
);

  (* async_reg = "true" *) reg        [6:0]    buffers_0;
  (* async_reg = "true" *) reg        [6:0]    buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    if(systemCd_logic_outputReset) begin
      buffers_0 <= 7'h0;
      buffers_1 <= 7'h0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_4 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          jtagCtrl_tck,
  input  wire          system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_synchronized
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge jtagCtrl_tck) begin
    if(system_riscvJtag_hard_noTap_tunnel_toplevel_debugCd_logic_outputReset_synchronized) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_3 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          jtagCtrl_tck,
  input  wire          debugCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge jtagCtrl_tck or posedge debugCd_logic_outputReset) begin
    if(debugCd_logic_outputReset) begin
      buffers_0 <= 1'b1;
      buffers_1 <= 1'b1;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module BufferCC_2 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_systemClk,
  input  wire          debugCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  initial begin
  `ifndef SYNTHESIS
    buffers_0 = $urandom;
    buffers_1 = $urandom;
  `endif
  end

  assign io_dataOut = buffers_1;
  always @(posedge io_systemClk) begin
    buffers_0 <= io_dataIn;
    buffers_1 <= buffers_0;
  end


endmodule

module BufferCC_45 (
  input  wire          io_dataIn,
  output wire          io_dataOut,
  input  wire          io_peripheralClk,
  input  wire          peripheralCd_logic_outputReset
);

  (* async_reg = "true" *) reg                 buffers_0;
  (* async_reg = "true" *) reg                 buffers_1;

  assign io_dataOut = buffers_1;
  always @(posedge io_peripheralClk) begin
    if(peripheralCd_logic_outputReset) begin
      buffers_0 <= 1'b0;
      buffers_1 <= 1'b0;
    end else begin
      buffers_0 <= io_dataIn;
      buffers_1 <= buffers_0;
    end
  end


endmodule

module EfxCPUSp1 (
  input      [31:0]   src1,
  input      [31:0]   src2,
  input      [1:0]    bitCtrl,
  input      [1:0]    ctrl,
  input               less,
  input      [31:0]   addSub,
  output     [31:0]   result
);
//pragma protect
//pragma protect begin
`protected

    MTI!#ev'YC=3VR]zU,'{]UA[2JXU{As+pV?pk=~oA\]"#e=]e,Rl2-2Uok2[]~B\r^3;^YW2~UV*
    rpUWe3U+a{@]Uw@oaaj'}muo_Y~@U_hw>WC<I{WU1n'a+-3Xv[OTGR7lR?pj$VZD!'GjvrDrk5}i
    {Zrjv!2:?+G<r^5}Du@=*Gv]WlR'JsHlmTJRzj]2OuK?a$<T{1$]^JJJ<E!JoTAvOCWnRT\]_e{s
    {->}jFxvI7tp^JkZUp{yJGaVJUu>$nZQ^-1;c*aV'^nxJ\kq@x}-^x~X}\2zf;YDn']J}P><I!|[
    Ja[uv@WC2Qn&u=ZKg3U$3r?R_.}-DEZE-nV~eA|Up,^VOuVu^3CCn23On5!<^#+5{l2pUI7K==!2
    -+Wr$ssZj,i;<zoDx'5UAA?6T,U-rD-z%<XQV]?2IW7]pYm=>^s?1@ED^nsz@[cmE~#C=TT]_<C5
    D~CkAYv#e[EFl-TZ7lY^}7QD{a$o^_;s?w@OtIiTKveYpLnHWU=]K$Y*ZkBY^KnaB#%Q&B~przx\
    ,DRAnnQa^mXr[$hu_@^o-7Qk=@^*]=BnBi]JD-^!wosQ']5v[]umICCn+}!;1_YOR,wj2vXxT==1
    1]HXoIrelT!-^1*EB~aKTujJE2kp7?CBT}G7*=j2CjA2\B}=Ao2CKjoJvI3B^{jbtwE!]kU'w-VC
    z2$C7>Gll$ZTsEWa3h^u-IE}OJ1tt:sI$ZVGj{_<<#QKo,sT>R6]e'$k]?YFTX<Y\<>TRpHOl$#_
    X]!r;UZ7[s=A+{CJEJ},swWA$!2^EmZJCe,vnwj=$ZWnP>Er-R=kz?EQ~!s~G8pCm,BY1pJ,rA}J
    {DK=Es<][
`endprotected
//pragma protect end

module EfxCPUSp2 (
  input      [1:0]    ctrl,
  input      [31:0]   src1,
  input      [31:0]   src2,
  output     [31:0]   result
);
//pragma protect
//pragma protect begin
`protected

    MTI!#[o$Tj!IrkR5nYBXe=xpn*3xBG$Gm1C,$|.><{[y*\Ua,;U*<,z^=wH5Z$#'xVOTpnp*yel~
    2=?*;X=kQ5='<,aWze+B;\rBC[W*?:QrG2}A!R?+3BLoU;Qp!7CyOgcRI[ol,BeXvDeD_W<ppCpq
    O;U!Yo^^oWY@'5YUsOElQzIV}iOJl'+$XwO[xjH,5B*=C!Q<HAjw<vuB$J3+9x#5*I?~JoaK~COp
    }IHDlnU~KC};?gN>[/xn'7^M~j[IA5kB^QkG<]_\pgt/Yo@oH+~QHUE$#'QrU1[JY,Ezpm_,#}!H
    1}aUcU|,r?w#-riJYBI}k++oon[.[@!W-T_7bCm~lm<U3,#A[3T{#o_m1+riH\J,~uj?#KaW!f=I
    iQ}$JCcYsY'|Az!-B'ER']A!S@5w^^_U[1,O~CnVls;]J=k!?yV-{^vvxosZoielK;=<C,1\$nU'
    Ku=1<X>vJOG7-Y9(lY-}*3$IeO+$O+p'ysJK{!{{R0X-U2l5i'&l9$B2~l3@H3E5=2jZ!w_mniEp
    lYX,uIUjUPvBjrVQQAoY,V1l~{elklH+z13E5'I+awaszip]WVCB^mUjUwGv1XC^BRr-K5~TnCvK
    7]2GkT][@Ui{Bw=\WYQvsmK{BC&kD]7n,YH=BXa=Q^ZWvKk[>Y*2+^*9Grr$AI^p{}2\IGJm{<+a
    mIK\[3{r7D^5,zS=mK__oA'IkWoVK<ozVG3_1[+i^'Ys,<zXssU_'Avz+xGo@*z{1rKWsJx/&1^R
    21+EW>B8B,V+Do7KC!7W'V*O}YA]}l@!~zO<x57?H,M7D'\F=^eAy5]+}Lpns!U{{\D,@zmnD-s@
    XJU<5pQao$s{,OW_O[)i+ExG_D=K$r!*\nn,evQ3'}HJsl>77J]HD7p93l-H-]DvxupoC@mD+Esx
    QGYp,5Hzk$[eJRVioZCT}'YKXrj{JrEz%^s$C,z}>#'=13s*$B?D{'rR+moWO}$+2vwTVsmX5YD<
    <[\rQCo5}e~A^2\CD^BQ?%R_\?JnIUl}<AvJKpHeG[Cjomr^{TJVxUEAl>,=$nmR3lHvsJ]_JGGz
    R?@&e@3BzJ]l,GiXMa+GnD*mZi{s*p32R"$%jU^Ds+U
`endprotected
//pragma protect end

