localparam M_BASE_ADDR = {32'h41000000,32'h40000000,32'h30000000,32'h20000000,32'h11100000,32'h810000,32'h800000,32'h0};
localparam M_ADDR_WIDTH = {32'd20,32'd24,32'd28,32'd28,32'd20,32'd16,32'd16,32'd23};